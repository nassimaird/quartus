-- niosvprocessor_tb.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosvprocessor_tb is
end entity niosvprocessor_tb;

architecture rtl of niosvprocessor_tb is
	component niosvprocessor is
		port (
			clk_clk : in std_logic := 'X'  -- clk
		);
	end component niosvprocessor;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	signal niosvprocessor_inst_clk_bfm_clk_clk : std_logic; -- niosvprocessor_inst_clk_bfm:clk -> niosvprocessor_inst:clk_clk

begin

	niosvprocessor_inst : component niosvprocessor
		port map (
			clk_clk => niosvprocessor_inst_clk_bfm_clk_clk  -- clk.clk
		);

	niosvprocessor_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => niosvprocessor_inst_clk_bfm_clk_clk  -- clk.clk
		);

end architecture rtl; -- of niosvprocessor_tb
