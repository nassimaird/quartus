`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rLaQPMZvFarXZMvrUWnIj3bRX/Yxuf2+BbmiQlMUR36vCoB4EQyjm7hU79xIBV5a
N7XdPe6/8mPcxIw8zL9+Kr3noTs9f9Iw8AML7+noNrivqZSl+U66uCVLUX2GZpvh
uZUajns+glR0v/F5Aq6by9ByoJweBeHp99JkMXstOtY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11232)
rQfBhSxvJwxFhvzumGbcUx6N7JZFlMkjECpXfQHgAsYWpVFQp4r+X+rKl9aRyO+N
l9latJKr2kLVw9u/mKXT6avVKwKTDdumZaZD/R2pyoHJomxhaA7Yu4q7c6wZfsJH
6wwEiTyxHRZjmJBa6lZev8mubCZLAUduV1Ddy7exmdOq7Wg9kHUApsSrtLHF6+lB
wmnl5IYOsjtlxSokVUyFQDa9/9vYm3Npah71Qc5zJSUiidbSoX1q9ggPym2EcDMy
5WKbfsyt8pdxduL+rT+gqW3TFd/caxikjg24k29YFwaTBnHMZyfWugiUjjugJQkX
tMou+ZM2/nkHWVFYJkJI2J4rGqGupc3rQtUmuDNVh+Vn7XHd1gFIWBcb/X0hQLhe
AmBpSDS2qyRtxoqvrHQEsPNqxFIQNt3xY1LyMM0nyDL1voPN/505wQywLmcQtcf6
Gu7B1PrNbXNc0AoMvnSzkz3dHdXqIjHC5ip5LF1XADsbzD35PfQkbeb1oHX91oDm
GyOBfJxn86xe8hO+rZDi10I5XyRatAR/ZEcXARDJIHmAHH3NlqvJEohdBHBmFTOo
u/h1PJHsDFk7UJBFeAGYyuuoM68bm9Wb9fzZ+Gtj6NBZT6Rf/r7yyQgOXVnAj7in
goDtxzW0D83Hi69PbyiVjBOpHfxfLNLUdNkCUTlTZ0Tbmr2qv8pAmitcVRhgr3cL
x4CGqxiFr/LTtj6HYs8KE0DV51cpyd55bMAL0BeqpgptT/BaAWff5cnmtEeIuEiQ
fjgNugNXVdW28I8NWJ+wo7HUaT1ECmPRETLSLtd6hQiamlWtxhft3f9kyXpTRoh+
90iAusVwaJVUqTePljyBcQruoboOL2EoZ655iy5ceAyOs5cL30ePg+SmtzthBkOW
n+nmM1aieDo3qFZA8KfvbFZLtz8zqsD9EIMqYDxGBAV4oy6Pdl86r+anzGKny0IW
o8ry4f063hr0vKaSux6wPV2InF+S68RLe8VLNiUd1DG4F4xnGaedXEdOaUbZJ3dk
/Rvfn6ljVpCs3/Mv7qMHngntyiwLiumg/is2JnuPf6HJDj2TYvFnNXM/Z+nL0Tuu
JAT+vCghUnlnWzLi1JKFDrKGuwtTCJTlK8hlNQ+y/4llEdCaGz9laC/IDzM4LTcm
qXFF0RtBugIwoIfXgDxbzI8JdnJEDdoz+6nCZ9RXvcI82qfI6uPk+LsXZxiIR4TF
N3eVIiQXOsEYhjzAUpQ9ZqRj5IIPryyc6dE6WvV6KHVd/S2SjwjCTwpNUZifXSVs
JWZ3ftB25MWJr34kRzImDBVV3j1Rp/wbxcRX0fGCzY5VrbLN1yBV0J16wQPx/RVs
jMIDfk0vCen5e8qYvoZQGjMv4QgYYi6Cc+bVfJnVWIYg1jndQJxgLO2YeYL0FIRU
+WgX/N5h7P+sm72ZpJn9xqFkooBk3rkJXgjmHbRrA0F8tFc6vh7+ZOVtYfFepjNV
BDH74vnOhQXxnWuXHf5aE6BVXUFH0v5cVdk4NKGJkFQsDB0hKkY+vqrMX15A/Ql1
ZRFNhQQ/kX2Now3WJjQemz24e/B2Fph5xAxgb05rhkU+6kG9oFnqcIKXRoJkMqT8
iLhFmx+FXYzNhz/43FAO8ZJr+/Nx24q+ntjzdW56t7xzmlE+0VhYB/1/Q8knuy9f
X4RP9X3iORqNJQ7yHdJ/xWQtqCKzH4uMC1C89OGoT+k9gBohRQlIMmvaz/2e+o3q
quRmSv+JEnoul8gvZ0sNEdGX2Xb3ZnHM+vf9yTW+MCZWelmcOAjyIDYAZ0HR4hek
s93CGdVXGYtbkJOElplyMa/h42TjMXlyCvchFdUWfK3pGnjyhI+r3XkHl3/vvNoq
bTEPw80/1r5RwNr/8uZ+LWOyyQvbzojSX8WpSeqyT9shJd9IF16BXN8ozR1PfEZa
3Qug0hjerlnB7o31grZKPDOobdoLmpZdVEiSvu9z+/10hgKbxkGwgK4d6JfP/mpc
Oy+m/2rmwaHK4SqZCQS8INFUIajYJhy0Ctv82ooHEY4CVl0S0fe3vpF2/tZdFC3i
MVUhIaZipMV9pM/iVSF0cegCRxkTZwmrC+ZOe1XpRkARP0b90L9Cprj7LbkWhkPt
qjTpm97OwpIKLRKesCCAsLHUB9PvsreM3BK+ds8xq+m0teU31upAy8xC4UnyE6CO
stFYAo/JIDuXn/q5EnZ+8Hn4t2ULMr64EAlPk0g0JZhuEosq2HmaxzNbF7T4sMHe
YtH53bAXgkDfplVmiLxU7zUNZwvQa0p/V3wF6qYYNU53LTljLjZn558JtsIzNHAc
NbIl70TuTN8ddk/svK5g9xNyjkiHgdeI6O2yK9RryHRe8Xq/AWFH0csashuyn+sm
bquF6v9iTkpm7k1k43SfjvsXzNawT1xA7hm41Q0QlgyuP5t3UYAdEFdqH1OvxGid
THV93QSiOw3iVm6PFSO/A1Fb7Bz6AvhvOe/WOV+cIUN+heJeSZEAlaH4jAE5sVek
8E2I1G/i2cP8+0Q6FTBefwU6BekMG9DWSRA1NwP79PaKpr8LSw63m2t+4CWMcMrA
64KBKUv7F1O1edEYPheOAeezu9LhDX2X0yLyR0qVALOzGvWYAPWzr6N9rWJ5AsXS
mwY2OPvVlX2AVNrnO9ksiGq/iYWFVrLDAii/8FQbN1044jWgws9cXcb666ICK62z
aNaNCu+kTYHZ9ZTNVu6NZGC4FrwbgnKQKUyah47jEpjfuvmmegbaOtV3/B4McplM
+yNkaE5Bxqg9zdNPyUEKB/fQuAenHp8MPGWPgInkYkw7uKVP31JZpUTlDft2aa9F
0c5oQ66pJ6o7tPYljQhSpmWXhsF4hM9Dy/5j7wIF2mZArkd70u80PmiAf0D1xSQn
T/k0R9HDhkz09GoKY017jLpWeM0sIfPH6mMtAY3OE/nm2RVXgeiU7v6jOVhdWNRL
XlWS8/6nW1LuKGBtP7xy3EcViYvLc7B38KFWarWul6NMi6KYfydJ1CRX/SRkrizo
s3w7CG18wWNo+BmV1YuqF1dlvCYKTZs4qFUvmdYj+C28dKlY3le5W+wxQLli56D4
Fpt0doShBNvu7OdSTql30w5VsUZw9nHevAI7QbXTgoJlX6Ejrg5uSgw+fsyl5g/c
nA0b4/2S7Tb73faj6qzl1hlyHbVe6IBbZRyyr2K02qRN4uKVohnEHrxsDeyRKxPv
2o5WSOvIOw4qJTttrh3KKO2kOVuXecLKTzKBybzQekEwkMJHVHGIrhExEOzNjFEL
Hz/8oiTFyxYr/wE+0VTg/gvzZmPhY0FvXrx5ihjMCET+SMmBifYsXwU/cUQuEZjV
cgDxTFjX3Lzmy8j5+EEt1ZeANXdWwaoqpASHFt1obfj2bd7jsX3MfFhTYcI5e/Gm
b+06tPloHmKpmUjUNOJMNELWua0oJh6iPfQqNdWhIN/y7MpSnGMNlbFEkIwiY/GG
4oMp0wxAPSK7x2P15WevizZaUTSmTdgWLyxMYJLecMgkLhpbx0piosKFV+JBo4em
Cb9udZLTrEfEa+t5Ojxo6ttO5CNMMI/RnW6w18j8HnMMu5xdSmXhH9sk4hzjmL1A
ce2i/+wTPdQoOXzy0JkNOlTwJo5O5lZ9X8msp5M+LOd+2VjotlMpqJowSDSdM0CB
cy2D6GPw/AquHhB9Y0cBPdPT5oOYY2kDkcHXyBNKKKWtT40Lm//Ue3bixk/SwhEH
bTqjfAbNr/o2r2bUUQfqemAwtWHYgbhLvBj7EnSmQxbu2aB+DvTz8oEYfU6Y0jfs
6mOT6fS5W9dHtuxwYcovN4m0/YCNczNSWKXujUKbUbzpQQ2Ql6r2r904viBWFsyE
dO9Umhz9KacU25IU9Qpobe/HoBApHQag1RW78/3Lj9yj8Ghy7hFumMKRUSbczV3w
tKCyTkZ7A7ftRChO8JiJOUVvxnGaeTnyaGmeE1bwld3d4PeHdCgKIO5LDWjImHiS
1V+9YwAT6dzNP82LPh7NNWYPomf+9Jdh9A8DkuNSwOWcH5mZHueV1vnW7OJqSKjI
ZuTf8m0i1aIeLE8lUve7zffuA0SXL+ZWiKkYzpv+/PGooJQ/g0n+5O/mbB/Mg6zv
JmDxjHlb7t48e1d6JXNoucDr3AHuHEzMbCP21X2gnj96Wigud+Hvx+fv3vF3bLdY
lM7iVDpjnP/jaUZLjF0hubYY9/XNOhfVQAb9phrcxDtxzhzfDEeas3b9Mw0eNeTz
G6CkyAAViRFnRRIucyWAMTQy7y+ndCTPUkKacsxD00M3m+hgikFCf9mqKz5m0wO7
huIwFnIg0YaSq5SAROeVUvFlerGl8WWr94znNEh51Qm+DNOHur6iZnVFpXLvYvdF
e2pAPMull6KxJcdBusyeWjVbJw0R023dyCAV6mEq8UxfDXfsaLTyh71tMfHTR7Ay
X3Z2Ee+qtG+XdyXQlwsjkCBDHmJw/S5RziFKB2W1ZChuYvxZgE6oQdHCDZDaQwRd
0EMwD29awz8B2WkgMoKjA4V5Gvp0ztOZN+igXc3xk99ARqr3HarSm2YLdcgssjUB
USSarDd/wZ1QY28+I3joCOsrET73X+CgJ6EVOUW6hHWr2lzacuc1htYcobhbfCem
toOb3CHjdVCpc+Pxc2A7RbZ05RqofJuR4aCJlbasseHA13SDHjfo6AHnLY3K3ZWL
3cK3sRgkslCSoleXJkMoIIGN8qFKAQmy1du1rHBmQAJWvo5Qvut7touWCodTP1Qn
FzJVuRGgN7QZOkhEuMzvTlnGn7n6hWJlEoZJibEUDaToVCPGlsFFoB6sA2x/Yhpt
bFfUvJG7iKiAljyn/bGXW2LeE2/W/hn4qiw71azBwjXvv8kw/JCrSAF+SKcTlzxr
wWLtp1u4M6QWLE9n+Q8bKWyyWbjMpifGN+63USXgjdRXk9Csn3VXfp5KHWTs5og3
SD83+mon4UnwlQSQytrR7eEpPeTGEiYZx115vqW3bT2T952KIEntlfO7eVptL2cA
MXSXqqmDfgp5tFMCpNnHLJ4rAV+5Gv2WYEoVC/G8TRXcFszre6kgONmO0wT6ciAL
ePt8lLNCCuhaz8MJ9zdZxAAJvg1z4Irnhf5siCTNEZYu12/ctWJ9eHBstXtTC/ih
BjhZpaGV+ywSzhQMcugF08vAsHastFoGg+h35OCGVH7NedWtmoPmGs3WXNk/FfIO
7U7JEInXUQOxB2+J8BJFpg/pwP4HP/PGSaY8n6Z64hChQQkdND4ZqKFWv1RZYw8O
UU07ivOgnu1TWH3iYV7+cFuMLgryphYVaWSQwZeCwsMxptng32HQLH0WJDXwHXFk
8H2O89P6lKM77s8zM3EfKjhntofo2DbvFurFdh+BrXb2I7E6MrIFjZcNqGzxcIUI
gbSGHU3+AB+8TDyfWtHAuBQeHQqWpU6Da5GodtIECQok61eQP2Xo3au3vokhn/Yu
rknPjFZGpanX4872a8q0saxnUIEndUBxjxpUcLT9dkDINkVQ1fTNLDOdNAC8tFDQ
VepmMXQOcFVd7RU4YZuwOQqT5PUQAaJC/ZU+V32vdD1gOvLzUfV0oiD92JSSPK4r
WPVqK73Da3WXKOg14yAPw7zKlSQHO+jbMjPJepVKWIwLq69bPgnk9kRkpV9ov7iE
WjmT3SaHxN8QQiVkQ9otyRFvEU2feyqww/jPVRN6Z8BxOisezjd04b/WT+ecppqU
knX6VRRw7mbeqmIGwcxRfkU1GjWmf/PTxvz3uyk/Nslif6jrHQMakpRy2hYnVmIp
3LGqVrqPHq2elrjzpdetUwXp6kNjtUZ5EHlqI685n6prR88jT9DJPcJNAqWZ70A7
BFwHSnvt4mtXBVMDpSY4RStaSNF6+CMSYWaU3u+TbByuYXck3E4DWeFr8pk0TAe7
XXIpd1oa+kIVwuiIJLsfNuRyMQOSQyrZldqZAPpU+4GKJ5oLksFCEHhUOOXFUNZF
AhwrJEznsip1Wb8XRkKIuHn9kt4HDnDZdECxhoYbL5JsXf0eWSGEBemMv137Gq13
20tddvhEHIeH/Om1IFZJx9JP+7XTDAHaVTj0lam48p94QOy9iaWuSjLfADAd7Cm9
9tSAHV4G6bE48NMEDb6E5//xwiYlLoAM+zXyGSElr/6LTwM2C/moXLq9b2UqyDdO
XatfUhTSyH3bIOo47fei48kajsiLPyOJVI/j48R2jWioLT3+0o7e/VbNtQp1dxjt
7JxgvBaB+adNjZxZL4wf/cZuCCSgvoiIpBHUmKxeEMteLr/Z6waxLxkkFwUtFMxN
3ixvNkQDAP643a+U9F2cd8ni9ZosuJXE2PY3RsSM9g3oRGRrHB+2juJQNPlKWsea
WPO+xHx/gKO10RgrR4w6GftiAMVBvTvBDB8WQoDkxIcVSV53MscLs4XA3QLKfbEU
jtTi2lBfEJEhljwOEEuconoI2JUy58Xu9itI5yKIyZvExzEMDcshFAfeT8otyXtz
zy3STHCT1zw/COw9sgWlwSJinO8LDLRtwRXEed6X9aW7q99pGFricWN2mFkgpbog
QigBpKY+Gd0xLig4EMdL7t4Bxz97vtPITO1po/sewbcG2g+wb4lTP5VYnzEEIXIJ
Gp7KVVx2wQqo9rmBOIQIOrzI8zjiK4i7F34ijUfwuMHDaaDbxkOOEMZZf+QBPdr5
xaUF7aZaDsXWvBGQeHPlWyMW51Mqj7H3b+BDU04ZIpznYlF0xAhzeIb+YBLc58N2
dltO5q/jEQpBtfVwpP6EYrNSNBRXVEe+sEJhHaN0bs9zLHekkOKwmENXhp0VrI/i
l4hbw/z9Sl5yJJ77vlsoRy5OTpkOimkcw0+uOfgmBnq4kRHQvjpeTVbV9LKdMLOA
gqqJDW8CKuDFiTsKFUlEBmn+JS9vFhNzOrnNRGEsPs5Snm7g/E+6OSwA3JwnTwdc
G8s37S3OZlc1AJ2o/qU2s8jB+gUiMDiAU6JcQXAtU8LJYU9nTzocXElU31pg3t1u
2GFYwOScllEExTNd1SBaCATOWDWMJy/TsUfHIX5PXnKqWk1Jwe067N7tiEJbOJ29
sb5nzqfH3nUBkPNYxeeaPVJcHR1v3C+STgmMHw2/qyeAwdH4OPKIpNuOR0+Sjoql
j1Col3s3NNuRY2v7azqsCjP0D5ZZt+F2mMJHDYDmB5fFuevsHEuhi0HR/6r+LkYL
umNxf4Ghv5qzBKIGgSw8nvRuW+CMXZb1dsMCMEDs14dshmtFK/OJ1eWuHnh+zqJL
hUYZStQ8VYk/xxU2f1TPGHXQT1MTgtv4548DifyTrvaAwS0EnJWAC9v2LkbRbSvK
fL1ZLDJFE/8rX3Gl2WNU305K9DRYjhEUDI5cyq76OC1RwW3EzQP8U2CqwX2de6ld
LPNIki9mS4gLhJROFsnqxHAsDDUeaF02Wd+no7+4Y0PEdk2FnbGfIbGHzHhXaM27
4bqaOiAEswZ9zWvpQi4iNxpl50EUDG1PSgtgfwiLz9VYpeWaugG/MYVTAfLdAv78
TZjW4jiF9pI+eolh69c+VtVuUi0mPRkr1cnTLHHR+cyEZcLZLr+vAC6XhJUaFQts
aJ2yhAzSa9SOY4vmPzqo9Fr5a53AdNjqTiyIzZNZ3EvGmXoJTBFoiLdeU6TXzLU0
0a3VMINFfrOsjNKkhwFgvO3WVO12/ymzQfMvweyRp9xsTlkGN+TntdE8f3egCKO4
jGV7Lkqb/Pcp9oVLRbECOSPKC48Zmufwy1xtcQIn8lG4siqmFE0WozI1IALQGjob
pq5qPuXt9Wb+U2z6sp9mcGy2Whff84OSkThNGY5tDEqRGwDw2Et83G8MCzNEfhwE
O//UK0c2ySyw5oR0CLgZgOqsGSWP4VS4Yul+98T/SkCMEEPiFFTh4QEGZpYzU/zN
aULVfiLMbOV2HiwxpgZdqpRWRog63RnUb7u5tpT+OEqhSimf+62pfWZ6kr3aw7TH
8BLRHBCEMMbOTkGUi5lLwh+h9bcKXvPebpOPKvbCKuuTozQwJhWoGSuhSe8Tguny
D7nFJ30NzsMvZhBuZVLBHrDuSRMcMIJMPNj/TYeTRqTvrSaq0OP38R/2VMbBEztd
2WWaNMoS84L3hJ22I5fYyQCx3gqwYeuGMYjDuseAoeHBaIoCDtPvMp4k1P9JGcyn
OWlRnUUTl9a5tv7r3xj+eXKi/LXZdVWj5ZBlqi9ZwAMwbE0Rd9u9lbZadANqYc30
4igcHvypt0SGwKzVU8HSFtm/DIIHDvO7tDweU6Tjpd78uoHDiJucu3YiidXQKzjf
AlgNoeLbXSUdyIShPNa710Yj1mRhc8fpdTPEnd1ASRDWCFPQsLLs0Sq71FODuxta
QCaVn/5xioQwGklH0cTUPdraQx+D69kjv44HWGc7HIhXQMLRKkJQ527wgpSKG4iR
oqOXr0/afagY7QiQx0RzK4KJhpdEmlu7PeNsDqFEpmpN4tJbYYJLC3u6TkSbIif0
AP6HQFGYi7Ca8tJL8u02I1Dv+/q1bB/4YYhGcDDJvspLHFT8e7x68hsAK1+sS92H
bj5BakFee8FFwNPT/GPMM77jIMCF1HHoPKxuvM/S/qZ1PGzTNUkqlZuT9w3bW8yu
8xLU30PeTYVDzzNu4vCs+RFE9EZjmouOROizxUp07HxF5HPppQ5VJvo8/FAFKCp5
7UblT7q0agBfS3UNN7n6WBOf7HmbIjair9oGJVSsBzgkW8cYIn7frfsvc/fbJuzx
DQo1YRRbHtCC7+iAgyNUBDErD9TTa5qzJkLhwHIFJdUNEMdLOKqAop1AE7G0ws2t
3+o37Xi2B7TFl5YfKi6//t5hPGet03IPMQqFUY6E8Bm3ArPGRSS4ORM6EiEZtWeG
lcp3v+MqH0ZW31OV03Jj82AhA5nSfPO4gaH/xwSeXv/UqZZ2Fyzcz7TmwudNgKjN
nCnxFPTKvpZeSuWEMWwMiX1Kmo2toV7DUEhAog1V2dax8V6zJk4iIFFAac6+pjaC
MmK/IOZWqFlwMGaeiL+sG3TBSvcrSZXiHFdibqiVsuX9x3I97LTwSkTMOlczi5x5
3+lMLZXRWrxmZ7iY42gfQO/XLgrnkqzLgkdaR5yex9LAqpoLG3/SSObmpBNdZRmk
oBTbgkhroaTXzHrvob4WpIyPs/3RspvmA+1XWbjovzjlG82Ei3Pj7yo/Bv0koiKS
a5srJz03E8fAfmHcCUb+tLfubGn/wM6HFMA/gai/wFhdx40PLgkFe39P3TgX3SNN
BxLbn2wsQ3aVfb/1Gope6GLbODXgIAo76BQkGWLPB3XVPer3XPNKSI6zsPkQwbS2
aj+4zxYuLPTo/K1mPkNeanlZZR2y+vBWN9Uz1fbRu/ofSxRNoCgwhXYTMdz2beQn
Hug8dRcp4IbtB6/POcVZz5elWzRGEm9OfQ0bXJKslSSVYZrad7RF9hfjYH1xgbuX
DhEM2pmyeqPA9YfIPCpQeHsJS3CuzxbGht50F7yK69BeHqS/SVwCwPsbGyN+/MyS
RWq0yhZo7erwjLEdhqxNv1Q1epPvk/vryh++F2UNa8nfCD8Rz28+0CZDaUElXQGD
8q+APPljpjMhROGq9P0UZE8lNf7Nfs7UQNwiO9McgPGyxlsPwRBxzLwnXlrDcahJ
896YY1BEL0Ow4vDLL9C7uND7ohOteitp/XIX8B4eS81srcBOIFWiEHF0rMqk4Z+y
EBkqGVrnfOFVGPv27+SCOMlZyMwHGaI95qG2NTCtte6lWQWX1rTMUTVPClKmh4LS
W/4rrPvQrg6MT2EkiXCk8Z384cDw9hbA4+mDgHWjDBOGhxLh2L7xKX8JdUjc5Lri
cUftxKNqM3eNIpajshh66E9NbkuEP8JkqpzQMTx3/FIRMHy3Q02muTuZHsVxYmwN
1ArERxRTDalVzJnto/3B11+j8xwfwaAYXp3YSodOhLdvYJRaRosthOYDvFB0yzaO
ptMaGRWE8kri9rOpbYmRlCdjQz4JlCUqf1IyDdyZuzmIDf+USLu3x6Z5EZa+Twzh
qkKSijbK6hdTh9PcX904XBG9A/8PxPDlw/Uc38j7qPyBaVtUYYQp61Dwz9ww/INQ
6v15cAMFc9ctlF+f+3tvBZygnuIdNQOJ7z7mnJhn6iKvcabQJxaSdzI7vDWPi9OT
B+4ONfu+Gl1nLIEd73RXLaFR+1+rtHeogGczqoC2V7iGHI5pU4atK/rzxYWZCpi9
GAGbomlZiWr824J49zA39pV8AJsgEiuWCiUM6xX0OC1ZFnSnXrieFZMvqY8C+0le
WHxmw27xhSXfRNWonon2V4jMfLqGV/EPLsgAKGcMQMXmb7admOF57b2gzOpSttmX
Jdkx8y7cgdWinsObcSxSggmxhrX1EWMDT2DGu8pbW3rwVkMdiaVBwVPmh2OhMiPD
TJdM8c4qoLLImZjNcDIYvvbkNtpySIbkVOixdbpGN6Zr5H9XmBrVBDsWMN1zWvlx
h8kWQOVAXRW5bLTNkKcbTf2c5GeCY2EHAi7iPluDYqWpN9LFhruWKDdeUdOmKt/X
gdsYoT2FTL32BkMcrAaSTTgIm2rSbooMhHfqEFGt1qiCnD/KcL3oanjBtIohsTzU
eWcs4kXa3LCTEM0ny+ZUdCwBL1kUeb/q+78K6lwaa3QXhjblGEA7Qraz6Qo8AK3s
e90ywnhUHrFv9lx/xv+zth1mXnnFzTzHvUKARCPIorAmQSJxl/UUkqBlqtxsLusv
RStliZbc8ll0UkfY394s1CEZhRv4E3RMT13xQDnOCQVzGjJhH82L0LvnTRAHl549
8F5VSxG2QrVEPbeNebLvpHnPxSaxS36VnZ+j+CT8ubdb1glLSKgLuNAfJVWuYw8Z
5S0EvXKma+1Yjym0XTVlbqpdG14bK8MVcmggDbc3ZyfBhHUD3M8ta4/XzmWuH7ig
vXrTAZbtoV5jirj77eeBbqBtajkQr0HSXmauTAe2h9BnoUBXTnjr1sVDAC/wdCwj
B7uYPfgnFO6uGoyU/pqBdf5iRzMzIfmkiHm6wHGRe8D9+o6SBGcSazIAjhYLlzEt
mZj50qINs+9nf1PGORudOczFSMrvSmRSC17zJA0tBcsqEKYNhrLv5yV4pcKyoAsD
shRLgLcZxL+Ah7kMmlcPq0aKAO+DGcA6FBPr802iyLNBGj9ita4V1QuvPDad7d4X
iy3XE7tlX6BoYVKYmJoKq4JsSOxYMThAv3BgEpjF8u3RmdpqzOZf5Lw65OrVFjPM
+N3hjrk1Soy19Xta0IoZ+STNiRnwfmqo44kTm8R08Jn4wLqHfh+6uempgS8oAW0E
s24OiPE/1ho5skSiaCr63RuqXA6muB8G49D3af5zYciepPX0L7yXIlxFE4PB9sWx
U5nEgSDvPQvqKSdaLyNNgdFyzF8ZpuO8cLdicIEcg8YJVaEWAxL/nnDgaDHLwIBE
rFCiUBGh823vLp41BK2SaAF0sEG6U5z+31Izso6kQjyRg9Msbbagczqohcc4dfQN
WE3xYOM9yD6i349H8bW1nxq7GSMFpfxAHVXNF/P0ilvyna01TPf8A8/GD/IUa+7o
0AICDyCCWL33tp6DOwcQTBwitQUDFZT8lknDCzp18Rxfqsur1cZZMZsQ872/V8HS
pkzLSXZCiB7FUstPEvOR9Hn3cgfb2yrcKyyxRLiIHf41jQPOg7cDj8GgdtuzoaL3
W3aFXT/Qg1ywcTkB4KQoGY5p3IBQUaVlIsSXOp4q35s/o/2KFBup+NabbPP8FqX9
Zt9SrVXFkABbZe9OfF5gykquiBsoP/7BoTK5dLz0YIk8VIipQs7Ruk5SeWbG6J6h
WpoSZN9u335sFokrs0P5MtcOrtMWBBXPyUSvnEy4FSbOPmmXDn9880tzn3b1BVJR
AzuD2JS4eyr6688aYAFhXOI5rVsYUzHtSeZp/4175nT0NNq+VdtZQRKJ/V9ybc4d
3FvPIssIK3K+9xXAdtTnziddECO1LbjfqoQjcWdRVq8d2jF/0aKR6vXpUPTtTx+w
6zSCR1uFfScWbR93AUaYOczCCNG/bU7lDMM6PHnavfq2ONlH6rgc222OKHw9z+No
bPgI075q9H89hG99uc/3MrsXGLm5RjUKnHS85eKLzyRMgK17o5TE/x7MZ/6SLivd
vNytfed/Z8ofyKF8SDqqcEM2vRxDDag2T+feqXRcCfZLFrQBq+Tpw2huS+F9fBap
2el5I35adMNlxLw1hNMuFOf7w4SenJyvnVEB0j+YtHVJ3RGiYY/dVtWpWjWnKpbQ
IML4mXoYQu7KLedKnbq58VfvH+IE1w27MgjzCcSJRx9Ig1PUnMLvyOHah/3mK5Ns
lCyG59nsXyQSV4iEk27vTpQm3qOIkCEPt0RJigUj7vzIIsqEsUcg41aXp7fh8CGv
d27gXgjMVa2tQGAJe9jcwLNDeqVI/yFIY0O8eSbAxtmy3AxBb5BsisiEKtca0RYJ
AdjHhWjsRIoLZNDmMPc8f5ZU4A0AMLY0ZT0VZ0z+V6D/qiuKHGAb95GHe/oBLXOU
wiJYnVq/w1TghG/jtNHAjlDooMLEZ62PbZkdfgpcgdO5JPQerWmVqUcLq4vezJFT
3LVsCRSClIHZSdmJ7yqXew76mBl3hyxrH7If06uQyoOlaHo7kWQNO450jFen8eZQ
5UBnOajptArlDP/Y4//PTT7PUA/2ekBR35V1p8O/ieohwZ7QYAbhRZOr8pOZJGjT
hZ95QtRUDzXF/U8n5AQ9X+IOceCc5hA9ET+af83Y3ajuMU9J/A4oYVxEWmRXFTZH
QaqByyHDBvQMxPYDNZ9liOyylLnIua2bml4u5d6R9+UMzPGn+RM/ZMd5UwjnZcaP
XJ5d88bqN8yGa7i5OyeH7TV0m0xxEsupmFxTcW334bTmDEIvo7wJJY8kT4cxVbi2
9IL0gRQLV1jGiv16uvhrRBTOFr7vXr5nKCmEyJ7S1VWPNgu4QFDWabsAJ3pgTegU
gwi6Ji1txpeTzKYyZrpr2kW7CQIADLASldcvWrhUHJFF6ISEn8N++xSKQCS+RFM+
MY8QCdiy70S47Rkn4rlPdneDGcB2/Eh736qklu3cAFtMvYpEnR677OGdd65nlkuO
J3Mrv8tO/rDtkM0D8NDcPwGw0YkkhPdiUmdRgd+/hFgmhy2IJBkJ+6N++Nm3x3R4
0LwWpcTu1j3d5UQHygqaA+2P5o1LbmhinDGqO841Ej61njODCMPY7rNG9yBKICnv
w5HBHsIyUStgPeUjIp0fGSR0Y53ZXr3a2Z+gj0O9tqXsRHtgn3pDuQJiJAvp7sn2
K8MsFI4vlk5smLikJ8Y+WoOe7TU7oFvlPsDDwcfDcLSdKhIpG77BGCiha3XJkixT
wVKp6TG6BffLXAsLlYcuKWAonwxwvLMwFc+bz1RS4DUeivpiwXssciBb91Jmrwek
QlvTPx/9gUcQLknGjVQciE+W9isn0+wxrEQadi56vvB1eIhCn3IojMpMzrhCR9GA
rFFi6OlpMiQGg1eqCnSriANUcoC/t3uCeTewdXdM0ITcwkzjFB0bkkjAjYoFh0zZ
iYkAb9n4ofyGtmUHp9BmPSC8yOkFldAul1kBHF/+i13PPWe0w9ubUF+QFu48YLzF
QS2OdQnVkq3hbmRjx3q9cGOHtWDm6q1FcPd/IcJwi92HFAisdrYAEYijFrjA8Yu4
fnP9Xssewqc9x4yHBLmMf8JAMOnElZJXmJIcBPTFUX0w6bX1IuwZ8C8blmm39F9+
abeIvmjO3944sf9xohNI8mC/2Wm5aFp10QGLCjUJXsQkaH0VwTO2ZjFA1PwlktlL
GE3/ddQM/QK8dLgfIShmuHvpYFj5pc7WkyziK6dBTmfFmvVPGw4R8waowfgACEcE
MbQTKLZX3EHinBNfaszsBfIDsVIdqbQoYb5GHMwCz7Nzpk+ChcurYJg++muPj0mK
3jc3SNLcvjZVQtM4MI4Hgp13QwVuKQzP2MMdbXYG7vhT6VHLAWiR9OVL8NfEXHql
191dTr97Qb4ZbgHe9o8H2vB4WAH4F6VeQje7pE38clY1BPY6ivEIPEfxT6xicgT7
Bb1c4y2OecEJu4SPW7HJhJq6EBuUv3uuzta3nKBOVDXxYlsrhvl2Qk16fe3cqsuv
kc4ZGd6GGqPRC+vIiaobFvreTYiyY/Cae9DhKOEJa/n88oJRdvZDJL3wNaDUYq3h
vyQrm4kpL1vFNg5aviTuhiOsL9WBeLKQ0dfX/a4irjSPWFEupRBUyNFu0hZMupgP
W668BTTBLyYcJPf7OGI4zCTgYmcXK7aE8REX7nriEr18Ah1xdA6IqaSwm98E3p8V
gOcCnYWlONGIluyknuZNJ8+m2302SncSVXMInOkwFIFaJZpNn/rZOvOWmYzlJUAg
KreyiWqOvA2HgvtvmDWzI7lIalC6uVxZiyMIBoDO8Bha3Mj3oSqjzaV/OV0rsZT3
2/Osth7v3a5iJD03Ich/gn/40H1pBpQ3V0u4xZcKHQc46DcFgQ5/MGbrdI+mFH30
9ZFskg3dV8ZLAoBMPjONURvqdHjvoozvgUV/8xmhIJrycBlXs7hxw8D9GMLH328V
TVdwWIQ9vELXx8VT48tiTdqsgi8gKCPAY2cnDa28PP94zFMcL8v/il6it3zgMSw0
6nVAf3rEcAuh+tQFdLEcB7WzTZwWKApZOKoJNz6V7d70pNqqj9+qXM3JwFrduA/C
ci1vgR8oyp3Rwb+3byyN9Cs8K4roRklddKQvUEBBsQxiIlnXBjthiiucmYjWPFMJ
B3NEa62M6fdWeYUL8Nz6qyvkP/1PtKlNFj72MTEifnKvJ7oP5Hy9eUKISBgaCeDA
jXRRnXOnAmhgD4FXPG9RDsi/HlvRgOveAICFslN9qqKGNrwBX1BP/30AliqGS4LE
05g0uFbCGncyyjE4gPfTTpDmzQqIQfAJYrnCG0D4lntYEigeZhbMpMf8lORfZQTs
ciIjDqbaxIsZq28nlQCWFK5IDBQvlrxJhb+M9B22bdy0OaipwgzFVTH1u2rA6G8w
`pragma protect end_protected
