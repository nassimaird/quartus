// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KtLDd0OdtXcUEK2iEiAOEP0bm8jbE/VU3XtCOgoYFqmTr6XltxkKqsgoOb9jZ8xCU642WjCROKbw
R2vKC73hn0l1PgSxOkTESamAS5mGpdjnXneokqUx9Ky4RYZKofuRpfnmnzJRGPSDVVVPI6R3BwTl
Y3uALNOYLwxclHlmI6yP6Ji30khyfgoWbtaIMIiqoXxKKMO/ssDLCntd2pp0MUSVJEpsfcnywib9
7UVnN/M7I74eAYQxZ2eDidXyC7Wc2/GLheC7CD2wuP4JN/S7HU/QO1BOMhpEq2mJcuH9AkmGL6LO
31UrsLNkycltWs4XOH78SzqQA/Bi2LYefJLOIA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2160)
Fuq72wZv5hrQc9thwFEuxXiixLSIfrdLhlDOcXPVvc0w1J2fkyrGHqlU8hOxUlTxOjg3ug8Qu9qN
bYOoFmVIb0PyBeZque2fMSYd1OCSkr6HbD2hLCWjZZt+b4zohkRkoNCRcDlRcCeirgKZzru+bvF/
7D/JKUDZGGyGvnhdXNWQ3GEIVOyRWRWqZiWxDAZVjonl8EJV7Oco4za5MMygzt+vh6A/RlvtmSNH
foLZaRu2fVzGzXOfZzbRe58dKb8lkRAawhbJwKDgvNLb/r8otnriR3P0o0jkIU9EtZyY8r8HTouY
W8pbsajvIojV11EZQ9WgDBpoJ7vNjjxHWXxk+IFfyKIPf3VVSAEZdqHafwxSafRUaGHuK0F0uv0v
SrN13utAovPaXEF/N1bO3SnOTZp7BDDKv+IxqNCZPc/UaKvy6F1eBTA9ulWLJFchblTDwQIj+MQo
YyhExTVjQqKuyJlHC4cQqNzVQws5T5uoEK8WZ5OxnQwCUBUss1r7Md6enrxaZ8wwxlONGlHZ4gdq
ITvrj9s3jJPDUZkwRGnovP49g6NZwub9I030owueVcp7hNXRfrxCuNsV+IlFtPJgyH6QB/y3ZpZL
9dPqXzXucpYZg8rSBzD16OyV4ZH6zzXswaGgjLklqRtgS+j6S9c4NMaCRawkOIA8+no8o09Qe31N
3XVD2I0YqhtKva6LF4yS0CGiyaJBJnUuwZVFdYoYG4q9GinJ/8USlk1/DFm7V90yKlOUfELuxT8A
bIahmrszsjwfU+ns5Ol9MpZnCQApraJplGarntxQ7g3GTYURqCs/0ww7T4/Sp77cgYUnpHWFUWx5
fE0bVVe+aKjnL/cIizqiN3ZTEmRH5aeF48XxlK52RwzTM92PKjGiWzdknlqCZ6tuhCqxh9h6eb4l
vFe2tHVGQQE5mx7Ve2OekUjCEnTzLXd0R+vJIH4HgVwdGkuG1MgCP9I5wPaST0YT38hsEEhieSlE
rgnfV//5RwR3DOIAMJ330zRXz3NXIr5T0cvfOfNUVQvSxkev42G+DKHwjmgnIzf1ZG6Fmd0jlZUE
MnaZmJLJJPkdj1sVv04xfI3zNypFFy2mEwdNwWU31+AhXJVHtGXuZ+uXeJmooTlu9Cn32gk4boRh
f/2k1YBqg0XtiydjFgehGUZE5ckXa0E375gga1MpjmeAN5ws6hnZjqMtYKG78POvq42BWTUtJL+a
fGmVZl93ApvxewS3SdKOGeFTytbdXWU1FO39mF7j2YbmGz5AEyhPpapKWP11S4ewTTs9fTBS69EI
ATaQZtn4Pl/0EfwV1Zw//IMEWxCqRJ8nDosZZAzf4k4MQu9Z2t9SdE3HJiXPxLWLqwNXx+6soO/w
Q7MfqzYf4wNMlVQD9GJ2xMnEeCCnxvHQNAmF2dGKDdhR6S/piLsb2jjo09iTWIBo97g4m/TxlEEp
3MftfC5eBkn49h+BZGuMT4dz/Xngy17MLvOJ95q34mG/R+9n7t7wedMsNK6+ZVTUOCU8XEap2T4C
egfM2gOGW+GYmggKTBSqW3WW4B50Lq7+mWtg9NxMwZjFWpLSNkJlTKOVTrlbVTyMp8zvyXrIXrfj
mXvPGiCsDPv5ijVFMDz+v2yZ/vFCANX4UkMpMLULsHAxl2e6pz1x85dVKSefDPpxZvH+uiV+GenO
NTML/0aeaa6vX/8UJ6wiVVEAV33xaOOxCTtYwjd08lqIBnbObi2sSNkzFS+cKZ61V3Bp0AN7ELgN
5I79VZqgA/VO6dkbCQj9QY0tPG5GleWj8yhDR/6ILfYOnxR8E8CYiRc/tou6rvo7wMeEiFgXY92D
qjb0+fxg9HEXrNTXhQIMfYOY4KJQarob5dQD1bzmEInZZcJZPQzraJlu7GgjjFY09Q/soCnHEzsV
vtngCHI+bUt0yiASZVfZRXSrmkgmfds5FL2fJeenNLetLSDf79EZrdOGX5JbAJjFhzvF8Qki2Rr4
kLAAQd3eQTzzla0Eh/SrG/I8ldc7jQ6VYDGlW5RTFKSo/12GO3uFWisxk3UMxunIez5IiiTg30xT
xo3fBdYAxG5L9t4iQrFxtG5mgoZe9D1KIXcVAOyp9JvG5b1nDsop8GtKHeYd1+nu3xjao9olzDjW
hhqIrvgJAQrNWS/4ypIqrFMz7Dv0kujjg3+kk9rXqpiDjaTC9oT8vgJnc8KpOIinaYeCt8MEUH0n
YKp2n9mHLcccpiiH6uBjpoE9dGorTvrfKSgs/hYon0DFwKdP3OvNVVHfK8aHIFDqOYAT4xOrAGAr
DjO0J4JPzqxeHwsyE6vvY1xf/chdOS3T7nfotfUZJtlL1REc9DQSTf+qZm36V2v5fTB6F3PJwirJ
PgYzo3uT9Mbz5TltXf+Z9EVPN1g88kp96vBATAijmUzCjVpfdnLTjqL/HKn+C03PCZINU4js6wsm
NQyFGtSgj6i6bLJUM6eMVMKj3nP7jUUEM1IuebmUyjc3WIn4ZhzVSjfj4v8CiZDbnLzsIs0x5C1/
k7U7mAFcRs2ShWKHU0CEOK5tTs/m9NkcpPNFdHNMvgce7adj0EnooymOmH3I4PsCnq+Bw7tEKeu1
GNS1NFkxC/obMAtAcwzhv09xz7Ia3kRUJ3qWfcWw/JGJ1HGWxQs5j0yCtevmZH5MNgyOcKQzM0N7
Kfxyw0eEAigzMnTppHsP9/hlgTIMcgrUer+fBVHhLvqmXoXBIx/gg+/cdC8zDGqw4zqpFm+x2Roe
mH6oviSar0eH4CX5wGrAWH/u//mHjOpH3d4XkkCF8VbA27zGVwVySY6uK88W5k3dtK84w7Z9FVPf
oZ+hCYQ3wEvkH+Y4q6SEs8NkTaqVHHK+Sb722wl+UL+3wOiosIh12w4VMBBxraz7/A5v
`pragma protect end_protected
