`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aH5SH09pvqe7ZJTVPAHrr7jlgOIm8eJ8mNzH2YBkyqC2UGfYOSPj8Haxpqs12AGc
o3NfNt2mCfObXzYVW057/3+t2g2AstCsx/QVDZwV80ZMmxIPXrhV5kwHCbX+GeV0
Y6pn2kwyKFAlW9Bm7bFW4cXZKxWZ2yYK9tEnNeCcPMM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
ka3dSRYcrs3vIOWqD9cikIKqZ5zglMX1KwuVdN2QLv99oAMFmFrkQ9TmRFmKNr1i
BD89X9YUEKLFkTlMQ3rRYrNHCG4njcwKZVoS1EmtDRhLOCJUCdCtdI8J3DVeO6mB
D89oWxXfMJj0Zg3GKYKV+IMA7conB9BRW3sMwoIc9OP3HiNisGavab3Ona9gRjju
po2AZmfDyqoeVLptNeKYca65Cbn6kL/Z6ipy2h9ZQI0qawW06pADLJ+Nr8AdP/5v
s87hvMWnkABs1JMWBywwAKAdrkiHpvPspuDAXcA2ARh70f38mt5jzeiUv6ToLRWB
R6yPjy6L8uPXLUX/9Wp5Hi9bQNtw/0VxTGZjr9Q4GUmy2qiAwSZ4s43Ik8O4OY8k
0lwwKFQiqTD4WPyrMZ+2hLm8klmxeyOnP+K6DobsQiDI0IHSGFN6/3M7fbkACX9Q
tPEr64wGngntpeE7PnlRcmTVvypOtECy8zBQqEKxad1yTkYks/8y085aSjRBhwsO
4j48rFJexi/QZjn7H4pHT0lFNhjCizC/zhKLuprnRhO8UR2ZQEAfJ3VR7WMXBLZa
PxIbx8MzRm0Nb/pWkdYVb2v7Aq2+HQBItE94DjBkOBwsLmuO9iDazWisPRKXBK3K
ZgHUvt5PpgB1Jv5QJoHr+dCBjJiDE6tibF5fQ6eSqmvd5DJHnrJGwyKZ7HhSzF65
8F7qcICR1gkqvefKjmRFxdO3mCdlGWxWxcZFd8/oYd+5mBMQFhPppyvyYTYufeWu
xpOiJOEsY/q+7iaRnzHRj2U7agcI61Lj+XStWASsevBVlxM1Zfah1KpMZSc4lo72
wUQvKmlaQr8orsqtrr9DxL2ypHlJDJHHhqWRsPPsoDT1HjlL5lQzeaDh+h6bFFPJ
UOk4x5WiDSTzJOSy89WiXrIJ8ORxtPH/zZ41muJLDp79l/r5ogtNSvJegzheSDN/
ENfZB80LQlexPh4qeI1wrY7/PesX3UdRHkAQvCQFXp+dnjsnLsM+zQThd+mz2Zwa
XFlpgdbOD4w/hVMvl5DyQ0vQs3c/MxZTEfQfpBbggE6DMDVLqzCKv3bnAOtX8Mnb
QROpUL/YfKv0atTwwRr9cse7UxwH8m9fk61JtxVEjbIsvNmys1RpUl+uWGY+C3ZJ
HHr8+5/KGes4aiW0VV5Eav/oDEKpTTcTHR3V9hS8BQYIKWvn/SxABCVYO05MEHmA
75rxfoVWD65Xl3S8suA9DbfcM/Y+NxN6kwNOYY3TbrNINXOAF4Ue/7vz67cC5BEE
bWYdDVT8cnw/Ugu7OzjprqYA971t2BLXctN4p7LnZcHPSMf9YPuwXlnfoAWenxbP
01A9S6fIzaE3NKbYzqcqhOmIIfhtydSmFRPBON4/7qYc5uq9viPXwClnE4MwuXRo
DO+HF1ABmeZxVCtgNaYwwT5pcXuVQj9z1laR+wo8vsG4clmTufPALt5TWbDESmiq
2im+7i5q9YLER5A+QBAR4l6jq2RyrSQvcUBTW4Xphra1kl0Nv7X8epbIISfCtp/H
ctZPyl2PzXOAiGFIRR1DJ83TnLSiMIgmXdjAwJ0vOecGQdHHk8UrSDgnTMLc5t3x
5RWzPrM4glEx4e+sErwG4SIGwsoS76AsUeFIfENVCD0sAS+etrJnvDFRhTT8gatK
8NN+tcKCICzwSX4OegpuyjcCIf29lQG+46PpK0jgLe+ik/KkJKT04En9GPDWBwGG
ELKaPIaLg9vB1Rb2gtHY1TWxFcoNOk8FF81hKDlnT3F9gw1SWXlogD3Pwq1WQaxJ
ZvpYxY1nJY/W51Z1iBM6TCR+q+oXcesMJkRDLYF18KJpxdq2xgIWmAyHLCrlvayk
Mg3HaUZ8D3WGF5OcHoh8tTrtV70K0SY64TX0gN5Mx/8OWFNe1TkJV6gLxzvej8Vd
8xaLOzd8wIuYv1pCc7eUmbrX7oVHxb9DhEJYkcN5JeBCH7zBKVxEktU1Z+sBsLQU
bJE7iE6xQQBL5uYEuss0hVWv76Obg8600slTfHvBbiEGHDE45vBl5s6IKgWEi1FP
mPxEUCzJnsv5Jo01f8VaBMjZrp4aswU8//xxGNTwYx3PUH+F3448RHcF1KbEN4fu
4jEev+90otuN+VLqD0b1HYqILRoMG2oVwUlF+tIAbkQcRGcLDYWHd+uzT9LaGXgm
sm0KKTpRrWS16W0/IKiC+D9jUUUM+1MGv10Xmpd6f0GR7SnKJzMov/xXfTPsgpOq
0HzJ4LmOuQP+WQVILl7yewUMWYWGLFcwHs/ivACx7XVN2bFSkvH7NlzrI7DCRwX2
B2yloCNItGQGcEeKxGC9kp429g6BkwtVXYUd6qxi1aiLOgUzfT9PI3uWqrAacgGI
Kk3Xove+vOVM+wyaoybmlds0bW4L/HWwaAohP3lQhm5mwxl3LpqxOqsDpfs8lATg
WxOAb73pvhv5hW/8QU3OEVumulQyTg1tChwlHAoau8ZgbuErXC0nfW9SHqehOaMc
Rt6CaKR7ksBENbzzYyvSBIg+9zLWfQiGXKstt5v22OtQlQnC2SvgLb9GXSVC4XQS
G3uUXk7GR2xxH3NihhvTPIfR09KtzFjfWqjZmeIavYmpQu64OIqGNGd9fT9ZBfbB
C2IuEO/VPdKLXfSSm5dug5Ht72UaCvmJmeTtGvCnNwL8T3LVbpEeaAbUznmsB9Vm
Rt8zLy/wKpOAupp6Z211sOdlEbSxN4VJe74iYSaaS1Zq1mP5Nxc3bUaGL3rmHjQX
MbVVR7a0nd2JJQG/wUp30Val56GK0isNDSYUv/xYZwb7veKH/1NunfqdqqTs3//F
DXKEIXhmwbO7pl6J6Z+jjxU4amNOIpz6Dbq4Riqsuq7Ft7lxF2KLM2uVoNkVJJE5
PVoMcECQL57r/zqG6hfKJUcSu5fyB2Lx/cwqe3W+ntQ+p/Jkfs5S7sBlFenU6A37
/vonouYlrwL6997dsb/mzZeAkrewbqICDVrVPUw7K29+mwxsRuMnDQtOo+jlHOs4
taD/isg0xuSC2kT4WfGIvBS9MaKq43ovOG7THw5mWJV85W1C2s/sctebVlZYPGi1
sEPwuqGiUXUrSgIef5qr/ZTEGfZEqxOLFds9NQnkvLGSTJ4nKZPfPZ8PcKkzkOa6
H9AcPsdkLkxJeHznlv21CLC8g1uQM/6ty26js82jhoPkJ0ye3Wudr4vyFQ8TkFQP
nGh77hLNMLO9n4emRXtVB1ZitvAUWgcao+1qtcW0JKDSGiRUtlpnOKrlzBvwSDMR
0yCtVQRW62PhdXJctqqQoqwaPR9oqO7fEL0mrHVdKIU30qOhSV/N6bri1FFFi5pM
0UmxA7vPA2GYP9jGXSa9Ih3PwY2LRLH5fUguMYhh9LknON/8uFs4xSPZsdV2d+xQ
lY0WQ5vVvd2da9XJyORyRdc3tvh1IviS9T/1DswrZP6Q3NwrRAwGX/nM+Op7AET6
R/G6ujARsdVoPh7RvvWDVjapD/BcgF3JaS1IR14lWgN0cbqcTQxQ1G7VD5Y7OGnL
WhEFLALE3Kbw6/nielrFMudY2NsmE8I8FT9ALFYsNx9iiNOROnMR0x8yeOXkGcS6
LsnRPxBIW35Smok4zOCCi29AIBfTyjSusOGUL6Qs0cSh8XaskUhpTOsXAbgjxQ1R
ojdPQD2JpnSRXWsX4GngbUQF2pDbpUzUX+5oGXdys8sFLNJai3nPK4im3vm9n0fc
+oo9s/1uT1Gy4t/kmmDqY9ZbkQ5R9MDhDnXF+qh47Oay6NAGjWj9AQrBwiuXY9P5
E6g+R5QS9BEnvYxVWOeMgOWUEVuCExsckWNx3SLY/b2mSaFmEw8hxIJVLhJdjjai
8OWgCM8Fi8oKXKUC2EKDAKwZjAf9A0ZRqVl8NbLPuCdfff5pBPKr83NZsSeXXLu2
MWa6AOhkUzCOZlLNegLqcPleFcJZKP1KpP6EuciOvUtpCeqYmaXaFvyyH1ImEHyK
XaUuga9Hp5pao1RMn/G8OFihZbDzG0Vzsim9g8NJ1x9gGW3UaKzyWHOreW9abGcK
NHJnBrBzYpBpmTloDP6IoZ2BIj3wTqZ6Z2jd3ilS31pJaLmkTndZy80rdWgokyDf
W4lee7WhSdXvgXV0AD2nqujH/iqYiw0ElhIZpgRrQtCoOdv6WKmSp+y0upUV1r4C
OHrElwSai3axyulbMAozHHSt6vpw0FsWucAo8n3qTHWf2j25ctMKBOj/sbkBHyyU
R+uoHdlRqMA6s0XaTuCy3zAt5HRPtrbzZt8oCkcKFkWF82rZ9rXEpLVzw2ra1uaX
826bggryXDFlwdHXQZXcHb6/0OQitYP/NJZK/7T+YEBP9HOcW0ejWqDBVTWgt8N8
TAMPjN70qlfkOFuwJX1njiodLTcXlSVKXjNgqEPOazY4I7eWmz9bEUwj7K5hWzh6
9AJJil23Utu16o3XtoZ4eRLU1zvIyQoK03CT62g7xl2fhhyIb61skWMslvvVozOI
X27RjM363eXn0OnSTKX4c2cNHPOhTTJOuqzT2GSNKScL4PBKP39thdCehLhJy7rP
+hWVFCpMIPapbJXwawnimF78JzIcf+jXtvP56kN3nhcX4nVAaw5pahdFAHbyevS+
xyUvJKJ3pSoyMqVSRIJdxYLDbZuQ6TjzQe9R4T+js8obmjjm3BUY8dCqnlTpv7g3
P5Syhbw/13cP1KXjQLD4bgAYD5TemGVw1/0ddVSZwa88IJkuCEcGe82pp549Hl4W
+lRCxyeUNRMcAPlRvucRFdWKfr2WBIHK7+1nXZOX68aQ48KM80+7EFIrVf+C6ymq
rikWYFEvicb37ANPy3T5RDfbpILkycsznG34BLaP7tjsi/E+sZQtXUpKLNMr2jGd
DFisYsn7NXmPZKV+RBEVKnMaY8yqLPGCxad2qD0VEkqeBXN3rAy+99vBPacHwP6v
uJXzuhDTRtG55yp9yuhbOPNZyCW5UZsf5dHR0P+x8sKqozWAR4OGVTu6ciPGabzi
vjQr22ERab8FcxDuXC94keSc0Lg+v+s6fGlhOV4O8V3t3DPJdRgAOeSh9bwymcTY
/JVHPogC6cHQq4OrN8W/srlGNdTlD1Q71K2ztN1OyU2F6sLGo4hZm6jdAA8wjBsp
AfRDJiCbySnH5qiFchTGQvUBVwxyFLoBJS0aVaRd1Ylj38+6YYWQsgppSF5HjTI9
NZ0qBJFV8t7rf5MKF7FFVHRjrk67kUSHWrrEoGHztLMwjeV6h46ecHPXmONTGANY
af+1qA9EzbN9G+/aQz8p1EshtMgBPjJ794BDzGhR8ILkPBYM6+bJ6Hrk2MzwC9CK
aL/vk7tK0zNadlvKChlr7PnvfW+k7FQGZT+EAKzmIcZNhoMmzpyZoyR87htx8d+K
HNA24ICtx0DMbtzC4iVJIf8q1C0lx4291RQVyKxy37bL0gybV2bKI0U9qLZcnrjN
CNLEzW3k1ezru+6THFcGkTy97TTtJelvxspzq2kypxtEzVS3RsvRrGNDIj1xEZ1y
nL4CYWau5FJPWxPkd6vzI0z6/iAQvFR8mUy6l30PmTooaKAsYVEVccqGtXEVxLkd
khnbxqvdliEDAMBnGdNcQLCmfKTfpDw1RZ42w4ra6burLIHbq0+NXy+H1TQ+ux9V
BT2Lm0R1yaH5khqwyTWHwkVSrjvh0Wey6XDPGfQenKbDG1wDEOcz68gJTu7gqltN
dP3cdBwQoSyLi1718s122eSP8Rz/STVrpAEoQ5xbbbBzKE4qqSLUXTkil6KUQFZb
px7/rvK3SMrLvuUoTjLUR309hxeMITC+bb5JUlYnPbZuEOBrAiE/gHNgvB33UHvA
SZZNxw4WpX1AzzNeP9H3JE4/HiQF28m2oX8j5q8MHmfTN/denndgLGkFW/MHV0Jm
UOMXcNiS76hEevVrqDzO27+GymKAk7I0bVNfr+0zX0g4cWF9QbPgAiYluAh9SybP
9vdJVrBvbyrsX/ZWR0hvC6FZjLcokLX7jKfrykt5lZR7A7IOfWzjovUeKIBxPRkc
A5linLHt/AEmZ2L/OGA9IVobM+isVNsYEdZ3G6yHQTQ4Nr4UBNPIDkw671j1UP0r
efadiN0jsP+/C4tXvpdZdT6NJjL8r79oXsreO1x4KD6xQXcmBIn7XtH8tnESOR5B
ok7wON0Me1dWwbcV2auGiOhbQrFmDtLYlduNSaRYi0tbNianw4jZd9Z/xOOzm+Qh
yQHGL+SqlKWgLRi95jlVWk7gLfpne0sUL9cVaZCysoJyfK6Cx3vA4v+r9iwBJNIG
G2UjhFQN/bIOYFB+KQO161jVEP6oyTmP/DrWywK3Sb18E35ILa/aqsKhKLHI1xiL
zhl49UEUtMWE6IboHkypR+LEJRf7fCZzid0uEdp81rRh4mSRfG03dyQdOn2qK/NX
El0/u4v8wbaSVdty8aIwRnAEF+GInmFdojFIYCxz806wMTEoaSrSc9qntIOYzCeZ
Zx5xLjCmsL6ImyOpIasppM3huw/UZ7n2JbeM40N8gsIDdXDzFvmaxs+LWP7QflsL
HfI3L9+WXr3VkgUSeXQIhr4eNa0eYRDCtV7uQfopevYNhN7lkY4kYm0QF1DSgyVW
NtNf1auSnxmXAg5MmsyS9HB0Q5mCnhQq71PG1JwUBrUbiuBbMVPxa3GSGan8ttE7
tVeELhI2NEAXd6QMib1OVPLWpJM1nm6dXPi5PDzuG92iBETpnpNztiUwVK6mW6hu
l1J6sXi2ewNKlGQvVsPJgN9qXyILa0fD+tnHEUqbjTzn87fZQ75rjPVLK2s6E6Tn
Bjoco4aYWR3VDAEjIlJ81HTmP8Za9il/58LH9CYBUYsxcWT5tu5LEp6V6CiKgcYM
MH9sH5PGsnbtvtjFEYoq4dR+cwkuMT3zND8fnh15MskSzF0Th2lYzl3dxY5Qvv2+
HajZpoQv33nYCOz/yLw2v4KqBR97ryoE34Agpu3ELTKJ7Ujmogv2lOaFdwteh2aV
26ejesczZjRfIx7wyVO/mIa97hbOX7NX0csjoktNT/PHsxyc/t2mMSCuWc8agdHU
EcbxNfCtEd8f/RcO+1Onlq3i7xM8xhWtvX3acRxmvybuMPDVi5hpK88nemwVb1Tk
XPFqQB9se3L+tCgoyLYQjXOYiQCkF8ix8rl4Akv/ZqlWTGN0xaZawQt+o6Hnc72z
ENu2fd1BwIeDx5D8Nk29xnGzdCl699dAu4t2P787/rGI4NujLyqIVaIQBdei+aMK
6JIEZ8oZWUt7PWl2mXpLFpN3+aABuL0Y+ktc3xSS7Uwl27im4g28M7ib6GN9MQXE
4OGcSJ5SVCc9np7OINpYAxwHF5cHWlCX3uC6y/nuyD5iKWfSdMqHs7ypuANH4FJp
Wci16nLA8agn6cgKq3Kw3VBVVxLtjj7+Vj2s6aRIBSxo5vAZzM9O8ACOXL/3i//O
h1Z1BAm46CWas2yNu4n7015ojPZxJgp+WTsF1Q/ZGdnJWA3z27A7fmqkEBocY2k4
y08nU44iG+J10ta7ySnLmQ==
`pragma protect end_protected
