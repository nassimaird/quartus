��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K��R�9��Y�%�itCy�k"l|�.���n�g�����P���y2fy�9���!��NUr�u��ֈ�Ê�k��!�b���sI��+��4����olb�Cǘ����3����Z-km��('�/Έ����H�����߫��[+�|
P�����D�m�@橷���>>[V���^��S�(-����(?m�:r���azBꇐ|���S�;����J����)���e(
|�3V��]�=CG)X1pZ�":&�~��
�L2�mB�V�c�A�В����&��χ�pYFx��*���ȫ�%����t�p�AVo	G�I6ȗ�Y��&�Q��Zf"���%W�������� x��K����4s����+5��"��q�#�JG�s�zVj���
��R�vj��&.xz-�+Qѷ��v���Y��$�����;^;�#k^\�Zm��c?�QY�����7��nd����N2c��n4�C،@�PP�*;츰zGD��{�����fQ��F�|�ϧJ�J��F��_�Է���o�t�;j��@R�n4*C{��y��tY�x�#�Ԑ�r�$�-�AM����\`R�⩛�ĈjjukEݛ&������ET�/�\&���e,VA&^pa���S�و� �+�[/Z�Z���!o��.D?��R?�sM��W-b��'���6��d��e�T���3�p��
�o�u�9��������ԣP�>�V� b*�v.,صR�g���g#]�Z��n�����ʎ򆤔�k]�L�I%�P��)3}Z~���ǧ7Q1���͡i�`5\Exdur��BP����cM僴��QOfY�9Z�sɓ�ݚ�I��5�>� A���);���gg��.~9���8���f6�M���i�o4D>\��ԘK���m��Esnb�z)�Kc 0\�]�<�w���Dv-��f�vF�36�����`�oZ�E����L���`L���1Z�ĭ�e�uǰ�C{�|;�)5^3اN�h�(�W����K�u��GJ���u>m]7������6�#�?��,�&�o�"cc�����ƅcG(@7�`�%�g�a%Ol�l���}g��vP��y�.|��x��$A���}�v�p̄C�L���O��%3o�:0/�M�e��Q`	������w�u�,q�*T����g#��~,�@�W71��9#uUo��_��u�j�9�7�j����f��8��=[L�����]� [A��s�hׅX�_���tYޔ��b��\r�;'D4H3ZZ��أd�׫�KoTx益��`���`?{5��_>���}�T���+�i����_RraU�5Z\y��Q�8��N5�vD��],q2J+�0�V3����a��,�@Ǉ^��bݒd�ܖ���b���Y��{���FB聝����) {$`2����BH{!tbѬ��Ξ���$̙���K�t뀞'��ν��I�*�؝)(���Wħ�����]q'5'LRoV}�s�2��LG^��0/ ��C��~��Mޖ��Cr�?�/�%X���;S2�k����B���/ҺV�~�r.[χJ��Q��`��P����"����b�}�dE�zIa�{Բ~��C�I�4�0$m�o��f�$Ņ�NO�g�G'd��?��	B::R���E/��rf�.�"��1:�v�����Ѧ쳕!�㉎(|�];���[3�4�>Hf-l����G�(ƻ��-�[ЄbM'�2m�;�Q���b��d"�1��!�}��P~�6a"��-#� {����(�]x�Ո��m�� m�Q�#Z���7�k4z�&Khz�0f3*����`j��-mԲTTD�(�e�)�%yc�K ��|]����q�[�a�yۡ�<`<�s��s�G����W�,��� ���D3�֎���	q	��)��;���0�$�������L}���H�nSG��eR�b���F�$C 5bGW�܋����E���p%cE�K �CM������S�l1���fΦ�����*v��UҦ�'����q�|)Ɋ�z�u2'�G���
�E�e�IN�̬^Od�t�a�M�n��H�Ym��x-����V6D�B���k&y��ʭwcT�x��?�ro��Pd^�?c�Z�@ϗ��G	Y`�1|� C��R����=��U���P���-FIм�(����s��GڔFV?�=��jz7Gs-���6���'(S TԷ�e��scߔ�5�����^wj9�g���:�Zb�3�� 6��z[���qet^¯�؝�jdx��b-J�)?q�L}?Z9I�o��	Ͳ�fʨ��~��wu���ԋrr"�W��x��X���X�7�����K��
�Eo落�`�g*	�>�p7��t��w�g�'M�4;�V7���"��7�"�6@�O��(��d�T��U�Y�䎏��*7rx���� ��۫����H<)y�D>�b��n�e��D�q돖Vaf�Γ~��-��.�bi)M��9KV���vw8)�
���	�ݢ9A�����[�o���e�Ͽ#�^9��+�mx�Wx?��2����ce̈�PD���Ʋ|��"���E�tj+�i`���،���0�E6�K'9x��U��-��D0�0�ZF��T�؋(;�>�ܩ�@��V�6��t����,�A�r8Sީ��e�
��G��Ү'�9��Q=��Ɨ�1ήeU�K)}u�D ԡ������j4�/~�N�!������!��EY����0�H�B�X�2���)��ɻ;�a(�v�Y�ȫ^ٽV������Y���J��l�	��T�`���[�B���w�s�R�6�	�'��Dg�-�vT��N��xA���r.N E��ë���=��{��.����;�����)S2��{q'j�Q�<{�^����J�N�U����l�(��)I`#���{bu�n���/x5sIK�ㅕ��(M:��ᴝ�YH r�r����z����UP���Z�O6l)>h���g�.�,��B:�Z��X��{��Ө�8�^Qu[�}S7ylG����<�/�j_	aξ.B��9�r��_�G0�����5���m�x������w�◐�^�=�6�2[hEם�k������!Fr3��);�1�A�n�3��l�ET#�^w����d$����|�x�����m�%7�i�핗�$SB�mM���8{��*� ��J�:�qT{d�DC�Ʀ��S�eJ�� k|Ń�t�����|R���@D�e��a�ʍJ���5b��Fh3��f�G�{��/V5]ql�]Es�)�ʂAh�H�v�jsj�PS��~�9�I�U�=_�t"�������K�$8��Q�%>�v���7�h���j��1�D�}7�^|"��0ݐ����.��i�?�����mbs?
 k���k��������2�3`�p�1�t�1�]�5���~�����yJ[�a9n62P�h.a;����Ґ�ih�g����&����lpno�)� 4���x���ꀑ�)]0-Sd.�K/}::��$�_�9��ۮ0�B4ɤ�c?�H�M��ȧӘ.�����D���O�%���ڼ�`�`��;��7ݾ�F�a)�"�� $�.��z�NC�bm�
�\���_�{4{=u)���&��Qf�L
�����Y�^9���s���JsG�em�se	����Rg֤���iP����3d���N'��َ4��u���G|���� ��C�Wz���l�>rz�Aa�)���w�����͏�ʨ��e��/(�V���o?�h�Q�p�{����a�	
γ4�l�IZHxU@�4y��^՚H"{|}"�0��s�|�j���.bj��u���[̿D�Q}4��V��Pl?�DGp�����u.;�+�Nds�V>&?h�/�ȷ��e��]�PC���Iu~Zbdќ)���[@o*OZ�F��jthVT\R`�?�&9�S����0����&v4�^0E�Z(hk8������O�\�����nY
�+�u �D[MT �w�"��?'i*p��R�+�Pa�g�t�O�%��|��7VP\�W�j�!�G �I�]-���
�'ѫ�E�8y�~���9ϷNrb)
W좫�M3�4-W�'��q�w,���3 ce_�qS�_��.�pۆ��0)ۅi��xs�0����S���S4��@�{�D���)w�8��M����6P�	^ZR�W!�W'�S�H�A�]�<d���H�����/ɨ@XU�:�>��m]���	�	��a�< �l�'^b0�}�O ��i��I�ܦY�VQER�OO{�=�霣=�|�S��Y�˄x�rN@���B76RD�C(-��z=�`��v	��=��<��#>����Y��I΂�/�P�!�(�}Z���F�u�au@N��H^0�26��gG�G#v)��k��}b�=9WO��m���#��d��8�Ѯ�k^'�p����X������u(  �	�*u&H��i�X�a�Q3v��߬��̕� �1�ox!+*���%��v�h-.�"���M�`��2��&ix�H��r,µ����f@��GO����Z��P.�d�4����i��Y�q�����CY�-6�(겨���O�|����G���?�;�`�[�v��D����u��`�Z�`����>F���2�X���ѽ��3
R6��WIu�E8���S���l��V�C4�FbCO�y7��$���	�yG�.ϣ,,fJ�� ���8�yw{F�W<�L{q�(-��24���7Bb�e�x��d�i����rg�^�A����w%��3I�@�R�?9tS���c�ǥ���|��ؿ��7 +�r�Y�������y�"�F<7ɽ	*�����(oÙ�ʇ��'>.6�F�i��y�#!����M��_B��R���yd��l�W�����)�t"59yV�Ŭ�� ����O�d�&w���z�7(QAF��K2�<�u[�
���β�	*7kJ$[�	?O�Q��в jV��.[��S��f��F�!�~�<7�p���2>T�3A��W����^Á���tݶpC=�\q(�/ u�T�Cy��1����6;�O�~1�(m�z�au��D�J���6��k�$\	 *��0����0�^�-ʮ��`֍��(k���Z�
PU��������ƒc~[[���BI�GR�l�Ȋ���.�6gY�p�C�O����"L�\%���'�Qh�~�Y������ߒW�:(v�b~��{I�}���<�F��	"�"��򘟭���i��!���H
Nb���qp��'�e�I}�~���f�3�a<�0��@�"��#wH/@�k��Z����GA4s�׫u�Q�37���Ϳ�K�J���:� ��=����;ܻG�f?���xk6_ƪz�.�YSm$k��ĥ�ږ����5���7ҮM��?.�Vs@ޗ�mS�B�3�oO6~��T��H̩\�z�r�'�n��<���{gAq��-O�Fy������@��),�]D�q��khЕ�z�l\�L_���͊t���~����p���/Z�6���7H5O��ZG�/bj��B��_}K(♜Ι�3����4K�Ib�j��!K���R;eGY���?0���+��0j�e����bG@�L	A���yVb/�Nn"°d�A�4��&gOl/q]�=��L�KZۨ�}�����u,V�+<1��V^~�`�@o�DAW�B	�
}Yi�����DƱ�4+���cLn�ϩ�i������`�XYaU��8J�](�vM�3��~(�a�a�30�~E�>���J(2U����B��ꠁ�y��x��"��@f�q~��p���H���mE*��Ϧ\9��|�a~�d8�i��r&lo���l�i��8���k�X4��L�hT~�y�vU���$<}J3Ϩǌ�@ #=a���US�Ib�xF��x�y��E_�Ҳs�����ś�j��+�ǹ���-�R���^�Z*�5�T���I��m��K��pZ�U����'�'m]M��Z�e��J�_���Gq겅Qt<�X�DZpV&���"V�g�Dnj���Ǧ������yܧ`�a����ϒ�Wv~��z9!�.Z0FU1��6����9��x:,�Γ�m ���7�%TI���\�3%��lM���,"�o�;�F�PyE�QO�}�lzT�O�s��W���73��@3V�U�y&v���Ỹ3�%�֞�VN�[n�\�<���ni00j+�-�B�³G���7\k�b�?>w\��̊���P�R:��.=G��%�0��T@�ZE��z��Rc�*u�y�����rq��yZ�-ϺR�h�TgA�2T���5����&.���V�4����qٚ���1ĉB����tXٗg���w� ��-�NRF��7+QG\��|	Ta*
���4$]�;�P3�[��0g[gy�_�,/X�m��}a�&v{����Y�P{Ȑ.�����i��FKߑd��)���R��{��@R��K����I4Q�����h�j}�c�)GD������������VG�S3�+|>�)3�~. $E*o`5u��_[Ш����2�Y�;�C\n:�_R���N?H���w�����/��������1���0W������ۖ�o��3��0��E`�L�	K�0ReNO�Sj�����R��T�a�NB���!��|a@�����E�d��v�f���}�,�R��X!��a��O�~.����a晤,�9�?Ep}[u_��le�ie��h��G�i[�t{��
�_	����-h.WJ��h�ͼ�Ca���=�����yց^�U�hn<sd="c�#9Cj����C��Pi>{�vm����1��q��n���q��7'����>��W 5����	��i3y��/���zkz;��emo�4V�B��ߞ(�U_hec�XP�?l�����u-j5�f��̂�zsb���6�Ob��=�@�Ur���q�-+{�4Z�JLjq�����/�'i}��;Փ�f:�O%��v�-r�҅�[�ʥG��D�@�bWK�=�����dx#�˴�M��⢓���DM��ݧ��(�i�פ`�\��Q.�=Ĥ�a�D�{�)�^�f_`��� ��|����r�
���{���Oik��i�����Dٱ�-\#/JMY�HH��'��c��m��Z��-'[,(��ڣ�s�cP��-|���M�v��gM�5�XR��i��H�ML�n�i�_1��$�oj��ok�@�����H$K7�/}�&l"Q��q,wG'��gNM�B�fs�亵����Yd����}��$�ci�WU����.�
�
us~Â��
.dK���_I����(��1�I2I��[�/u璬M+	*JaJ�g��>��Q-��w�'��$,�Z��#���+K�#�}m��B��\��G�p["��⾮d{��� a*�C����K�oݷ��s�/�B+4��w P?�ҙ�#�TPӮ�ix�Fն;ّ���O���J����]��U����YQR55�G���0ۑ�d���v��z�fpMU�K��=Ar�5��\@�)���@nO�F�2�`�����≌�+�����3���<�_��Y�)cB@�y+�Bo���8Z �K&�A���Ql�3�kǬ����.�Hxe$ ��ɅLb]H�w����[�_#gS͹������~)f�'��&��¡jn2u�Qrj����>\j���[5�c�Yr��C�7�FU��S#���©ꞷg���ګk�f��5��k�,yq!t�ƼN��Yzn�hƤ>Q��ܷr�f�u.N#ht�AX�]���Z���X��t��L�
fcM�����J���F!��.��t�s�^M
Gu>�mi����V���Q����mZo���9�KI����fpQ?ҥm�DB{����>�x�S
^h�����p�u��"�5�ihJ�x�t\���9m)�Q�P�G�y���;T�W�ْ�,���LHfH���BX��<6%2n�߆q��mO���1L0~4�6����'�>/�����E���s8���ic�Ԣ��x��H6M�w!���.���'*�E��k���
���z��(�D�+�@�]֚��	��;y|kw_��]BP$*�k F�㋲5�wZ��p��8��~�$Nn��tvG!"�ZmL��&(�|���?u��Jë��@��v1ҝt����,��a��Y7T.Van�=k��#��W��_�z[����>�_�T恈ae��\7����2R���W�����ܳ�Ų/��B�e�ߓHhũ`MT#����)�T{��{�
p�7���T'�5*3o5�R����En�!R�|f�� M;���-�t�4Z$i'^[�<3qʿ6�"��ն����Ӯ����Ml}v`̌�D��`c�SH�&����yŻȻD -.`�Γ���AF]�H�7i�������eEgE���c���z\B�G���ڎ.w�*M��L��T�׵�¹�&��s�G���G�z���n��/,��o1���:��=��q�u;����A�8FXS3NU�k??�����%�K~n��e�4���B?X��TY�^1��5��Y�ژ�:g�
5��	�!��GL{֭�h.��q-�����)j��M��HTY�G�=�~i�P.w_=��pB�|m�C"�Oů�/�O�Ӊ$e�wy����b��k��8(�;��T�k���_��^���W6�HZ�!Y�td-t�k}V�PY�f(�TxYڟ�c'�@�= �^@D2��;۫���ٛZ�>���+�:YM��J��ɇX��C��]���}
ߘW�-s�N&��O�P�r>��j;J��pb<�� ��S�qOn\��\����3��
$��vD�\��mn�1�R����d.8oA�s��<aC�e>x�Q�G��FE����/�|'&1Х�޲�qc
��<�"!j��� ء9�������Gz��c�Z�N����ް�P*�v���O⬓�#	P�l�v�B��SJ��7������� ����ʷx�p��=*N�B:�7��L��D���t�"��s=H�s"���T�N�S�]�3@%K��5�.k`����/�y�P��P1��s"�g)�oF����}�~��N�N��7+B�w2�p��ę�����;�¤�S��oMP�6H�Y�WU�Uh�ڝ����K/���Mc���o.���^E�{e�������w5������0��/"��~�����\�SܤS�w"U^巰9��2t�N�/^�'��?}�9����	S�[��Ps��{��5��ɜh�3��+,7]D�����+������'����jn�%� ���i� �Uu��hx�i�2s%�L�qP��ͦ����_�qB�e��m�7ܳ�+,�?�9���f��[4�Z؎����h�,��'�����J��'XW�9X�K��j��14���~o@`k��;�ph��m����k��"�M��s�wJn�91�L)��� L26��b}�l	OQ��p��K�̻���Kl�0�$�!� VP�CY�Ӱ��GO�$��ɣV�r7�Ww7�W�K�!3:_y4�Gt䡾�_��I�߽9F���)�����"�
�V;�	�<�����h�Nsy9no�/��M�0�]h��D,��Ԅx���pDe�V�I�J�~~Z�9�ڗ����nՊ�JG�Ĉ����+�E��S(˰�*_Kac,O����&?L���ޯ����m$������z� O5�(<�����Iծ@P���e��׉0��-��77s�aK�H���}�D64�t�u1N)̀yi�r���3�S�1���2���h'.��)*D.��_"]�؝���p��2C���n�ZL�H� yqV#������1�KW��ە뻊�X,y��h��!sE1ֻ�v��|�0<Ҵs��;����wF�"3�A�ҷ��9|�����LQ��L��Y~�����)
�]l�wd�����u��  �.]���ߏu �^��G�Erih���������/�+�oj�����It������u!�ռ5ЅqTZ�q;)�z�P���L>k�Žڄ���C�:"�9���G
'ϭ=��p�Cvz��o�2om$���CP�L���=f��]ð�h%�������}�#n�!���#���&��כ���h�I��+N�Y�t�"3W�\Eo���jO�||8���?*��1l|C,���>��|�n���Pw#�!*?���#��_��s�Jg����*�ۃ�_�-���t�H�t�tG3Z�ِI�����&�X~A��D楲��X����t�,���<��@�x=�dn���Wq�l&3�e ~����<ܙ4��z���i�����9ٿ0qq���@e@���Ae��3ކ5�]\�B��`O�CT�,a������j�7b4�_r�����ʏ!��m���vÁz�uTT� ��A�/�å�����T��.<�*n��Irxq�)m�*�^��"�z;�-c"��ס���{�a�UK�1L������u��	�q�	!��;M��1{��VA� Ը^Y����/����M'7m��]k^��� ��9
ř]��5�y	U��/�n�a\�4��T
��{��:bg��Z�D�^�v_�"�#�aK��X6z����,Ϻ���2��[�����ӹ�d�ќ�O�I��(%�f�dS�N������7��h���|�W��g'�>Oh�AnaOIpX�X��1��6Sj�[�X#� �[ă�q�Đ�l����)\��
}��9!=���Q�8ے]9��M�_=�D~�aX�2�B�B��&����dϮ+��̴Z����ZQO����g�5T|y�AU��� �fUH79��>���p��m��M�=��>-�iJ�ɲ�<[���Lj�{3˄�vJ`�&=�8�m�}w��m��!,c2N���KR_���ʺ&w�R�Ds`2Eqm�n�~�7��S*�{M�e����y�A�w|tG�$na]�0|ɚ-�`�V�+��(ᇉ{"Y/����K�O�
�	���OI�z�Hb/��x�_��iq����/N7I}�K9(af�M��aC�(|H`0��,@�o�e�ǒ6�xZ=ړ ��Nvi6\����OfT�a�ͯ7��&�n*�y��5+��U����g$��ڌ�]�`��S�%���%���)���gd��)������і�B/|6�7<�qp	{E���64�,��aM�X�s��-9f�H@��'&��툼�e?���ecY���K��Pn�I�	��R��f��~C�QK¼B��C��n��W���%�R1��� ����_D�JA��+rjd�\q.��WD�❬E+�ZW}��{5�ln�Tu$�*�s
�1'�9t��-�wx;�+��e�9!�M%�\7�:�fw�����`�~�D���)3qo&'�5��E�7w� ��C�wo��O��F�����}�� ���)�oY�m˄ ]�M�,�=SE ��u��"wo�	Ι4�؈K����Xe�Vh>�a,N���2�m�E�t���>[i�"d0h�@��lxU�H>@[��sv~;��#���!�m�v�,����С�T��P��c��{�R�X2����>��p��F�׉���е������t�q@��1��ĉf��G�z�C�p�#̭���A���gv�n�<3WM{8"׮Lg��8l�C���&��R���5F�	�݆���,g�-g�7"��h���t���I%�r�+�v�H`+bf��tH�`��U�ȵ�"�^�i�Hb0Cv/�04G}�'�Τ9pR�D ,K!C���d�Y6�ބf��j��]I�~)�S'"VWb�g�D+
Y�)EK����f��U��q���O���vJ��œ-�"-��&J�-�a"�O��B06�B���ӎaJ�����n��?��j	"���9��JI��w�r>�A\+r�|ֆ����.J��K/ge���Iz���i�ǴN��\3t	�O��	�5$ԇ!��F� ��QT	r�}.�[�(�������!ق{���u��wwe�б�=�8E����8n��-�_�¦��L5;!
��԰�P�O����Z���AR]�r�[�؝~\ՠ|˼��6~<����rik4��N�H�|��ZAZ�V�b�/d�qҢ%��銪ԝl/QҺhj�����e�(�P?\hj2���|E���K���V��-;3�N�YDk��ܤ�+R�����k��i[����c*�r�{����*8�9���_��P�޻(T(L�.�/�G����ʑu���O��Ƶ���瀰�(Mf�P���hUe"=��������/Ҩ��څ�_0�-o�
_:��?i�~%������w��,�ߵ>�=���f>�!����C`�c+
�Er,b"�wֺIj��0�����쇱3~�쭝��.�� 3���]Z`���G�
��݀ob�hr+��[9�J�0i�Ha�?�T���I�AZ��uq������d^&�w��M"VѾP7'$!��e���-�a�=�Ѵ`8��8�΢Q� U�AV��y��t���z�*6��	L&p_�]J�j�Nʃ�2�!pM@Ph��ea"����v������d��/���y4�@2�ym�������]өå����o���9
���\��g��f�ޠ������Ҥ��9cs�؎���)8]�G�#�s"�)E:乵�?�	�'���8���r���X�������
3�z��D˽6�R⌅��~&X#��R~ 1A6��e��0�]��|i��l4�S��N�N+q��bx1�`�~Ϡ�fzK�{$$M4j��	mX�A����RSw�
�bL@D `�%�s7,\�c�p��&aM�����fɿ�|�1��^S���{�OU��]}2� ����}�W>�-�zn�}��A�
_*wt���V�R�wK�:|j3�A�������l�t,E�ǆz��w4�F���g��hM���X ���@1�gWS�l���.�2W��nG�����>�r�=O�I�-s|9A0#������}L����F�C��2��bS
<J��fep"��>
v�������;�»\�Ԭس����D0U�kï�����ڣP۠�|]H;�Id�����Ļ<{���R?5`i]���c@���M���gq� c'a;�hw���U-M^N�>U�P���E�&I�5�[t�m��Z�*�R����	׀cUϋq}��0�Ul�N��"x[0޿�\��B�:�Xan������cDTo8�qO$!8�	��� ��ɍ	"!iw}}�����-�y�ta�����M#�d�0�H��|��*A�Q�|�ʑ^!��h��r�DC�b�?V�$�.�u�+��ϧ,�e�1Q�v3��wG2?'C@�������.�����.�z��ÜS��p;�N0TA0��hL���f�8G ��A�����P�4��h���aS�zp��z0C��Iߧy���M�hC�l�6���(�>j>�w�՞�o�	5GX�</��7�`z[�kdN��D����Ør�/R�VTĦp��1�ź�|/�%5���o}��s�� Uʭ�s��?6��"3��"iO�W��[��[E9�Kb��n��,�a6A��q.űr�i��s_�����y�4�M���ٻ��_{4�I4�()�1���%����}P~��Րu��Rw��	yTZDL�u6H�.b�k'Mu�~�O��D
~����vg�pp�ЭxO�(�]�\�����u��� �RӬ���欷���DXm[�xN��2���S��u��&Q"� �#��"����tGؕ��&BH��MB����D�"��4Qb��,��'��S�О���\6�rǺ���%>ømW������ܤ��g�B�l��,��u�;}�\��2���,!�Ҧ�m}�☚No2��!�&Kr֭3aʢ�F\�+�&�N~ߔ2S7	����m�Úw�E���9=���i7�Z�kv��3���c�B���0§< 0�%���*��6q�>��®�p-p����Q�C�/m��x�L��/%tZ��H	�/����E}z>�����V	��S�k9%��z-�Br<�le��Dx�!Kmd|H?�LjH�*Bx�Ac2�v!Bv�㩈#��X������t�>[��kj���Z|�p�O3;�Ԟ�ԏ~��eNe���E1 �� '��%|'���^�v{����7���:V���WXAPy�mрf�|������ɷ�+�:j���a��Ic��X�T������8 lD�{#���.�s�fD�x��d��� �I�����8��|d��>�P���
6�-�R����8fp2c��D�9�l����7�M�G롇qnPd.�������kY6mOJ;\��櫥�2�P��d�Qg\��H0�\�V{��]'	W�I��-��������o|������Z�&]��\�GG�����  �Q0��~�;��W5�?z�Vt�$���Ҭ~���C�R�җY��>頔��1�ϲ����*@��tW�~��n�Z�Ok��e�+�p: �T��t5*�Z5L6�AwOX٘!��:���a�<2w({�O�h��~�q`x ��O��z�t�E<bo�t���\�A�"w�Xλ+F�1��V������ػ�Zy��q���(��3�M%e ���*"�����m��Z�J��{�Q�I�G���=�*$Vz�w�ڭM�x�o�:^��04^�8�Ԥ︬�O�F9��8���A��4bWs��<�o��Q�._.�e�&�HF���&�l��a7����=�v�Gj�VNm�5X�1��Iu��u�pÁ%ٯN��e�N$����O@H��X����[W�շ�v1�g�V��5w����L�� �݈�`�~�7�]h4&YƱP�]�������X�FBQ/U[�:`��r��
�1���J3"�Y�qaXj��Ol���|��A�쎪�=^��\<4\��俼1 s��<6������Z�HB*�\��gʁY]�Er@V�x��_��d��i^��n������yA��獳0'P�4�rפ�=��u($rt���.�WN�R3ʳ4E]�Ь��g��jj�����+m9�Vi�6���탘͚�R�7�7Bq�U0�#�=��%;N�5=Y��)KvJ���"_�Q�2 m˓�@�f��o�>Y�4��L&�����Ꝭ��O!x���������H��[g��n﫽�;�ŉ�B�1�P�m���j/M{� )*s���4?7J+�-8s��\?4���a�:�[��Z�1���
%E1�U��	�I|�y?	��>�c�����^�����t.\X�kg�m��!g�T����̀���}UN������r���Xpd��L��Ԧ@TOgI���-�ĶE�
� q�3��"߃�z%��$WGRߏ��>bW뎍7�+(����|M� ���kaF9і-J�na�yn��U!�ݵq�EJ0�������$M��ܶ��@^I��I0#X�%}�h��\�]������%}]��m��
2�%��K��Q�L��gy�p�J�Ǐ|<]<�/k��r�PC��jP;�� �i=��(l��%ވr'�4'�[���#E��F��-��DGh�0�p�{��-��S�����z�E[����r��zɠ#[j�M����g��(1�p��oVD��w�H��r�OƤ=�R�"��E�p�½!-�pո���Zf�i���8������QK��N�O�щ#td�p  ���RС�Y�qz��t}]�W�l�r{���3nm�E�W~�}6�������A�/�0�t�5��ň���l��sT	j��)�pA�TҀ��I1EMjD.u���B�ZT3���n���B��$V3�F#�.���d��:Hu��a`NW9
edڙ]W���-{���T,��ğz�ֻ��f�ӑ�n-�*��Ҋy2]5)lPK��1�Vְg�@����9N�o]M8l�'BEn�c�þ����۬���@]\�d��I��X3F�E�v��}y8���Zm-�_�P<���;��C�ĸ� #���(� ~�՛�Y�d���T"r�3�y�x��g�CF������j�`� t�hN��51���en�!��9&���!����.��AQG�-�%�U�*�'/r��X\�h3�% OYV�9��6��-�Bd�yi���f����.I�*��Q��.��}�F����z�<(�tԀ�'cdج	P%wj'�8�F��A�-�m�;|n��|fNU���f�W	e��"F�WP��ﷻ]�Z��E��ٽ�)亃��!�yѦ~����`f��ك��������.l�B,E8�5� 5
۝���9���o�r����(`�*�x��Z8��ge]w�Db���O�����]�CG�^i��-�9��s��?-29ڭ⯧�M�v�(
?�w�<9��~	D2ǥ5c��׸�XT-�\��;DN��
���]"q����2!��/��y֓�!���K�}��H.r���F9O�f�C��fA��~`t9���\������I3%b��W����Z׳p�w�s~�������npGz��A#�ğlwZ'#��7ť���l�y:�g0x���[��RO���a�G�˞��CYO�4e_�+c���:��*��M��]����w8���o�[��b���?�Bd�/mAWY���^���$ ܛiWH�q�@g�L���ι�'������S���;�d��I�U���r�1C�k���U}˧�G�����'����;�3�i�`ˬ�%�-�ѥ�^8 c%&�]򦢁|�	���ěG���OۧE���`'�Ѷy���yt�=��0>��@ ���݌2�m�Ʃ��YD������I�X{0�8S�~N�!�j8a����F�e�0'���N?�.Hn�82{-
��s��4���/�c�G,�(!�y�,˙3���`�����*f[L�݀��*�-�׌c�Ԧ��Aj���d%Ȯ ��>�.ER�9��?��^���>Ѷj��n,�K�����3-M\��ݫ
|�h2f�����O�,����Հ�J�߇��rD�����uB
U�*äe~���K��B�j;֔�߰�`�;�x����Ę <�����D.��bht�N�U�
/���{x<#Z����J�PG�m��&.O��6B�� D�B��!i6l��*Q.����gnO?S���A����]��;r��<�j=�3dK���D�<���M {���ל��3���*ӢK���s)�HUCQ��v���C���d���dB������Gq���;\�D��0��n�c�v8+β:OOI3�kF$-#kޢ�p
�P��a;��a^n�>I��ώ~1 ]��^o��clR�@�h�vX�Q\����c���[6�K�p��y��G�]�4)�4,�E6�ň�����3��;i��b�K��,�qC��s�&�����9ҙ\���đ�Ȭǵ$��R)�s� �T�3���#�YO��Z����b%������tG3uu'�q�\\�zQkZ@q�ٺ�״���L�u�Ԉ�<&���~Iۧp!�I����KX���Bΐ|��mF �B���F�hA�؞�Ō[�6�zn�I��Z����42�G�Ѝo'{���˝����_�_�Ե��N�%���ps�O�|Nvͧ#�Q�~X4w���>������=��N�ҭ�s(\�\��=��1BγS �����_^��~�q��S�F�U?G��릦�y?�U�� u�ǔX�٘���Vw)uxA�S��s�G9V�5f��+�꼿��oS�������e��a�����6.�ݷN��hR�����x	 ��5��X2Q����p8�[����~��(� ��� �y��~�&�uu�H����y#�?Pk�	��=Wȉ�R���}	q0��,����vt1�*�#�c�3ecCo���2qεu���%Q�k]�v�R�S9�?Q�H�-)���'�]�0֚�.���R��(�_��֎��'*&A /�ss�#֨d����_S�4����	��*q��-?sȠ������4�@f�I��q�{�1����h1���ɾ��z] ~
�-�X��V���!s"�v�q��.ev<5��u�����9������~@��^�q��o�v����#\�B����Wrh/8��N���)$
�L&:ᔵ�\gF��{\���C�����?�K��sM?O��59�i,����@��`7z��	i"�Uo��5����ZC�C,N}�:@x"T�k�<�x,e&C�%/ng���Dkad9��~��_�$�K��.E�eK��|�X���F�� ��cVH�ǚ��:t; C�=����c�{*�� d����n(�G����&ޔC7˔�d��&��٣�[�A����}[޳�3b��Z(bk��q8�1#ai]�C��'��)z~�#\o�\������a���0�g]�Q���-p�
�/D+o�5?c���y�UM���J����,+�%l�J���j��-,���:�_��ɻ�b\�~N0:�G���zɝ^x�^�gD�o��r�
��Rƛ�Ho�Ț�(߶�k�h	=�Kyxaf���]�����W���0�|�d:l#�u�Ro�n dG��`҂�v�Q�$F��/�>o�9�����T��C���I�t�vHV;�ʙ{;�GB�냟�4,�{��S��.�H$R""��};��&��
�o���v�s_�"؏L��CE	��)���͵�{2�<�&�����7
]a�RD�ǻ�h0�*hsL�ѳ{ɥ3�I�+ko���"�3�E��@�xgR�����>����L�lI�S`w�����g�3{fGFh"���ԱhR�&l�̘�Y!�� ε���3������e��k	w����*��߲��9=���Uy齳�}��N��Ao���":K��D��R�E5j��m�x��z�����%���($�T6�y��ܕD�W��-��ޗ���D��Ez��I� a�[��CT��Q���a���0S��:�t�wޱg"��.��Բ��
���xk"���1�ﱴ���B�Y�mؾi��A��]���*MN��ݰc#���\G=��^(���k]/�tc�B���Y9f���=J�������cx�h1��E��\:Z:n��,�)����ůb���D����I�T���ɀ��o�ni�1���"�����rS2��l�7�,t
*� ? u ���V�3�xX7	}�b�����/'��m��:��$�iu$5F&A>����$����o��~l��w��H�rt����&��K�j����"��LAn������L���s/�x�g�/�5�T#.����i5�b?��a�*sa#�~�Z@��CAt���}�p����@^�5M�t���D��h�1���I��*+�A�1�.k=����eQD	��|�`��:~[��������oR��M��B�ُ����m;�3gh��[�C����	�f���{�p�P�0������o���������t;��a�kK�ġB�D�L 2�I	&`T{�5�i �>���{q�|��;,>��3�@��	a!&�3�bH�fo��C��ğ�_ُ�NX��d*_���΅��X�QoH暝�%��2��.�:|��m�)�Z�ݲk�*�o��2,����xW���2��M��Age�o����I����G�%<�F��-&%��
a)$������8��� �*]��w0��O~��ͩ�I/-��~1=z}U��C(��`j 8��p �E\}�,;���ԻZ �⩯,�'�	~ۇYd��-͇\�����+�@`6LH���6�l�@��N���S)�m��{�i~H�F�L�6T�<�K��l"任��췶���E�2��Ȉt���3p�T�M��}!�!�T�zCƶ��Lyˣ�bPd� �f�1�{r�t�~�(@�^�8k��M��푻,��Uð���H���V<����41˿SMѪ��֎}G�?4�j%��2���,s�G��}�^��{@e�o���������#z��8���k�� 9�d�|Ű;�;�
�-�i�+�3�q��`$#:�3ى��q4p��l��a��`Y�;E�>��.XGY��]<?0x�\��"��=�qS���o ���|�L���� !NkYS��|b�ĸ��f�s�嬍�B��d�߀�D-Ւ��6���!s�>]���",]���9�!U�C�exئ�ю�^e��6��Rs�����(�Q��[�<plK�}!��=�+b���'c=�@�NS�Dx�gVaᑿ@N���o�"şG�Y�U�dٯ	��0#�x���{Г�t��߁Y<{W����n��r��
E���� k-��Y�_��R������oܤT۟W*�KSP�6��A0�,�Q4��/�FDw����������g��.��0�j�l�@����e(��K3@y�ਃ�>J�R%����'L���i��g�$���-<Yb	Gm��m��$ٕ�.r�S�x�S��((#�6�G�����RbߺQ�ޑwB�s�rCG�։���<���ҚZZ�z6L}^�J��#���د��0u�s�0;�z~����!+5һp	�Hu�
�����m���n��:�7�e����4�����Y���2��N�;��e�{��>�o˶i5RySZu���J�.i�t���<�ƭG��_�"��p��Ô��wMO�&��ÞT�f��i�DH=$M�g@���H��$���QplAa�+s��8��"?&BR���h���ˀ��S�8�j������A�-��q[ޕ�g�c9V{gR���i��S�ē r5�gY��<�_�g����:��fkE=5�b䣁���
�����*;c�P�8��T��{"W�G.�x Vz0z�IO� �����yje��ʗ�8�D�fU�.p�:��	-�5�骷ު�T
���<��]!�Dݣ$7c�7H�J�!'}���AiIW������D��]je�Ph�Y���\�h���h���2��\����|a�z1U<C���z��-{M_-�)U2���s�?�B$��6���5K\�t;զ�Q4�޾c]�O�@�d�/��� ���n����GP����]��͂�|���p�T����Ę�@X����u�����-��uX
��mb%0�	�y��ej(�ૠ\��6L�QJE�ꗒj�@ў��+\��'<�n���r}�`>
��F�<�����e��7N�?�P#qN3��H��M�|E=�3;�~*Pg����J����^Xs0�Y�G��Dm%�����ݬ�laa/��������!�Ԣ��ȕ�>5Ӛo�)���\�����j}�qxQ-��5\����Fۮ2��;PX\L����ٿx�6�]Y0cr`fǕ5װ[?k�Ț�P�/��ض���w6D��(��d�l�6.�q��Z|��?��J)tl�5�b��3�����</�L���)��l�|Fh~օ��C��t��-ͬ��1<��Ӄĳi��d�u��90�`?�嗑4�˖�8^�CߢF�!�]�kH#[��p���F���kƝ���q�$bz��q�r2�
]a�9�ԣw�=T ��`"PG�*�6�{~I��%��,�$�G�h�4hm�!	������
c����b��DY�[��v��&`{���fb�+��5r���vk"ST�y�
�m; ;��x'R?��s�I�Ϗ��7�^��R�xeZj�ۈ�
�)*��$G�d>����^���?-�	?
?�jVq����э*`5D.ie�A�I(�FX@��ƪ�U�����W97�#gAf���,`�s��9���j[�� ��D}P)+�?՗t��3\f�dU�˿й'45a�9r�/!�S���[-���bv�~�.ޠ,-T�hF�%I�.q�_�5xq�Z���3��Zj�M�I���ǿ8,�)Xv��!o�Wʰ�[ �=
�d�-K�f�@���*IG��yG����G3ka��$f���.v��ںDQP��'J����.��P#ҁ��4��:m��ٚf�n\��^D>:���`��6l��k��-c�h7��Éx�k���hck68I*�'V�g��R�j��*p�4��\�BG�Wh��6R��a�=L��ҿ­8�mi�B
�8�BwX�Qf�6�.��z���o����O��_Z�^ Ε6�B}� Ԋ�n��ȝ��)�U���s}5��'	��q�Y]8��:��c!C�O�VPO�$i^R���e�"4C�ҧ�du��V�v�kE��~,�@�#�<��^\i,�0=~��I��D��p�0��mR��@X�=�㽅MS�AJ�Ft��5�{r�,a�?�n�%�"
d�;锗@�<8$	�4�3���vD~��I
*u{�Ϥ0����k�OX\��iA�Iݵ9����/�6��}q�>�&l�`�5���ʵ'A��2�>}:�]w��C�U�bz�	�KJϨ�
�4�Z�T_��u�����ﻹ��y &X{�rQ�V�5�	��P����3�U号��}��P�-[Y�y�/<���^A;�lp�͵,�����n#��~��g�������E[P�W��K�����ѡ��,yUA��g���γS��Ƙ6Z՝A��p<Jщ�/W���\/&���\uFC���8�83�|���1��폰},�Q���lZ=��FM����K�E�A�ߪ��jJi�����+�]�e�έO�ς�Z��	o�C?�M]fTX�c�J���y��z�[��{�ݖ|�.7m�Q��2Vp�3�$;Î�:۪����`ީ���:��l�����6��ɮ$���K�s'+&h,غ�NP"	y��Ƨ���Z U���u��L��{J�*q�4�?�25/d]�L��=S�}����-=��l���y�ʐY����t��t�G�	���<�uۿ/ɚ��Q��厷Ζ�I����,i��p@�PMe������<�[=���w*�5�'\"�����&Z Hh`����O�N�·c�a�a-bğ3�����#�D�0���3۩"񡮟)l�G���a��!�Bg>�)f��}��sG(�� �2ے���zȞ�W�C�����H�'9�2��Z�����Hp5nAbioP�*��z�͉�F��ue���L!1O%�T�ŏ�w��/�'iqm.FC��ɨ���u�u�<aj�r	v+a��'�ڨ���\j6ȓY0���Lob/�Iɂ��i��R���Ɨ�����4Z;k:����l�[ g	�͘z�W���:0<���:5���e��A[��zE8ȕ�T���Q�s_3�(��]�3���8�zz����BGo��ُu-0T5�Ƙ�M�lp�t��!lO�b��8`�:���¼�O��p|�>\��u��ϙ��P4���^Q�(2�pgp~�i�ߝ�UH�Q��|���\�W��)'�I��ֹr��~��鼺},�)���u��\S7�����ҿ����ԥa|��1ĴPsO����B!dI!mo�kv��/�Ж�m�uT%�l#yI�p��C�����2Sl�M�e<@���Pߎ*AL9�b�������O|��m�����YU{Ȧw�kd�\� dq������^0��D�GR7�_1�(J�IZȵ:E�8�j=�v��� K�Oթ�?��Ê�3N�����?��r�s�����a�TO)��5c0(���ߧ;v��mnh Id.r
�*�`A��k?'�l���`^�� 8_Y8����\@$9��XX��a5�+��Q	�D�C��߫"���ݚː�@T���h�����֖O[Q���3g���8�z�g���õ@w�Q�����(�[�9,F��=�V�yYWޅ}��>g "-��W�IC�H��������D������zG
���D��q��B�n����z=�����'�'d��f�޶��m�Ǳ����t�<j�وxk��fץ���B�iȎ���W��H�L��c� ���@2)�/����y���b@�����WA�q�}�h��L���?m\�v��&�t�f1�~;���l�FNjD\��-kvmM4�1����(����7S[L(EO6�\���\RV'�3�D���T��*i�6�3X�,srk���ӗ�FZ)c���LXV&�,6���(���XDc�����ZD�Je���)0�;}��+Z�N�5��&K8ŕ� ���� ʚu�9X�\�Չ�d��m�7�  ��� Z���|0�brdQ��I�yUݙndb�+7.z9p.��W�1E�H8�:ay�R��IS]f��x�{j�o[�Sqܨ�#MeF��и
�w�]wJtN��vX$�X��e1��x�l�1���?�yU��ol{f"����ru�!��_��5yDjwv��0 ����T)pI�6�#�]s ��I��LpI29,��5"�3X}]��^� �ƅ��DO�(]g��B]�Y��O�ٵ�f���ӻ�]�k�S_�`(�kr�����̮?�����,{��:���qrc��(�P}����h�n&mF��\���u�k����5`�#ݳp����z� �9�VT$����Ɣ�A���㱥b������r �]em�׉\'$�9���ɍ�`���#��Y��2g�_T �$������f�瞽���[�vG��!���Y���̏���&�� u��Oy��h��E��V�fV)�����	��c�;xֹ��$�+	����̶]��ndB�Jj��5�ٖ.��RP���!r+��ǲY�G {�@��Mtg�^1���b�E�*N� ��OY�����RE��)�H�t��c��ʿ]�\U\�5$T��Eb�U��o�@	�R^�s`6 ���h�V,��iJȥf�)�	���� ����}�0����>ޜ�� &�6ʎJ���%\���p��?�}>����!<���� ��C�{�ieڃ�Gz+:�|A��N����f��>Wk~S[O���?�~����fVs@��_�6>���3��}���cpc�DS���FN��0%�I���q��O7�~���e��׆��Jf��ݜ�8�Is�Y>�2��(ܩ2Zv�b�M�Q�B���^�Yl���ޛ�e4���k�̏'ӳ�����wsgvE�[�0�OF[+����V+�,{Q*��S�����˾�R~8F�ä?�5��jc*�$ˌ������P����Yl��c�"Sj6�_�H˾�4�A���k��t��&x�/sG��t!x�KX��9�Ǩ]4����Ko��_1��9��w��a�������$0s�]'���wQ��������"P���𺁤 ��jC��^j뼃����Z�	�(�ukJ��J)8S|jEB���� ���a�L�L�+�R��$C�5�6FF�j:k�A�y}6�U�@�~�o��߃��G��ղ�b)��nӺ�{��1�Mȓ��BS�ESY�?>Y�FG<?h]�%�;
�
���z�X.�2��9W�����g�B����!�f�'�x(itJ5n0g|R���">���e���1s��^$�&xZ�{���&m��]tJ	�/W'���<�� -�C�/�yW�g��~�\P��ߤ�G�H�$8E�eH��R۶�s<ML_�I�j��=ذ�KV��	�y. T��>E4+����$=O-��B8���5u�b�	�#��u��0���`��N8��'���կ>V�,�i,^kB���W.�Bv;��"�L�Z�U~���Å��Cdϐ�4�C�¿����
�&�~42\fU�N�!ٱMG)K��y������U;,�]`BF��[%���OD�S���y\/f]���i4XJe��<j�����G�,�r��Y�-A�?$�"�����*H�Ŭ�MN8�#]��h?3"����`�j�� E�x# ��M���T�"B��d͛����%v�׌�rVGu����ƨ��. ��r�c9���:r���#�x�2��>�\��LD4����2.`Z�>U\����α;���v�?,�	�E����H�6:2���d������0�"^g6<n�@b�f`O�W�U�_Q�.�Z�~��J���9N/�r�[{��h�{�@�*�����lR�#�N蝡k���u+�s�gMu����hq�����T�b��(�8!w��	�~��;�vR�j�S��W�Nh=p�x��|�)3	�a�� ��F�_���mS����Tn�*����QS��ʦ�4ʲۇ>��Nqz)Z��!bF����OQ�> t�v�?o�w%��F��j��6a�U�L�\���u#-�V0�G�\i�����8<�\��Yp��/fO�����e�����ŭl�Y�l��x �����F��E����.Rͬ��1qd�݉�-���c�y����\��@!i2���ZFP�5?�^�x� ���7O�s�0��Ϫ��s��e�˖�V���@���t�����X�\iTz��=�Z���;��C�O���H����S�rLʩ��~��x�l�t6��bU�ũ�Ţ�f����n�0W�{�(4>�8�2p/�&'�����/����/���>�fcc�n*�%u2���x<eJ*#u�-��q@��@��3:��+.�a8����:@�Q���J8� �ݜ�(�����F�H��0����#E*���_Sc8~�;�v!25.�p�Cme��Fw$�|�F�3��N��W��͗���9��.'� ��Ds�.tʍ�^�v�2m�A�M�y���-n�v��0j$L�̍�o�� ���z�h*���d>��� �J�Tn�T�(���r���6���)k�j������/�N"�����z9"�ol.`Fp�ݑH@��r@L�E3�b�T�|����hr�JNƚ��QMh0(�j��Y�kL��wz�}<ړ� �Ԭ����<��p�y8	(6�s-~�Ll��r6q�����w��ݛ3u�����Ϡ���n����&[8�`-X-.��(����(z�ֱ~iC�����C�%,W#��j�9ؒ����e���a�Q���CG5|m�ޯ��A��*�*�_���I(���+l'�EF�[�t��܈u��ie�R�nx��-4��?ڶ�kn}D}�
��-���.��.?��h�Q�����bz��Q�5R�6qd^�.^;�s�����;2���M����y	�6���L��A�m~��M6��ʅ4�p�N�\Tહ`�`C�K|��˫��y4 ������Z.I5�����.F�[J���?͙��? 2;W׍���~������I��X�[c��/wt#�ـ�Rc�1��_���:ih8s� %l��J�@:��J�wDZH���^M�;��P]/�������;vN#�T\8�Isr<���A7�0�E-�����4�d�Dq�ir�pW j��
�f�w(d�_&��3>�ݚ�0��4���gl7��CH@��r=^~�qz?�lNrE)7�kuZ��NBؾ���e��Vy��@�9�l3�I?R�{�Y�*؊�G�4��5#_�*1�%`�O2q�U���8��;5>�@�ez
:���[(��v�`�V�Ŋ�曚˭`#��b����ܾkC��/��q@r��s!����E��h�ԯ)<�n�j���>���&�i0��F���֊Q���^ƺgib�������i*|!����C<>��U��XBF�`��_G{%]���e���>���x&����W�7U��k��Ț���<ƒS+G̡�w^/��æ�y�CWѤ�І#$�w��p�&V��Q�f:t��Td
�J�&��	��W*��j����~��������X�t@���mx���iI���m��P5��D�A�:��/O����^h6I�E������~�#��ߙhO�`��A/'�eO�O:!��lə���|֠������L�����4I�ֺ@>8�_������
(������T3�'}(x�GK΂������X���v�O��� �Vc����D0pS
\��&�n�':��qԈ0b�4���]
��+��f�S61qK�9qzc���
P?���VNY�@�,2|��2٢|6|���B���	$_�~l�ցta��5��՝�a�$�p*�H�B��S�,Jׂ�0�,��'�T�4r��.�r�����j����3�7
��*#�qN��e�ʍ��ik�a9HC���+5]H��䤪���uS9��w߾����	�tQ��ICG�����/G �/�	�p��2�k�g(��<ǿ�T�m�����p\��	�R�Y@�o����D���&���g���{�������aO3'v��[����?�s$��2>��Vf۽�Jr:`s)�fhsoԉQ&��[3`Z�Z2�B����P����<�7�����ǹ��-�V�cЬY�s�g��<�Mc`�]�_I�Ef(>�4)����b��;vӀ�P�W8a�k��9� y!���~����GCY$�.|X��f�*�N>L��/���T�z��E���F�t�jB-���u'5����a��tŬ��~$��TB�Ŭ�j`.Cn�-�Q�P-e�5h�(?���coDt{=mS�bEMf��X��|CTX�j�9�ˍ@��H�S�~ר��U�R�������3��=�r;��ky�9�r<�NִgJ��z��s�4H��ܼ|�w]�0U��D�;Y��G�J-�D>�nm��p.H.�_p�C�j�˾���4'U��U���?mК�.�y�����	�k�߾S�>b�PiB�@��>y-�zHS�~>�LG}ƺ��S�[s�Z�F�mVy��<t��oJȒ�o̒�X���V�,n��k��P�V����G�>i�Tl �(�ng؉a���m���!Q�_��H�Dޣt9��{�<"q�{��*�d�@�*���+ᶁ��}��B�f�	q�9���i��;�[����s4Ƈ��
b�|��	P�s��V%i��[�B��鳗��h8�־Ԧ<�p�p��C+��#V����(�p��i�j�m(ս�	F���?�v�Ö��PB��y1fp�<�g��FOcW;:6|�����
Kl۲�*�r����:���}?���{��V'!����B�˘I����^�[M�۰l��g?�*���ս��Xiܷ�#�N׏����N�����'-����y��}�~��̌_��z���ϺN_�
Az�qߋr�5�# �Zp4xjb�#�<����*͐S�����W�cb��\�×��M����GHMe�@Zˢ��L�����M�6'u/�|\���lG�����rh.{r����+��o9��֙&l��+R(G�p�Z�Q�ڀ����H�$5-J9�Ɵnp�~��7|B5������v��,�t��Ϲ�� ���#�]Y���@����*�T�z�˱®�Aޘ��h�.J���[3��˿/񣄬I�:���>/v�����8�cڤ�'b��ٝ`B	��ἴ�J��i�� Ȕ����n��q/ڸ���ҏ�o�ȀÎ�~��D�*/�I�<g�o���	� D���IX'(sOee�^

dge�����I����5����� Cd�>k🥭g@?W[�g�Vaµx��*�s��A�`q%��u�SA��ɺ?�{�w���݊d�I�HJ�p��UR��P���	�o׊b�>�l\�����p�'��)��`�i���}�9�/�j��/MI�X�a]�դ�W�����FY~�~�ܰ�$��@�?�@�CH�O&v���D����ܔۙzj����5��r������7E�`4ٰDS=���=�-Ǒ��	���ΔǊ��"Ԯ�R�g��h%! WI�Q���RQ��6k�~��yN���h�<��������:�_+��KPm���2r���=@�����B��ĩ�G!D�$�D�Ө���$��_UͲH[-�<D1�F��5���\��.�e0��ߴd��@��&ܹ-�)�c�s�/�鍓��(��!��I쪘M�d�j't�i_]�l���1�psN֖aF�P�ws3y���H���eJX��T���m�Q���sr�fxxW��OZ�g^`�L5M{G�米}F5=�@r��Og!�O1�sy���Q��1a�R�����{�ͷ�[c��s�=��f<�u��t� �R���o8�QG�+5/�KeV��ۚ�_J�*����{%d� +��k��[w���a~fߕ7�6N� 	1�Y�%Y�t��3��6�=�FI�9����y<M˔����=3��7�Y�~�7Q��Ү(���K�S�ƾIRw��Md��7��H�#�g��I~G�J3x�@��,k-���>�+�������"��G���bQB��BX�<L�>`J��l��?�@�g��d�RsE:�{�>��x>G�d����]L%�y��Q�6V>@���ui���~�'&<�S�ޝ'�D;���O��O&����o>?��=QSe�YD���_�q��a�\������a���d}��K�˯�L��}<YT`�q�ۜf3W{s��m��Nn"uC�����d*!1`q�zߋ�2���f�Bj�rD!�p���12'�
�'l�Kټ��|��������+�f���i�p��^�� ��_�J�Q@����@?@X�1�������7�h�b�-�Ad��~��;��=����-�}U+#�x�P:$�(�&L�h*V�t��$�>��w;��Х��(�;���!�ݙG��.���0})2/B�P�N@�fPu��)F�B�uЂH*~�����)��C��gy��/��[�`��d���^t�j�Q����m�_0�T-�C���������G�pYYr��OՔ�R_�4&��8VsE�Cu�딊F��&5�j)���^$E�4Hd��e�݄�tI�C[?X���H _�AK����|�g01u�3f��Y��'�E�YD'�x�O�tw!����x� ���޽���m�'
}�9 �Fo�H��eSI�P��@� ��V9jbwK&��1ݝ҈K�y�&���8��H0�>���a����(�VDZ3I�EH��6��a�׫c��W�*e@G����Y����t����=+�]#���e�H����[�������㨂?�H����� ��B~���(��װ+� ))|$����.4����÷PX.�1�
ĕt-R.��`kfE��>����}��Oj.Z�^������U�NwH@���@М`s7���J�t}��P��q�~ I�۬{)b��
vp��ʀ�-�(%m��LB�9����ᗰQ��>�<j��a�&D-�Y|,H��/C7��D�]����`I�˲3�3�����Ox5CT;Tni�uQ���;�
@�<ā�>�_z,��떨��c�HvdB������`_Ҫ���v<܄r%�� ���MB��4.vq��2R���z������m�]�ȂZU�64�ع�y��s�-U�`�)�1*�0]kǶ?μcȈ�!Ca�w�x�~���1��$���ָ�kb��M6o��f_�ɫ5���?��_�cyk��>����Gɫ�߫�jʹ�4E�k�a�?�V(&� �oɢ�����/��`�kè]-�2��*�X��҇�8����\�����z9Y�c�^�|�lU���E�Sv���!�X���n�w���n�b[aH�3q9�C_!�'aথC�����5Sk�_f㏽��l�ٔ8�!���$D3rGYeb��J�8�n*f�F�<m�&	�*X�o��71�Xa}n}�OzjvvTB±���6�����7'��-�d�b��,���4Nl���� �7��e�oUxc�P�2}�#�b�������_��NU�ZJ���^���s����|���DҒ*p#ې�� ���,��J�b1��o�tV��E*��W�	i���)N�%d2�F�/��q�����ݓ�����Q�d,���Rr�#�&�p���и�^�aS ^��2 u�� ������G������~��\�I�6�@����M8P�]y�Wj6)&��+ݮ���2t��7+O��R�"1'����-�cu��P��床9���M��$+W��&Ó��Ylp}m�X�>O����@f�J�#�D6��^!���5�Q?P��n�,���t�u��M���4ţ���� �60}1{YD>W�}�f���&�G\q�� lni5���h@Pd�W������J�h�=�$�
d�=3���zV�������*��D/"��o�*>�m�OI,�>���j�-f�/�t�ˈ���D���d�#w�lB����wn���y{�������m��n>�,nޏ��R�^���Ԗ���VE��<�"����� �z��l���KK ���"t蓬�Q8nl^'h�^.�ON!6����*����z�����O"��|�wZ��;�_=c�[Ԫ�V�z�����:$�ِێ��g�
i�?v�A���~�>�-��Qs�Q?��;s�m�����@���e�����n&��ߑPE���ca�*9��V��������w���:'�㹺�qD
�}�׋V��6i�G�N����u����v2�	�����囱^�H=zqԱ?�"6z�+3�?X�#G�gF�U����y�5D�+���z�S����4AǪt}8�J.�����6�G�Y�/���$��SM�M������������F�"�$����&��R}�2�j�k�W�m����%凚�&��Q�Y�!�^v|k���
6Eps�����*�ݓ��d-�/-�BBF��0������s�ι��M �_�YkZ�(�=	�A��|�l%�������?�M
��������"Q!��O��r�����n�~�|���|�4ӛ��x]�v�:��V�����k5�!:�� �ĀAp�x�ƍ��~V��42�>d�Ǳ��){�8b�[����!��j6*�����,z	Q��o�:,c�/���js"����p�u�]�{Wxá�dg�+���=�@����ڜ���'�{\3-h�&�ǡo�ˈ�wv�:��&��ٷ
yS� M�\"�O����9b�&���}^|y=�����*�쀜"�s��pa"T�
+��/�$p��mw��Ea�7-I�Z��ܧ׬�zʲ���g%�b" �`̉�D���K~O���Vb9m�?�4�Z0�N �W�"�ƥ���P��G
 gr5�M�u�3ƃ�@�m�G�D�4r ���鵉e� X0��ۺ�Z.�s:,���I���x��`xH��@o�o׭њ�l��>�����W��K��>�b�/:�7�A� j{��u��I�,׮i˟��#Y>�A�Y�0別+!fF�C�ÿwC���|T]6V�����Չ)�5���.��F�'=?Lo�s�I�MM�X��	��Q	F>@�ޜ�H˼a��=T����VU\���m=6��G�����1�q\w�QA^�
�馊�Z���mi���3s� ��'P���*��Ӣ���6Pqn����vʕ��1�ak�[b�>�V#�2�c��g���B�5 ��g}9g[6�X���w�ϷC�f��R�I������Vn����غ�/���O� �Î��4��K���1���d�σ��^?r�T���2,�sR�&̛z���r�L6����Z�35k�_6���f�����8�@�G�y�@(��ϗ���}{�h��z�bX�-;s��Ԝ'b�_kؠԎD`�h��.���?����v��w���1a2֑�G�d�Uʣ�X��^*��٬_�ܑ��!�1�fKZ�������t�#gL�F��9��D}���8�7���<[�[���Ɏ��jh��>��&Ӫ��Z#��-|��i��4&v��!v�f�.7���H�S�
F�
�:��\�h�'x_��z�f�Ƥ���ot<�Ѫ)�^"���G�+\�"�ڧX��M��XHH�C���y��Q���m��?�r>wE`$�;L����э~4�����*L-����?7��M�A�����R������3m�T1�:�ܭF��U�}�M����7_(z��O"���S�Z�4+�d�#�]��~��s��'�HLԐ��`�G�m(X���9��o݋	�I&��Ժ�'�Q'�cu]䥨�Oy�|���ᦁ�p�G�8� +��V����NU�3;QY��nCi�i1�T����|/U�m��!vY��w��%�����;}��������!���O_
,!]�B=$�^4�!b������x���9�I��ek��u��n$�1_X2�P&C�����f||4����;�Mz��E>��!�n%�LT}	y�\x���aPu�\�v��O���x@�nY�b������� �{aUO�q��� �L&�u�y*��(�˄jC=�R{���<c�z��u��.u���]�@z�el޶Ñ�yn-:&��z�0!�������u=s���:���އz���0P{.����qF������'�kT�^�X�`�>�ߌm/EEwi���/Z��PJ]�]���H�H�&A���F͵c�\E��##Y��4�������|�F��
��q_}./�,��EN�2�O�~̬�ˣهYs�T2�ȼ�����+.|,�� '���Ѕ�`?լ�]|�<ƍ���QTG�!�k���@�:��8�����de3��m^`�sL� 41�3�P�M&��7
��1j(&/�Ua����`7�:��DOWW%�fz%C;�F�csF�PE���rŻ�~J�ap Q�ڶ��͒H����R�G��U֫*��n�1>��%��g[(F:ZS�?�vy��-ph'e��/��}8� �KWp*���2d�@Vl����(��i���Y����n�Z 1
�i�vBj����>�2�Ӓ������ه���6DcH8�U�dd�1�N ٫ÿ�U�q�t׭��7@jՅ�+� !���<>��5..�=�W��6�����ky��&:�F�q<�$�?����
��t�m���{'�mؕ��u���{z��bh���0`˽�a"���
��K/t `�|�]����-ڽOSޗ��p��!�Lm��K8��l��<�$[�30�^^����L+�.g�Sϸz�e�ɣ$i攦�d�rm����+t��4�Y:�����N����3Rn��M�7a�i�҃���A��!~���wH�᱂w�6�
�S�����EL���4r�����Kg��-Y#�$o��-�"+�%:��2��H��i�����Ń�;(R�fj��R����*A�q
}XM���  ����ƆZ�X�H�mPk����8A�w}L�5or�1�t��δ(��J݌���^$�1��閷����\Ww���O�{�g�uf.�IMJ��K��.�o��Ϛd�4�-��(����K��m��{����+?���%O{��xJ���V��w!���&�%G^2�M�M�1"r���H7�_	�h���"�Z 1��L�FN�t郏�,��
��*b��O��^6���U.߀`��;I�³��d�����,{�v�iT��`2ᥘD8��1|:V���T�5*����ꅧ�Fz���8l%�g��Kz�G>u��"h+V `Ќ�y�ܷ�.����(�J6�0U[+�NG'�y�S����4=��b� =3��s}h$g8�<Qv?`��U�	��[��m.̰�V[e0�).e�A�Do��A�E��P��o�:+s�E�͝7~�y�9p<�{@��;z�7�J]�Q)�:�C5\I�����בV���	�R��I�炖���%�<d���|p@4"g�h?��7B����y����B=@��3��*��BN��w��4$�oJX)�$$�e���8��)ͺ�}��5RkT�x����FF�:�'ܶd�1��3;�(�a���%@���9Se�PKh�$G���[���v d��!�Kr�`�]O�9<�����G֛�(b���&*�{���SEf�r�Im�o���Ò�B	�/䘋Lط5��w[�X��Z:Fw7K�@{��ytz�V�MR��3*����t �_p�!�<�i�]�ʝ�mm�3�Y�+��of	zi�������Y��ۭU�<#��@I3��-��y�sM{Xa$���N�+}�RK�S��C�~v$�в��&�#tZ� ����O��w�f4\�:�Cb���'��bny�_b7L ~�G{�<��tV�{��E����X����w1���3i0�ʫ�^����,�ͅ*l�}L}��<u؎��$�.��v�j�uTYһ�9�i�ox����D\]=�[���b�ڤ�����4��u,A��m��5^׫�Y' ���>�$Y0�������΃�����b��V�ػy��yJ>H���AL�|�@)γ�������`QL��}hѭ �KM�b_&>@@����'n�zt~�2שHEy���yw�[�G@�U�/�� _��F��Z
��Dw��[`�tNCb�4�8
(�b��[�w���D릭 ?�=��Χ���fF�k^FnB�g9�H����yǪ7������ޜ[˖��z}5�����