// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GosY70Kuj6PNUihhf8Iq0IdjHgdX0xeK1UKJk3B1YaHCqyiSAwUuZNcm8uIH2QP8XTc5L3UY0Xd1
YyVZele4N7sI+L8omOxfZTdzQF9xBAyyrXZFrWouLU89fuoAlNXbSRnbAVGqikZKqZD8ONqAvW5m
yoLHm3RBw3gAECMWjRdaOKjjzm7oXb2sGqRvEmYoEzIkHSlinaqrCP/HeYJ8uj8NIWejWdsMzkmh
Qq+EY+3swsPiORlM36hdrJ4Hz/tylRMyBqSIWHiy8qqdUMsGp6u9fmFgQhzmw/Zzz2DfHEvixLvZ
3nhO4f8aX9SKVlZXHm8FRrqUqHPhYv8NxzOZug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 144896)
jcZ+ofL/hNyihCx4HcD2N0GAvexb+ZX85lgsLgB+vWU2joctD+Iy1E2k5VuufXAxliCQ18KihaPB
8QRMXXKk+SVRxEIn5HaXxgGJae3AHTxQqiiwukSHdT7/GlPeEj9G6cAhUgYEYplGM1ieN1xax0uY
aLl+ruG2LHV6S6LP+OdbxoiSYTDcrXr6Tiz+aVmXX6pOGZSAJUFloPAjjor+BASntm9HsOJLLi7z
L64c8NFD9CxB5RUyrHPMJmWol1xvvabjPBHunUPOtN6Hi/XeUeXkTa/PGMJ2gBAls9kl0+TCQvtk
YmIZG3XnyCJrtj02zn8IHCRmBP55HBNmKU9b4HK3QGespbc4lTyNE4x6bhNERWxqW8pjexOrcvyT
5Is79EtV9kK7xtPzyzWUUZRXN1rF8MMEy8seApWg9CbKMnQHDJyTqnXGwAkP8nUSVHyp6pu5wO99
T8p8VOKkQcvsFmVyAWMFsS8bUzajjPUaL6lpsmRapektU3kb8E01gvrVLt+wCFusB98+9KixpF/k
PH/q8s0b86bwRacGGnA85CAypgD+C017PbmvTGDhLxP38NNN7QERg2gSQasdJ2D+nKtiFNksx/Rg
r9JUbUKOpAhetvmJZSbF1IrZUT0UJd4uVqNhRnEXYaCtqlyKT0RL0y7KjCzOafiFzjz79uMwljem
dxB44H06v1ODamgAsqsIMqJsv4Ivwm5yshaQxcRtqIMPl8UHBSxvQYHIG5Q5nob4IkndxVrymXT6
4wTCDkLpC8esSzUi9TMnTDPFZ9tgzRTU4kjsxmPwdz1RG0AjqpYRnKxP605sMyOGpUB6vTndR7CC
r09/6+OnNsaEBN68a6O7hQQTTt/bVTl1myq6fRjnKJXBjUvdH9Ps5guPBDNnmbqFMN+j0j1xoe67
ailP5EpPUkQOB/17pD0+X2n8YGXcvDdhXiTWI8gXyJMAZY/10VHoFewsgvC0dLvfdUljuc7WnBLI
j4yQNvDzni8tLvHBXfMq5oP8L7JDe31aJm7JRZMD3vFlpV0xhu/W72L0S+9/2g1QgRUVzl3iFAfS
iv5HNRIoHYGRkaauON51wS3nLxgjxFaCKcjGQ30LG2WfktzPq6Fjm8inK+DQDb6iuXjm+c11L77G
glNkH+/Ktu7WMzasFcZV0CF7W+AHC4mAgLZKMPTUWQT0CIFFwiifesWL8RPGhoMdKpauN/lNSBmU
2WHiN7YmvQ7X2/X2NOlSqbjdJ1M5+vgAMQGyrmi0Pbj+h+niHqF2n0Lm+0ckQZUkwUNI9qs+1/kU
PqwvVzNBdLppqonV9+oH1Ew2/GW+GSN5a/q5zbkgbPS3A1Ejfi47Qp2m5/C898zmuXC7O3wYaYHf
+371oGDVcgcI9ewpAvvzip6XKoPJc7PLGtTxmdhIJALuU14BWej9YE+U5wpPgsYxxh4eGiARV+F3
tCZEsw3bQh+rd9keom/WeUvbmoAvLUP3DUIEaA6h9U44lrBTWflk7A5F66WHZu84xSesne/JyO94
7+k0DymRNllJeVGAfuFluXgDuion5rUQQbHuKt3RdCDw73elHO0w5lL4Q580Ult38QBUNLbwCR48
fmddvD9cQVKnGXVZDBvjX1xtk0M9FZ+OhuD63y13OjyTSQuvr782+K7b49pxit7dWFgT3oKc+IYc
X/YKR0KOR/ztoLONc9xZPjCYk0PL2YaQyyHUsiVQV6+rrytCBeL4GCbbzdau/xgPm4RTHf7jEqAz
MAFOY2cROlZCmjTPvcct3sRWUd+4GlfR2Xn5wfqxhvYFfb8Jph1NL+IXbFlEr66k5vcLANPasMqq
zNziIxJZzDFrmz2GH1Ugl3R0Ta/Ic6ouM6SpvG7erlRYGKF2ijrWBvj5V/jgOQYwnCmVyXRkBH+a
LtrUpXy+W5FbuAKpYI8ymAExFN5hELgYjU/4bpWOpoOUG41aTQVkhXBaRK6mx0rHEAQVaWT1kTiH
YD20bJqkl3T1VQZvDnsgJzraUrgSIGZOH1iosqPGON/uIae3OWL14/db5+mRfSRbXExYDnDcd/zx
Vv1mAmziqdWrT0Wf27wPAvZhSXeE9CR3kkxe6qWfuxJLuC3OEX8PT2yc5Ktwpnfh2vejHJcr6dQe
9cYlS2q46ZkJ6vJBHR8ynaDxRTMOlBOb88gbyv6M/BBbUpMr1BKZg6reTed3k84yN40BjpojTEUi
13S5DVCGEP4PeNpyFNqcbzEO/azNsyeaVs5T3Zverzzw8CESo76CrYY0gVU1haCiBAhl2rA6nEmL
TJoWCySN37xgfHVpkoUAHIErqUyLhq8fxXt9peIBODOqXv8aViLtuKTzQPNIf4tqtjiMK5/5ITCm
4IOiDy1qPtSmmhxFr9U8GtM6pwUIoR9ZjXdx5LzP+dGiPGFXJy2UfADK54QvHzRSpzJsn+5v+tEI
rbDOVs3mbpA2PC25EvSNA3lFYvp3pWXYOyhxDEffBHUoKKucd+sVhNvWfm5d6drj7KX+qJcYX2JQ
ixpEi/biSx1mo2tRKmeIS0AmXALmnvyLkfHaDSr8PnrtFo9vX/iQiK784lOAYG8LxE8fW7kwV+rY
xKgMZhn26iuECDqW0nQlvfnQmPoPbti7/yn7xY6OQGjbZYOdYpwFjMDEUnVqiMwVd8wT5v1pY8tq
qVCbirlwyW+jl5skhSpQqfSiudQCnYdyf+GWFgBAC7hPfQ3ZNdicng9GVeb9QsRQTFRmBoFJDKZR
U7z4pkLDeFSuSOZn00DCdGw2FDfOyO6v3hm6PgI4QKOSBZX8G9EXLmLbEYC3UYmWJrEu7I/3cMCF
eSjQ3cyWgBoNRmSRLC6mmGXrKV3KtpDlRCNdbNOLv23itR8NoPHCNJKPZadlB//RcQcyHcgZYu6M
RgkpHhaTksdfcY0ATgjf9rw/XWieueHznGX8dha+jgFEmDSaNoyAHyD6KgVi8yPQX8KuIDAdt4/N
/fLQXISC18YdNMG15aAoZ3MamdJUbuGNf9dHcDynlMYrt9FYVYzgX67nWQb4mulI/bsTldEUR818
VjZDuoJe4Kij3A9Xz9Iedew+7TlbwMgrjIazP1FDJNPmHDuGhlXfsJ6tRaSb471Negi29/OZJzb5
FnOJ5cxBF5X5XJyCC5FPTN7PbTTlRsYctwq3TwmDBH5ua1VFUtuEfGCe/ZdxusbG768eeI9x3U1s
BTa8nsYTLme694+lA7gk0RF5Q0TCXBD1FqVBG8/WxyZj80co+fehvSXGCeaLZj9hpfSbpEmbznpz
EVUkZCBS7qaMDc8uQSJBuUTWHqNAAl5QPyZqHUWdwpBhb3yVgX9c30PgJYkNmcgpQvHCwa7oK6RA
E4lBzp+y2+pi8LW9iyhPirsJ2XPTgASbMFuZhiJ8CgIFHpqndd8qVS2T4Pz+0sc1XLMZA7aNF2TM
IwZAdsK7IaGoeG6NFU8VcQkjWpyDxDHLEALXUgBJbJ2IdgEg01hZT+W+lim2rVqsgbll/BhB7jmk
8hGzCO5Ov2llpM1LexHGlwkPdUP5LhCN0Wnf8Go7JkPnMc3YEjcT48e8XpGO7b9sd6OVmC1Z5Ee2
ep5n1DRLsIUIBVZqoq1wIDobTiuGMgekJCU/DrrmF0OG56HYLNMzeJ7BZ8K6MChNx6OifUD0e0YS
s7yAiZrUkoXa6w3FDB/oWjzusT6WlepaTg4fceU4FND+Ccdxn/xgSEZ2EbCF1fxQX9w/QuiY5A8f
8pyRYgtdq7YMUlf0776z7b3hVPQ6hgXI7Xy5GdYhLaxnnXdxmTlzA+R84LtkOfay51LW3eX6Ik78
mDBNOJCIIpv4cD8fP7Gt/KX5Cj+RKV/WB8KSibwGIkGdYrLVH3+yEbj1mPaQZMXi65oppiCw6vIf
+oDVDrnsSiVuyKeAuE89jHRr9GAhxSl3Wdl9kmzvKgWl+OOxJY9udheEzmjrTpnSlpcDm+DaiYbZ
4MPcFjs+tVu2zm6Xe2xdBrLiqaoL1iF0jHoFtLoSmGhEnb7decQb9JCx5Tj8+bSbJmTwWdyJsKz0
9y+uW7csnsgp2tD067SVNPIUegoXrodK3JVDzrGMnTlQHPYAw+KOLfobJqViSKOBiaKcgCqEbwlm
SSsowJOjeOhUKtKgxX+hSxZg1AQzmysN52Cr7ph0Sh1Ci/cPRewTi8HbuDKR5GjUBN0+7JJN0cBL
wxo/4etg/NDHoz3vVmn8ziHaN8aZrdrYYZIsf55QoZqS+ZdEnFrhxFVsiFXkaeE3eD2mlWZtK9ww
qS6nJTvPCKtiM7re1zMLND2TCzXfLD+i2L36bDVTC4lKltsbueQ4Dfaih9Wk1fgqP7iyQDMfgaBj
J1/xSHH2hUo4cVIaSPXoDyM66TpMdyzJ04I/LTr28lDjuPOrlVKiI095EJ0lHuulp2uDuS1WNTOd
CN2nJ6P8oqrztWdziMTZyNJ9ZsXlZE7Yyh6Qg4b8qAkr7dbpLBkwC5Z1a+2QcqlH5I79Tnl6XG8E
zTtC0xi7hFlA/L021z/iBSjAgmg6rPP/ejMIuixPs8KWBOJsDlyqiSgpjzeMBndd4VxH3QydHGuV
Q5k+RJxjGTmZ5eRqNxUJiHrRwMvDKC74T7oNfoVSi1oVabrjVuyIpvkiQLZtsFVVFZ3tDsyJ9hbL
Q3Ghpd60SPfIFJTUwWJC2IeRgixQ+ADqO6a8FYAOD222YluQfWVOSwGfSkZhTwsaIEeo2chWySF6
VHVlZLj4Kf8dkmVWpRO4XMjP+eMKxC0nLNa5PtBvdXuuYN7Yfni8Itn0nreqw2DPyU8qvQeh5SjH
qdNeuzOgfiLrLF2TYPdgskTTFaTzQwb6bwZUJmO8vqWAaI/6loaQv2CM23WbGkCEyHsZbsm/tETM
YiZRq9UpmO8S5eqfwnxBV3pKdQzkwz8HLby+/LOh4cWPMTfZfLOg9hxDz2HR++gwJKRlAksyBB8Q
QcrPtcdiA2II6XuX82hrPXlEU1EusLV2bnQUfv91Yi9Bz4QTy0v2HyEO5Wcdz2lMJEeJsWFVE8a+
Q82wEQ5x98saBZ9QLX0/cN3Pg44aMtPD31dXkFFu07VFnPX1JwUXSjuLv0dsLIfTftIUQF6mtqX5
xxS+Z5VBmoDl6VQKeu6j0kynMKx29HacyZwZgzDP3vDjH3+hEhNYh8ZrAUBRljHFd7PBBYbnjDca
h4LXnO1eMmtABnJITvcCVfphekK9nuLpvczNf1Fq1Yy7epsfYhzsxyUchsTwK2zCOAowovDC63Mf
IrbxmN1hW0MVcpxB1hi5+kscaKBy808X0nvaeHmA7JcA8WI9t4qfKroEg5Wy1uYScZMGe/VkLxVt
9Bu8gwqd8za/LkgZG8oFXNrAhlXbS36mUzM+WmzF+AJVsSL8lFkrAVlMTUwPNzWDjBvtjs9eBpQg
QB8pWGueyNqJLf5j5c3j1IFu56w4J3w//cbeaVzdAGGYUJZw7PiswMjJrn5c3XrF+WOk8oyLdK2g
HbjS3cS9cXMZ5jYI+TFxFfmEi+q/ABg1SCyFIofpncGk+0cuuTh60q8pqNaOOT8c730qy2Rley9Q
/TCkPCcr+OBcHaaZyiij/nHlW8+DvY+EgSEIjWOv2eiepjKutrDUlh31WKDIRAjNiZETEbwfzfcp
B62G6ASAbPRb6GQSmHbh/KNPMVVZSxcwjQUY/T9/9Jdps/NC3JHF3WZOt0Pfs0rXiTJ5DIO5YyZC
FnJePMCstyh1J9KTyiSojmgP9a01n5W0W0Mc/TbNO0/JwNhPD4hYZR2eK6GwaC46uOxbVomgJ3+B
W2u/tNt4p8LDIZAic4ftQhZo/vdPAXiUoHvnR6sgk6yx092XT8XHBFlCsmr4WoaKbNkFLcAwffOY
CshalsbT2y6mkAiYpfh/V7WthAwemdXiN/U8HaDBKSfms79tiXhUmjCLaThRX60Fq1ieK8+3kW5V
QJtcqdk29PmVBZW9YDNQRZnjRFE7AUdmwoAm2cTyLnais7he/oH2CHSLAOnDXPWH/wHPj45kvQ1A
BfmcSoFVs5VsOFyKzSuMf+fbuStG4xnylorEPfX+PMcOFgMUkJKlFEcYJq0pgqq3WoXmF5yHb//1
cwmR8GHbMImGShsrlGZnlIfpyLH9CoOsf+kA/TfnGmHZGGAjMTiYXfPLG9qPETePiIPGCpkp4Sr8
6IQTY5peWOTzqwfdNpCHUCbCJaSxLTAeBJPGYx/rvW4dukM26vZ0HGmQGVANMyPM7+Indg/7tEQG
7dR6OHvZS5KSSDs1jYhnctwzUfTLbvXINeosxVu2LBUxvTHD9qRV3K5WhZ4i9MLrYN5txheomUFn
RpmQ/UR5py0XT1Ihr8nLioqro1lIVItw9Tkb/2zhPbPK31LrtkLi257skgugma8S7rImIEHuT1/m
oNyWGdUypFZxQVWIFpBAV8LSlQit/aad5inPfmu+bacyEre56X/Dk70bLia6ti1OxYmq73zMDoTJ
8RXCsBDkNVNq+zFczrrj1ccHLphvdEoe0HRDwEOXyZlaPig/ESkoPpKaxX8EGrlWYfq7z593mTKw
HZzKGf2rfkBRKpb115tRfhcdTVXuV/DdUI1Dq2BhbJKVP92DKBAkmfp0jX8xJ102/P8I4Z2XgI3r
+Sbszps7O3DPrOMNPUFuE93kITS0odoQhtROUOJcaAkRmZzp64Onazot1Iem+mM6X7/5QwwaqbbF
epwrBsID0EVPF9HosOWve6T8SYk7Y+oHynZLPQgbALlXoXsutYsrvVnk6x9B7ncds3IfnXj6ZsAH
1rLkkPD5RPyvj1fiaiS6qrpNNxZFmLEFNuSfuSP8MKBAp2jNdkVpIFzr3o8uhgcGKeKHon0s8NIb
2xXMBYizr3YtfCbz25O2pAZQJ7GnWwt9xLKV7P20w1rMXlxbvg0qH1s9vhn/rayk6tmkpyoqMyR6
JyO6AVko0qklvNUPZ9dVKo/enT7Zr3VWNFOMQc5aw1xXozUL0eRKiGZWuaXLr9uaiNismGSjbIlD
mNpueysstdlJYLWL+J0GJPuOiS77Ka5/YxxDGiagI9e0pWYa4H6R0KNM+vXtamCkPlXm16vPldjZ
/9K9wg8iuszcuBhoj/JD8kp08GG2uowwrkG48Qia1YnJdNQEwMnG4vQLx3WDLgGqzozeUcOWBp5/
LRppmyH/P4xX8tnly312ivcTcnncqHPnt4eJpuOHvgOFDFb23vY7pJBIFZq1EfuvyjCvAxV/Q3A+
UOBKNu4sHHyY1ERREOdC/Bve34IFf8nRUVRnmNVbJhCfjD99G4nVFu5VIbh+9OsZawdLWAjGJPBh
V0iJ9SqHQ/GOuIRPtzri4k5cioHakLdqEQvejeguikV6hs5wCaRpaD8n5BsIXhslIrGVE08otWHQ
j/MV/bZRB/DH507EtVgU4gDN88WS6KwVZwkzp05ApEJmSDSDls272FBwwKex+0rldyZkIWClRw95
nDheVSu9mE0ZYB5gDAQDtWqKFhPmLawOe2F0TgDDeMUIfYToO3pYY2vbY+Oxdqbgjyb5zmGQSBy4
TI0K34pd7iVq0pSVjLzImrzWCSgUgKo5h/VniccBbP5HlHaHUJs5aClR4Zo5WGseXbCHWewrxMJw
TIa5BTlMfb6oXwVt60+P8mLA/h//rg4mAzEeiQSdA9U8AtbfcSNnjCxjbJPoAojvUVzi+CAvmbWS
Ev96VkpG84VFFY0yRvRYEpFkcRGsZprpqRhsxFz1My8x3PEwVx/z9gvgPZEQZHyBZMYDgmtDpCbE
UP4+XzrOHZUPxT2A5FXgHujSKt4feeSod4vX7h3fDqmOBwiAmo+EbatX1w91bIu06+/Cn+1sgWZy
r+8ai/kg5GRzrS6lUvTcV4qclWE3tVvgx5NLyvbR+CDYpnsgT2o1MSg+CRSQow6b3JK+NpToT1HD
fUQdebmuYeLCYqMW+moBSlu/ztODnbJAAe6hAn/a49W9MCWVJh3PHYje/kNZw3xpDUN0dE2V3Ccs
Yf5KaU2p7MXqJ65MKG5/odykaZR8EIyRs8DayMbgCY/kB+6O6NEWPQidLpMMOj3EU0YrtF634+dz
pnF+5vUSiUzI9xTQaNBh6/KWNf5HuvLlJrPey7P1C+qnsOwfrev/zeTNxufPlBu3KvQRr9CAWzkX
MNdkjVOX550b2vwI6/q0On7d10GQxGDQL80CzWoC/PIJnewu3eaj6kaL4WLCbvn5NgZP49+3mGvv
RK0i/U5lyE/Zbne0a+ifj1v6JLygrjEIfIUHcWENckMrl5jXxxMRNOP2ziZq7XADwMkCGgoPxyBQ
VMyK2D9TlSrxi35EVhf0Nuzk8jma0JaB7IpgeyC++oTIxuwTa4pt+V13P9QeUMYXHF+2zaFRyWc6
wmfWrtqag0+7Ek6tDHRFfF3v1Y87twjS/9+KyS27WIIGUcV2fxEmAb6SEEOWfW0NP/Zk/m9fW3Jk
Gw8Bu/8p6XRvGMU0nlKR9lewBhMnDGtmkE/II6CfS+nKAiEarj4N4U5O69cRZM6YvGRBPUcCPfSn
8w6QnfMl9oiNsUn7L+Kqg7kWQfYBaBgJN0flA2Qac8oUo1ZF96eVCUTjLt9kmzYjmIKNtNL/guFX
49F4Q7cZBPBrLYxjsOgzSCEOYYpLWkyd/FezpXHOW8enso/ma5C3LwIJAxaXz/URh8o0w+H3S0ia
T12KoYAYL/lL9Albb7iZ/rzCHPI/YNMN0OYE9qzCuSXOipKLLli0nv1QZoOPqbRqHP6ygGf1qy1v
rAsHUysqCaUTephCvITfDkckMfi/ktFvaKAwlRIq7PLR2CBvp5qCGkokjXsMgUF/r92M22PCd0Jc
zqvZ0yYid+HYZJd2IiTGHq3ldEXh+02R6zK4S9ATJfOgMD4/Q34Nu94Y8p6MO4zcu5QFazAScML/
Hdn9Le0/ovLNJ4iiJLW/fBZwTkb3GeUoBU47eJU1rcXP8c+3bm7IhqPeLkX4waQvLHZHvNguZY5V
Z1sHXz+mTMoyzu5jWj1Np04xW1uxG2b2GVkrdO5JWEDkfckWk1GE+7MQ5MdMRI2FLRnWdixxtgb7
YeaHEdchVW9kwo8wYWkzakQ6Ditxps81jGkCQT+3hnhzmRAXTQEOnE5Vo7/MSccRA1EEolZqYfzC
YXHG5SmHVNwB6bFlpaL7U9Wh2Sx54ZyNNIoESvVR6BaI9XGgCKTWl4YGATQFZ2HlkRYQRO6xyvyY
jdJJmeY3vsaXKX83FBP9RHInIWWW6HoDoTrYuWpQq8Vh7uDTwKgiaB+4UVtt297W1woGENmosFvw
PAtsCYfYm8CnhWnNTXVYTxKBVi4svIK1TfIkWdFMzkdlkhcMScygqPcnMO9P3EPTwhLcw3LAfxgr
DSjpc69XdxYehRpqh1rG8atTxPhDS4CeTMQguUdxbxGSeyRFUBIT/KA0SWwmzZ7MrWtz7lsP2jhC
uNsqwao6lszxkeYZwdS7X5YAoO+tUxnjCrsOsTw/3OtgXq/ADYQPODRRyR/bx6DKXu+2cfHrESnf
MWpjeHHtJTUYum7Y9rSOOLgWod0ZGk+Ky5hHTjfoayfK/AnixVCuHShXV/OhFsGqgshrrr6OY230
G/ZHE8XRG0A/xarqxun8RGOpMTCDqcAV9SNuuI7WSvCaHr6ZTeQfWtfZX+BVmiSrFvaVq81GLkY5
soVNi1yBJw5qcxYUzBTVfaBQ0IXu/7NPiYXJQqAHSpW9r4DM3fwYdGoGNJj6/9JBHz1++IBI3CYx
Qs8O+K0xy7fzB4DCsns1/Z6AmQRbbD7a/xGiB25qoqdv3OFyTkRl0auakeBNfbalsTtMFW6ZE5ZI
EhSJ8swwuUCHOVxhnInWFQRMAYxRoITTalukoe+2pDqKqVSER9l7CC5xIF16FS6+9uOQnEuKbU35
5TbR6q9W9GoOK2l/HQG9x07Dkh8zmxV1kJ32Cn6vlfFOJez1GzWbeedK1wpCgVP4O1RwxG7K0m5P
rPZVrHLYAl3ix3IZ+9o/VeFtR1oBdbgqXbJgFz2gCi61twSFwR2juKsuAXTFRbJ+dpqSToR4iwlI
+6c/7tSwjTBzMxLAlW9M1AdEAswwKrPpLKLNsE92A6XlS8xMGg9fQnpU3SSY5HhTKxau78oBMAqM
9duDdyfwobVfe8rAxaQamzFfyMqhIPBc0Xwjl6K8i1cgUf+wwHXHuhU0H3NNmo1SSLbY3xuAwvRx
9jpcuc6tFlv9gwWIyhD6/xSoG711EjqK3J6uoWZQfk8aPFhubOKYpR6McTRYDuqwBVCEetx3l4Bl
dLEPUk3oqG0/FXAq7oLd9AeM0so02X/6pJbZImU7i9lN/mWosan1Tpd1Hro+TzZLcq0u8I5/yHIt
9icx5dx7sdI5V9KEr9wFE+URmJL7OhsDGtQG75ZfOJI7vCLXwauEdUuUX41qyku+2YT0zh0Tmp9V
c4YIXzL7JRhATdXlex0OojNzyqrMLSVnfmFGZh4n2uWbjfcQHm/iOSikyUu5TRxALWJiNIUc4Tu5
B+plhvuSzw1YnoPKaYriGc5aKJX3afFeXkLJ/2Fm5fcVFIPxypJI2ViSJI+2oGrj36JRt8PJalOA
/YHspv8xwniqVNvK0ed+anQ2IEg4Hd0ZJCRfKHk/qV6xQzC5QJXfyHB0AMH3jb9TMXq5uY0+7TwU
FUt3av1vSJohY9r2z8zYr5XXY1nC4PuZ58BCi1nqc2u4XZE+46yvqTG6LjQY67NHwNujgl8/GJ+x
0OwpFHTxLi4kIGyiE0ua8Vl+nFzTggXmjm0iFsjxbxSrSY7c2I4Z3C+57s6XWNDGrPe/l3ymR8Ys
GqW8+UShvWOJLDv/70tX9qivJrXhmS3R/v+HIRl31SImYiCqh5nBE6YHe93BDqNqhSsQn0UZB+6a
0tJFvveTGk5kXV2mElhqSc1apdNoZih8gUoS7CE57Jg1I0JJ0mM6G/WvH1NrRd9bOucK2OEE7vMx
MsIot2J6bupqHKbz83+t5B9BMlmwATVQ9+rs8itHfzsXGOpkZT2IThBCBaztNSZmjKbHq3dEE7Jm
+poO0qMs0LomfTaW/0RVow8wnJDSH/Lf5/YJ+WHHeCo9fQZVOj3pf4rxdgVSpXt99Y8jbvUXCCFq
VnDhFJB40pl0t/k80jxXxjiNE23AN6K+3QXs6GSxQBveq6kZGfjAKvvBWk3m2UqD2bDA041TIQWC
YAHKe7SbDUPwcA822fqPYgBIQPT12Edpz+qpQU/YflzZvhxIo7whtnqoxkhA59aONiTtLz4gDXZx
FIM2AGsNfx2b21OlUCoCFER1fhCh5DEd14irmpavydmENNvmn+/F6y74PaCI0Ot+CaZz/KOcE2fc
DCw/RMGd79hBcPTxaNbduSaU1c9xjESTMoJoALE1yu8blYb/Uu858n9V0Jswwe4BfJtcKXL8p8uT
72pwEhf3uzp8FE/8VrgV/bEMmvABgD3RpTLeM7TS12bFt6brdZzo1cdbLjDBVHg2kQEBvNrOOX4q
3+2HViZxFN9mHShKBaFcios/k8U3pWwIK9oJj4Cs91mJNYroiwzWbQDUYXnzylcm5CnDBbGoftRw
5ruv7OWQPOQ2Ei0ndVSqQkmqY0W+/3KOO2nu2rcDeBvDTJTpwmsg3F7ZovV7Whll8obLAMDovFM3
8h3ENYQSSnfFMFpuMlOGmvnwfVvqfvJrNUgb61QC3Goai97T2HeZvzNEiSP7NEF/SJO3sN3+qRxU
L2Ye7lwwBkoEOh/BnfCm4RLdo10zDOVJApzZHCfBEwjEU3CrCuJrhp0BAneLZ4Tw3K/V4ayFDZ7Z
mEzyL7Gjs5moKuwUoitGr5StceBSNmhhPVQfx7mQF3olIGyZ5n/fZMWKe6tstIQMRdejKfsfk7pH
+Xy27ZxchwAq7sWU3gSQ16uSAMxrYpJJHSWeM2LHKkp87bLIgsO6PVzzk+ngbCWXTvlr8bn6RE0z
X9OvUr5hpp1Y+TCFTD6YSxGWLyTS8rcXVggtwbVgOSzJnKIGiht1tbHuuD35NIibFF3DCRarM0Z/
tu2hHRKsd6hkIsuolKzPIFMANLxDED9HbW7BxiwzYo4GTgRHxBw2SEKl+RMGWD9N16gdS88nv9fd
d8I7fJpKm3A0fnJqONHEA5oGQlV5yTvkadAJBl2A5LlDHigRZKA2sGq6ZZFHLXf/o1UfFpilFtNe
NK9deIw7AFS5YZ9qBLWg5EQcq6OTd3UN/UM0mkywX2YJRAyDYrbfy5U5+QZH3vlHnXXk1nZzcrVX
Cg4y+w/LfAOc0DSPPuitwTzDmD6f03Cy/0byujjAx75eDM7bxduPdIr5IhqvQ+ol/nTqPmJTkXty
Z4ZlG5TbwISkCwrwTRFkdSHoXvfP1vLlANKYVmJHkKTOfNdU95QOK/pq8oBoWe7kMKRTHZ/X/ptA
uWW8g0hEa31jEVZJWVKS3aIsyGzqJhKhXcS1hLrTAd9oA2XbJl5khxYwvLOL4PkQP6G33GPCVTlN
YoFN8JUKG1c3gqVIkgebX7BGafh+OxuRTGsmJg3glqaFWpgWGHG2ghXKzkkOqgIRCW2NnxeHpVpV
YjOuW8RXXmobyj9l1rg9wA/Umq83k4ULQmWCZU7Rihs+jTweBO9mQbqJjNLPTI12tNRjPRLJr7+6
FWSq3Y5CLNb09wxAglcXkw56v0KtVtJ1r/WpECy8tFDlArImx4Bq1UX+npR2N629pX8rx+Ht/K81
045gw4Yv3VUxtM+6hFf4+BKIzz1tGitDto4PefVlrkAUELK4wY4Rgn9Ip073Of+xVmMQFh9vPzKT
vTEEWXYSMYYWrshlx8MQ35ZXfiKQ7P/J25TLoU24SDcl17pNCQJXWOSVJtlxXzfEjXrVl1v4ZBCM
tGc9fZypP5Mbufzo8JUweuU9v/S5OFcPrwcrQ5jZSAhriNz6AfkKHyFUGx4JODr7wUzOJWXWbhBt
ljO9giFldFqdJ8IIRMQ0si5m/EaJSlk+ZWveo48TyYFWfED9GJwpd9WPDZzenDm/XaforbvhaWvc
7eaZEx6mwTp4XMY33BlApeAjFxi/0Dbr87MMc8qFRvu/EGwGueZTrjhVu2UE1D6SKdryyXDVFyPw
IP2ehuvozSKVmGUawQrB+bVXF60wgvTseCWwWYmePQud90Fchl9Ackd7WEr7opfAc+lFkeLt4Y/Q
QqPS1RiskKyAznO8kPe7s7mNJzYQd5izbH7pWquMlBmdi7ve9WdfVrZbJbs5BYny/EEbVXzsHgwt
ZYpLtv8gsHR7M3bDnyGpmEaKS9jCCd2St7QE84oENDhMN9q9B6YiaYnzgPQ4ldpM6jkhSL6O9f3F
0EWfcLmNeBQ/quRma1qwmoycnsLk0OWYnAmSeUOaGHIcL1T7VoMXqB3gRZkRxPitPni7gYSf06wA
jDzhMfntmuA34AIVzSDiEbRh8m+J0mxKAPtQdGY8gdNJKqiNbwsjGlr3Y141iP4dxnTdKGKinciZ
paQ0bXmqJadiDQNuZUse231B7AFTiYg1BZWFQmfgT2VzDMkwAldukyzkOgx+qzjZpSr2J5XzPQTR
sVpo6YGpGV3rY9ScnMNeOyC0hzFv22gfp/OK3Trs17mmJ+XiyBQgT7HxybfYMGIRzFvyK5bbwffM
d4zH/xi0EESzAJdbehXwH9xf9M3VTqr/Lr8IqYD7WvFlchlrLBaLi1fBYuFB6PCTRU2vrnw21mz7
F5bYnY4pV+kkDaPtMw9XkUrKp1dqbVcvCqnTar3ddAZUSuTL2/gDSBR21CI2ovruIl1A5Mq/XDQD
+TPqu9zJ9b0LANCsvRIb2iYqdatVNnfYWQrNZbysZJqa9X/Few/JIHaQEALqDADxvweCldGbRqlT
OSjc1ofmTZnxVpNgIdXq15+4fQZByeg7BIiZKtIUkI53M0noqn40/c4ghIlWyTB/lpg0nsrQmcyp
TGAaZ9GrLm1dGYLotWJqPA2qoYQIFhP7csaBNhiYEILVg/VEhGMwkWZe1Ivrmw9ZXSaljsYpImyz
WI+0qPKIAGU6xo8Jgrrtj7FLb/efSf4sdpJ/9QFa2zbRykj6/s99L29EIl37Dy2pgkjykcPGZNzm
jWDJifeWqxH3XIgqCGXmV9wfaG6Pk9YRjKyJ9Fn6vkFY1UqKSqT9zojqm/a/x8Xn5cHvyU0C5iHC
4wTt5FZcehyvxRX3OYPfKM92qrCLXCtI/b7Pji/RSs+FoANqvGqxW5oQAf6FS5Q4DtLXAxtDFoXv
t2MKdnWSyaUiBnbpmvR/0UxctPXljKmWa5GzjjP8S+0DjZsjroQC9xdpN0Sj+0xbRjKemXggIFqv
Hv1GuVuBMgeLd1b5xzgJ3lAEBGT8vYtqqXvPcpntybVYNMAzXRaQ7hFmXFaVWhw3FRefpKQLrzej
CDUw7RlZVOIr43x3FKgGtOZgubBXtQwXAcCnQ+DjP5m3dLsTfi7vMRT3ZO6skINsL0GWGKDEx2sN
4EURNv4ajZvCN9yEEMESzvYiXYcmSu0dxBcrSBAlU78XHwLdWKVrYcBRowbFtJ+xU+14Co81bfIb
EboCL/wwzy7OSPBgQuEvi/L3pDDTiqDVLAR6hdhPXKCV2eXVX7xUb8/2aT1m7otImW4rvO4RhQxm
b4XXxBE7ofg6Qf6qJo352pt+ET1qfF7SttQTLEbQJtt2UPeDJhSsgdYL23zLj5X9rbgRerXuB2+j
H+OOFewMDC/pOIXyWEllcHEU6l+DL8/vCh8twf1/t3BmuBnWrENRleGhT20Q8wdxOxpxF8M7vIDy
O0FaMKZ2p4+i2DhmD/atZ3q5VcP+c9z9TOo43rYW5abYtWMqLaAKTNopQAvTvmts8AJ0bAFkaf75
IU0G6IbJ5JRSk4t2zzCxPmaswtkdxFIaZSTuAPlwh2I0naCvBjUmGWfVklg21OSD5flFE2O67ieZ
6fGgKaKi6jp5V+vGmNMtXDrDXGbVLKxX7CnpfbCH6+JX3sfMLFLGlKqAYCqML23JGgYS415bDEKG
zazkrVqW4H2Rl9SmnEsuAOFmdnsI8Q+Lt6arEhToVZZB8AflgNDfR9V2kN3M0xL8FkRnZIvlDpky
6yYniI/6Ctg1Vc3/nwBWF+NV65k19nQQWKZrqVJUVAr192pJhIvqrH18KFvRxtF2SNV325HNjeZE
/KPYHuK07Dzw2pLJu/vRdoExzpQSwh8BNT4p3ub08Wa/owCHSXiy4aNRUyAi/7vXHr/vEXPcdG2c
xFd4XsXhEk6/hjvQmJgdimeILgQkwtq1xWMrHLb6kaouRWhRQMkfdfmoH5fXkvj43O3VoDZ9q6Qb
unBMXCnFKyxvyEfPEwtLM/LM5n+sTnhD/QSyb9TbXNV3rCfLz0jTD+jf3r2LQlvPPSqWY/ppYPQv
zMW7UJHCzt/16SpOw0o3QX+/vpmTePtFVZ3NKse9XJnsg4BCEL+5+7KD5tNkHllTOax03zkzQobV
5LkcpCOfSRFFUgpmhKmxkWnCK6A1gamzqM9zodCLqotPMNq/KZlWIBtusLR279ihnqbt+YvoYfN4
CxgJJscdPfRsvMxGN5c8m+aANujHr064OburWyvDJBs7sLAucINTn4n1c0mtJztjRFD3BvKwAciU
cIYv6jBuYIVn+VFjt9WssBgDaCbi4NOEYxEa/cUZmwLLkfQnh1dFy64Jh5Awj4PNuLV8w5jmSxlL
YjxXq9YtM+MCv+HK4pE89/xmGgiekj9TI7Bf2VAn6y09LC+CdEjYqY3hOU+FUnBFThdlpbIsaktx
QV7Ig0y+KD/5KeUi1YzmizUoHlPTyt85EoWnyTNxxuxFlGlTJRHy6c5B0rIWAIGLjLlPbTUWH0Vc
Mafy7bh5ptkyMwQCWsOXH32Q+D5Rmr5inBEUPEcTmi677SKjHqu0qvlbPLMO5ptXXySnPqJ1fUjv
d0YdFNznUzw1/3aZ9IK5hS0RfEMrrJ3eVfP3cz7N6Dw0eYfRGhp0pui/r+aDVHm2BH9nD+gFgyfQ
YBh3qI7EjB1tqdLYbiR50C3xO2nP5ntnfpcR94bEjwlGJEIOEFGl8VkLMdsblm7eIBfGxzUVR/Fu
3Z6jT+Uqdrj0Wko9dsCZFMI4dZC4hn9TTh3N9Cz4kdF107jJ3uR0JvF8VfnG58TQALTydc1SUngy
cz++zrzf1dAOi2QSpDhsNnvMMmnVR8wY//TjwyYkf+M7PpWkpZgYcUGw5p1V6jjlrcuFAAAwlH/x
8VSzw425odjjzC7pdxd8sOZJLoFO7bD6wK2djwnM52DUp3/WMEPunW/HjTDE/wPbb+FZs+/IW1Gf
vN58vDkqwEmo5CNEb8iOG3z1rBt2eYE4Pur7i1vrjqXSjR5KRaIO1ndvu6yWwnoV7oitKlb8Ulky
MdKw1QT2o8W0MIfWXnxYiPmpH+NRIaigdnH+VkCLxKAz0MKc76GjSM/RWaTH8v/3WZqoyXm8f9QW
lx95WCedpdlJv9EScdYd4H79IB3gPBCcDogxuqoXHSMYog5TvOouPYnd1xQmMG7yWLGF+gd1HdDp
o/yIng88Oc6iDGnuJ8ydGjfNIc0nI2+mwupTlZlTTZSiQF7Mk8PB7OAISnoslhLJhqERERdVp/eo
j1LzcBrQpXIN6lGlN1n8MJKWiG0N8DzVW7FVGUTAOqkW9tbi+4xZiwZYjp7M9QkBrSHull5xpCOc
kcbWLKYkSp44kJhlLO+Jn+U1pBbSYGeKpj6Li2H6Vd3RJ3n/9Bwm5tAvuThwQMUayD2LGFttfTk1
Ikp+QDRVgtdjMkNNPGMEvvGZTpo4raz4xim+gOWkoRubGi0X2bYulfLfqI+7DcUXSN4rkoUIkLSn
hhNJDushD5s+kjMIZ4+6V8rI+WOS53ndsED83kQx6I4lCqVlOLeBkuJ01A5WG/R/U9LyKV6wPscQ
M6HbvchlJ/IgBntmuBVlhC/qaZVic5yEJLWMN81dHZF3qOwbW4EnYnCsh9IV2AI34syo9njzBA5N
fo46aCvSClQdHgqG3CbBjz3r0UJTDVp8yu/mjUATofS5K3zIUi9UiXGmLQ9E/VM5OcbxfvBNDgs/
nf/oyVfoA6Yom3992KN1OtFFerksuw8laFQ6BHXphvjGePRCqABM5ToEqGAPNZBqKzqrRt6UHzZY
RQp68SfRAHIkPWnXwzZ2MyDgyeO3h9QFeQrdztNrxVCPoX3LzK1sVx4Y89057Z1wYfrfchofXJYS
x4n/gePLHGzmfkTXIt2ejAOjDIU0+IY87kTkC3IDoaiiQpV1hKs4y4rW0spgOeVd6YNdV/ja3leP
BmHI7bqPibl5jc5QVUC+XASPZtIwoQEiysXM5PZZIo6TOp6NbI3W0P6H2L864mxhzNl1cFAPbARg
/AcK/zlCrDdClmR7qxmHAQdpMzz4vbNWHzIfSCmL8q6mTRLYXBQbgy1wGOi3rOeLjPJEOFjZlxLP
nTmW1GKWdn7W6L6xARwCKRUteLfWrKWxG+zoaH3BhA39xeqlOSgp744DwVcXbDDY6Eyom8C4GhDc
oSQpZG5MOjaPo0e7Awoo7fJSkSbPXZRx80Q3GEFEuRvVaIzY6MjkTj7DutptO/8fzvY72zn85UyN
LL2JhsgF7K132AaT2YwuUCUDnoEaOUoMVsRwgfE5KIYdAgIgmmghbznIybO3HN8oVntJMN5Z0foh
4/6mhVf8GVbvRfdZyPrmj+DEX75l1YB106KXMPb3X9/plpateV5LM4n3Ft5whyMBVkiMfsYbiqRB
1Mbg9PB2EheH0K/ZQ8uA30ttzEPaFLsdn+Bak7EZOUybcCDjTsgohFbA2/LMmhSgNJ8Nam5aioDF
8TSyjUj2yqzsjXXHyTKfN7H05Ee0zi3pHCf50kMW6LrkTDczQOOZceRlcdJ0xqecriFgxuWaOTy6
/LjJv8JqkNOHZe2bS2qlYf0IBlrLM//1z5atqXhYHGG8paNjLg4m3t3iVkTtnPr3SgKTV/SHUKoX
Nag5cLMT3e9dn82qUyt5qTTJW2Bwm9p38ztRSGNO5VtRP+XtKSDzopsPKXuXXnzkLUWJ4EkPIXWn
azUgVgrGwO5MGMf4R5ySnYh1HC+sT/ZIoAXUca8cExHuiMJx1ggr14XJBC6ZBx4mO0mKR5JFl8rB
PPhbxD8d8r/yyGJyKnEEGVCvb8dvG+UEYabuO5HZ6bDW85dTV2EsHcPvqrCQVedL6yY4liFkcihh
byaYSR+i22PCmIwQsjuoNQizgCYSPtRHedLZRpIq1T4A4uasSmXtpiSLP8tSYbmB6Ck9doZWhL96
s9aRsHDTsJj4dHIzvL9gYjOvTq3q+OykQLPfWaDWvTwNxesGwEUUdp06YEVL0BRE5ZFz8+W9fIZd
hOIMtsL5N3BRwaSTgv4J3U4kfBbIGfpTpI5nJ3tIhgFNwXHI53f8zQuCbhKG5/uFkcRVqYb9fvmM
x2plAOups/BaTveuRbYeb1SlFtSuMb0Vflv028VKUey/gmiC8zIIRNZs1/br49Pv3iEODG89Dipt
GSnvFB+hcwPPzrkHfVXHAzSlDBT2/lgpbBgstul/IDrjrD0loo0LslDhJ2fvNXrjql/sPGWpZpho
DfQ/s+HsAUT5rEuh7r0gkyZqw1h7zGVX6NYignTPeSkTJKZawOiKaG0zUpHejEvM/pxuLsU3mq+K
M6LSvT/K86iCOiJ519kGWkDoRIU7khncAu6IB71kDamaqMsLW95ZroxXUJINUq0NJka4eJCWqLEK
+R0NDVT4wwFgasDzq6jBGtmydYp/o8p+MvMLxBq9lNU5X8CvcQO2Xl8UPTgjpC+kCrw643oMWoyV
2TiCPmxy7EsbKfy+KC13luO3pALwye+5DVaCXMpo6lFds280jQ1O+Ckq1Wj3s/ia1pg1L377TDOG
QorhXrIgUudyM/+p+ONZqkR2GnjvFGRqpOjvwiX/+/XcMvDzVti2AnCCVWu1eG3FNAd5Rc0BeZ8g
NMTGO91iKROulzBgpbxz0mwK1uVlRLG8dQa3onkGMC6PV6RIGyHH60CLNAM1rdYrZGJp3R1lfZu+
p6zkWHmf+WvKp6KsA9YFSrssZEtHBlvqZyATcUwaJJxrtLJZaHzJ5oqW49LqJhIVM7uOSVjjOgbD
VmGGReY36schy2fQGrZ5YfT6zN+xf4nkrOR64MCr/3QvRr0WJseMTke4Ju4V8uus+c3UqD6cUUaK
sqrwwbUfto3tLo3pvI9yG7mjGICoGs4p+OHWrqphzD51EXF4jTn0zYqAPMP/oD/kyoOn8GZkXsqx
5MLmvBAJfB8YXxBkebHg7myzlgZVqDwT+HlV/i3Rwj6VNNPNXOOm2wXXZLJkwQPGXr0bkOT+O5aV
8+UAYccRb+Ce63MHN9acez7buNTQWuY0Yrh7YkqprlrH4rrRgAM/MiWj2GaPCRxZs6bpoe2XQurp
75Gh9B33p8WCtgMiJFymTJfIQdux70F7BufGuf9oLOmI8CdomwIHOhLfZElmc1tfR28NSQ+G3iNh
WfcvzPN9BsX1RNu5/+SbXdk+oCgSVx37Vh371W1wl9ZdT6yE1mTpCebtnHVcOA+drAbvf4zOFF1A
UZVurch8gFXmvfj1Fqnd6FCwqJKZexNL5UdO+vWlQAt5Ot9Mg9vbbNhIAnX9ozkddTOR3nyOPQLU
cZfNtNNhLKBREDU5OD4wD0BsQLbqhpKQQOeofzyU38UdDYHwjEGngael4X7UVKoRQ6gkWtFPJ3h9
4kD23kA1FrBf/OCq1o966C9mU7lXhyymgdSCTp1Q2y0CPKHyPERzpLrKM3lkFmtkqsVsM95IVX4B
+JYSzkjqC0kqSIkQqOszLB4YMS6fRNvLIMt/yVnAHws3DKxE/hjM2qXvoLk5Dy3x2fb1c5iNy61f
0qkvf/epnH/E6NrJUmSUrGopOdM6ABm6IxMWTvA+TrSSdtYyhTV9VHlchZfN1tFYwgHTJHgCg5Wv
ihMezlIR4SAS3bR//4819M3Jx3x0YGXTcd7l0nv6/Xsbrh6Qatehh3koDZuvML1ybmf5vvid1FMv
pYWJsbb4wFdCzWmJwH3xAks5rbAb1nATKD4agGlBgPW+dfEJcoWiFQstsK1qwMuAaupFnknQCP2q
La6YucqV2qNiX5Im7mihm9WunwQvMo3OQnAu23G2YY8iVX1IsXmYoDjat8MncrZLUHFJfNeXpFNi
PS+CvCLKNlFk0wy7pIzV/Eym7J99I9V7wDwFL5IuJ5WfGmJ3E27TH4HnJeMTVtoBQiz02xezM9aU
28TejASEkUI/cqc4oBPelWzom8XewYBpP1m5XHgKKC9I74xi50/Y4K7xYVO8e275bXrJyA9N1ieV
sH2yMaWCu3Y1WH3POXfkyKnSLuLddDRwXEv6vsdwP4zG5nCgzy3UxDTjPTedhpKThIj/boI8ODsw
dQCIGyuCrdXSO3MtJGN+MRhgRXRRGh6nigBvEApi884Zp0Lfo+V+VOqDRTc5cqqg/cdsdh0HgHCf
RSDLIWzGWfXF+Y/nMrPa8EduW3PxvJ/7ZVo4joJow74/rb4IUerIFrJcz9unUdxyFkMqjLD9Q2hP
FltPjvpoxTcGVVpWKncsXmX+m3kBA2+mLzercS/byvtyaqyaklLvmjzzOr/2cymf2F8VSokbI1yn
GXpCEYwoVCjJnAH45DWC/RV5MCPRjPO7MxE4Cu1SHhtK+sPTujM5djMkhLRlEONL8UArx92nGS+W
xCIUciLGX9OOrCkRzGdLnsSAjyW5CGK1tWx1vSHQa9kCzQO4YXyDv5sX2ZwITgqA+McwvOdhkzWY
l0XJKxR32vkqwCc5txb33rVNhb0IHBFloOot0ibinB+lIcwPU38OwvE9LUENBG26MMmYU5m+mCCT
NoUjX8IpYtmZZlmyowaAzxddKI73rJKYvoO4+bBdnIB0btfxIPp0mnJNAdenlnhtrWcMJzj4hSID
NX/IQcSgYoMDW/wLQ7nWMmPJIzVo7qErX9hHmhMg/wVHAyQVU2YqZiaRmqMe1LrpXK6p79GhbC8j
Yv8m4No1zkNXy3FtNyY2Tfoon93I2l+0Bobgz3sCYZMkroGaACQ93Q9dlvXUY2HsbSZZIvo7d87q
z+JSPvDG/ZwgbKAcIqYt6UqYJYjmNI2cZZ/wSZZiYGcQEIU0RTu58UHQXXM9bewnmANtt/R3Ixxh
Kv8Pb16KPiCB8D4eTfvRoxBu4/yh4IopHQKqxrm7OCUn7xsPRatE8cyiEgdVyOYHNIFRuVQpXoRW
AWJfmP5liYQByWlwPmiNDr5KZtouZ1pJa/eGTQ1Il9lJQMeQEz65xbfe7aX0U4xTCy1rQHuzdMyk
fwFI7SkCInp/VyKc2minuajUezLYwq2Vf4uvKUw0ZCmeaiJvXlQoijDmmFX6onF4yQVBFx0ITqTW
cekGkj+beYIHKoH6tFNO+Ow7ig451n9RalgqsGrwRdYW6qo9mpk+HGU+GDPp6EcXgXzM8YDcOKoc
TbC9GF+cAQAGU4nHiD8hKikhDxlwCWjab1IZfvhSXda+5XTBC8BqfrpANZPpoF+2RssGf1YkGc/v
vYyMUt+y38NEefb+30mxFI5JZn+BdH75y4t8fe1MzJzz0sJ3aLnkJ5InN1QBw0xPPXBc8VV76U9j
oYj9Jh2WsBAt/gAgeUMHgKd4jxXGXukg9jB+KCPzeZ5kv1FhmD/1WxwMxGiy2kHehPDfW2BvKvXd
tK+LXMrWH7yLXxlhJWGBX16o6TID9LbUC9Fmy2H78dnWpozy7YXnNFKoSxjia1qajcaaKMC6kBrv
C1bRJtP7GZ7TrTi/kDlHJGl+SthOpBu2NhOPakA0kgEDsV7TPIEm152Xz5lCU6QnHhyAB5n2uadS
aUzNGtDpEgFgEsxO2WA/JLssb5uP1gPV5tPTkhJVpBWR0TAOibard+V/ppWSvcVNK/EDK1JFQt6d
O03VbHU1j/4VlpJJc6XD7HF999AV08YdSqeNf/OE6/XBJw7OuSW+sjBnCNewzbsRtH9FtffZ0bVv
wSKDomBh3k8tJB1OpsA2ESSmdb8iAUSJiwpj6EIPlOODdE2DGGYh8frlpsBMXOdW7LNP1Se5lohi
ASEGVYOs6V/EPM9TohMJfla0B7xfP/eJh6pGBfHgByC0KejnbPYuDHkLnPCL2pj2CwPLDjtthatQ
fWJH8cy7TYiYUYbY+cjwKssLgKPHeVtGJPktIchSh7TT3mjZSD+mm6q6+GfUeTDvgCRCemLSL3TC
+YaGR0hcwxDlxiDVnadRTJLRxfuVzytE8SWCSO5zzDVsxiq4U84yEuIDmN5RpKH5Lnr7ShgB/8xY
CWJwZTCV23NfbAC+sHSb999nm/OGT4Lh7VNST6ChjYWlD3JehrO00FIUqTx85bQ9e82Jm/IoqFpv
MxF5KvHAyepBTC4YrxwNGJyeJlT78z03fHfZgCXbyOWGj4LFNNuOTDIyH+DY2l0l6M845xGSY9AC
uE1HdVihx43jBzoQBu+vFflS5tDXF5gmStDH93GRlnVRFt0y0IJFGA+MQ7p2kqZ5uAfxfVLP+7xV
6gKWyr1Y5XpsdqpX3NeAht/ocBko3FHTDu7rYzQNPLFfrXV6gwimEhmVZnw4ZT6m+e7bBvwXiUGg
N5vmm6AP15i27C2jF13buhpqi34dFGKZjgjfRpqNAjQkYv2LPliwtsOqcaXzR5QFJDyPwcJNfmN2
x/KkZmKcS8ENRpEzJACIgI+bTQUBDcLDeEQlTWQVKxsMWqQ5ys6d3fHeO0Qkpz40OzTQe0ImVpmy
aKsOzdT7ri4lR6eun6GBU9cd1PQov2ZqcItb7sV7FBcl1kfjkAmYDjg7lBxkCEAdRkZZ3NqMI8Q3
ftEIRwiWjh7V24sCUmGiBStKgodw1QYdF2j5cEdwWQ40/SfNZYfmO0lW9ufZJ/obNc+LR8pDJMSg
pb+58rL9s1AG9F27j942i1e74ChVi7M0bGyZJ6VdSxQiu1dP7qEVngZp5BexO0JD5TQmrwY3mBau
Md8x5+l12iKww9RxYH3+mURY0iF9kKmI/Iaz00GwE2NYmmEHxykbhG+4zPut55+kllVKKh2UdUl7
mNK90nvLNwiUZAan1BIzhFzZVcqVSqXfT9IokzNW/5H7pJUnpR9UeUlKk2SOR+v2R0dMYmCNwYxe
1SlOjKGXYw/Wn5Wt+aKfiZHPvxLmzwxzG8aAsGPtJwEylV1lNF+vjFg/3N1PEKdwyYQue7eRB4Zh
JV3Xkcl1o9ZDvtKIG0IgEt/5/7KbDBygM8HthW1SVwKgJ017ivkv5YBRi/M2E88is/+pGSVTaTKR
z0vCWqQnCD46hD3MzQ1g5LqFgw3Ont0KpLi8mg4KnpsfiyvpNc7e61UbmwrBM5aVgUUgFUriUUcU
RTG8/evsSdV8rZfb6jEKZmG7o59MWELMjxIGsJNxYkPbRtgbyXuHyeCMoSOsZKHLiV9H2jmepdRc
ZT/n0Y0jQTY5kFIgVKZWJPlmOLwx+bYayx3KUluuvfPXFIeUazOSwv2Rj1GyTdJOFfIGPXmklz0t
6qKg58PN5DdMB5zfrXPH6uc7KbyHyQDTVuFql/WroKXKjAOE3+F79DDIcdjD/kr5nmBTCnd/PWJs
7In48iRCzKlqP+WNSclCmJacAxJDsCEu54FRzOHlPReRUaforzlJJ7grg4fbjvDnAPzpA0CzXtpp
TuLnFIkUZto589DegFUIO47f0D0C8eR96IxeF8WIDf6X6sC5Axlzw92rayQIxnYY6beV5+al2uTw
vB4Sdhuv1hvZyodLlu/UWfkTG23VaTZQ3EpsDQBMrYgC4V3SrBx5fhqe381IY4JI6EkZ1Cw3xl5H
6BUmpEaQEjONNVS4DhuPL32+UB9j6lEEkoGi7AX7I7azxqX+horjIge+ptpNIjfJyJqAhwN6+HYu
I7/f+WOR1uc9wwkg3DCBWx5/trZbNTwasfxAd7bLlJ6lEweR3pXAIvuU1Hg0z98rtKt4xPbhYxjO
uwZhYaGiPSrUTV5TDfKPxn9MHuGaKEUdbOU5z/6Oa/ragHxzL6gf9uVzh714EpU2Y2Z9nBXSiQWA
OLfVpA5+bKDWAgNu/hhtjcRQnPBYNgRiEPXQ6483Ni4u2rX1LUmR0403hTWcS96uPao9JacPfiU7
FLcKD3bNaWro3yl4Cn0CyHd9CFIEP16xWNlUMOJs7qP9eQJpgnxSbMk6kjHOkCXne75UXHUX6Msw
8j0xcG0xplArmlMPmcRmW/aQPqoh2vThHliyz63HGIOaB6/8KCDHAX+8hBn1HbA4EpdG0mKOROIE
GjJD3s3HxrkeITA7UQehCl8zVv8N8fB8op2io/hwu55MQ9ixadCnXvsO/H2HWc4beFJdPQnTzbh9
MRxL6qR+uRU1t3sD+Gao0jGtA9OIFZKnMLgQp1QnWEFXfBlzdSWheBF3muSMXlJ5GokTynjFjH2D
uNndl+sFbPUwm1tmd5B/c83f3AGRzOJSmcC3V1gpOvroTXCfsQI8jNohXr5WtXX96/WOXjgXbCxv
jrk7OuBFUhR6Zv2v6UYb8l3Ear5Zx9qK/4nYjTsoPKDJ//upbNK7Asqs0xkWX5gGHHTp7JycRLiW
yG+9LvoQo9Xu/H3eWJ9m9MKXFHToQC1+NiwEPvWETjQwxhgLTa8XqDD8+R5AtFcIsIG1EolVF14b
xpML8zpbJuYAW09E2LgFs8qINuA0mhShF+UwqT9pRNIZeIZ42R9uBS9GS7vdGEnXVi3LPFDY1ACV
oly39onopMaQdhOad2yvaVY8HAcDNKtlyhUM5xqZqCGplvZNZ7eHoXZ2BkhL60FB4mi1MLcKFHsO
T/Rg78EBgAujxlNyrpHJpMdF7KPyY/YCT2ckyB7Auv7pDf+d7FIovlnface1aR9F9qDXyXfV2DDt
3f5VHTloK8eTpH0mn6X0bnxAplxJ5RrxN9Xps1TEyLBbR1gM/1TW7zyQG1CSd33VQOJKSAxoo4bE
2sXONoaOLy40xzXxFhq4ZSV85hBkBjcM/LxG95DnhvnH2Xzl69tpysGRblQ1TjAkqyYlpvXvdKNI
BkPb7JF7M21xWimNj7t1K8SKzXuRHDKkGj+gs3mnY7KkE5NfOX29g7dnhk4rfZUf+NQ+Jdszfi+2
8T6Cy9qYsZ6STgU7cwFHLSk+V8iKZ70ZEv+KJljqOZUfg5lZyLR/I1z9MESYhsDkSd8VKwQvEahX
jsG2F4bFqmbjfx2lY/iYiLmwlYgKVCXLtx7+w4B/y04Tp8Y1XVL6afUGPlIXif4Hg19/k0Nqwwqg
fAK2Tt8f7meggS4VZwVAn6Yyso8vBbAckCmOWTGjOuCOFHBElxkwORGU+y/kyu63nxqvw46oRWzm
T4O9L1vWpVhNls6H0Y3QzCtL86ADlMPnmPBJL8dS0YUwpgUOYaicv3KzyYLnttGkGEAYcyQ3ojLw
o8+XJAKkW7s1FF3KEswyeAX8hRY7l0lU6fUvUBwlxxN4VzprX1TRi0FKdL7E/fApQ1FEyA4ANkOd
92NA6Ape8KGS+7HQdJOcW+id3cbHdEXMQS1BMQ8XaQV0wdGyE2SwtKcV08wm6wa/ivaQssg4cT6/
zxUVytGZhQtFBE7O2Ihtc3Vw4QUQcw4cqx0JjK+b7XMyg99yP2X29jQzx1ZBxGMaG9wetMnIZn4c
lduApYYzhC9lXOV/6Mx9va4Njr5dEvJ3g0AJND/a+imO8Vc/dZqUnYYp1fzprDKnNmFeJ0PtKlHV
f32irO6QM4euK2NjGOJTWChIh1qt7uIiuzV5t5U0ToyK2OxnwZ9G277jzqU5rVqIl1vnES4Ez+V5
NDn6xEWgcE2+9+YL3YnqKjxAZoQVP3FFqnhjfXehaiyxOXPMefiT8rni/c/oDHW2MWJaeGW3k0nV
ZwcUxmG/92FHP7w/cJ3Q862sJylZuCn0JSdkBTq/y5rJkjZObfa3GiLlvgEmdUfU+ybIHXwccJQn
ER0pjbtzMUTQd2sjCUfF8tR+6j5W16BIgnky4/JklzgrRxhg8NcN9z6cPIoz7abmnji2ZaC0HHCl
MGHLMje06kGkXHkPbUweveyDjTB8IQ6+l+cy68xV1Yr/IqFMkDLinu0aPXgvpbb5se2w/sRMV+ku
52NiAFAc0YXcYDyuB431vXNxpgV6/+zeW+l+PUYvxcNkzhadMVIGLeMUAieMsvsiUnz0vG6D5QcU
ylpMp/9ES4VtoLPK9RK+mS6Wbdhrps40xSr6IGG9BJz3VO8QMPXfl8rgmkUuIu1oFWHMovAGRHPO
V4BhjFKNE3Wkbi3I0OxOaPVJf5ZK0mfVQGBWGlDFnwFJ3311WiVOzQC/WK0efIHtFOtgwH1J+/CM
LI+JEedDYKnKa0qnXOPSk0EBsi5NHHvfd3EJr1XcyUsRGaUUOMONEVGjqzOw+4lAKw7XVpQtLBuj
frjrqN+GtJXDGS2v/6fI3QoZELEVfMdRtFOJ3o7vwPi5hm/fP6JnAW2Zbz8THzR1dgAD9/q9+5Ss
QRLf4huO8/vYu3NLXJyGsWVnU0wRE0imoyFF2Tp9OGTYDdVi5A/yfqGdMtwrarh5rEwOI6uqHP0e
RDUF9XBzX899Zgx/68PGzE6PtEJdSKK5lEj83Zc8/pj6KVQm77RxczzjY/fiLXQwWFzIMwe9g+Vf
0mE+I02jl+dPggoCFbxg3O/vPnan+idKyqjoVloJNlBdPlLygujuIEtvffc8EOJSQ1JIWKZOzFAz
sjtjjQ51iFiEG+fnhA7sMfi3ZU8WMrgIB4LP9nBt/nit6FKtHnynNkZ0ZtwuUK5UARjdC6Pw88+C
aXyV9KUpOTWL96c9D5molUb3/fqE8tKQ8Pg0Wcbv06QqzgxLqTvv5q7QgMxkkW1FRD1LrIfvOXWJ
2SGJqBh0zMu1NnntDhWZxhBYQtPd556SF2RQcDlj/3E3ZexbLRcJ02hE6fRa/NW0J/Bj4Q3UCIKs
XCQUnb3Sqk8nhmtFLO668LyegHZfjmxJ7O6W/uvRDN1qsNZzvQKzmzcbDqnKdehTD3Q2nm67QUn4
p9QOLAsDIGfeqWrygS8KesYgANoNf/gwYKJ8Nzo9RSsua2EMwBkv04DnIT/i3S2wpLq+kx21u50x
mrPQp1X/KkL+O6MgYMzQGisRbIkghPs2f1rE64xFj5gV3GHpEpc7fswdAUgQOxLC1gvtnSVKW+gf
Y3ihbjlIFCU/WKTX/QuO/Gz56sjV3AmknNX6T+F26hRSzJk+e3XkVDqH+9EhyMcXEmqqe+iYatEV
hHjiyD6Apckci+PLhw6sO5ddctFLstaVUVWMnkAC585M6Spt/14voxu31AXhDfhSBGrNTSPh2kJ6
sgQg74ybl1O09uaSi30VxDtdgd8eWaSaKKZuxRZsSFQjTHr0qpFnsPBacLnReuLALqOxd72SRpdE
0vm5fiNdYimKUDt3Otcfqex4omZ0KGoR4ybaTTiYG1mLKgL2rhkQ/SoFItw0LzDCc0eDQ8w5Xo4w
Lb+6+7kWqsRBwcUMWhpE7CqULNfFnLHw/q6QZyfj4JzSHIZXHYzNYnJQk9/7E4VXp62Kng6IEEZg
KpgWOD0zom4JSCCn1lxkfo5lcINXdP1FvcBJ96kYDMn0DocMuCUUPWn1NxfwJdTxS/PigAcHc1np
frAf+P+XEZAY/6wfEMAeldmfTSLUugRbSCZPuOcxplk4ByMXjCfillSDLGr+52xak/kxQ+wnR5CL
Yt5YMnkY1URWm86lFVf0DbROzcjNor94Av+DDX3YwU88CJbxc2UCFCaMuTn+KUgU6DrT5el38BIv
Ot+hbqDDq1an98Chidn2BlStBIMM8eQU7LLJAldPHEZfgmp3x1Bg3clbvYeBkQc1yzQ1Ayk0t3R1
8kOLIVSrOEc769d2tx1cFOIzFsDOszDNPDNxVwgWYdP1SgcJjqFLsMxkws0+SOR5MMLFL1AUAAH1
uEIZ/qgG/eszlgaIeT+Qus4IgOs9ISdfw91ormX583VeuqR60pkJnVnb41Q5J614ExafdjOgJXFD
KAgRyFlnrjNA6Wqq27L1SaxgNY9RlAL2ZcnLqL91HncaVTzGQrAKBQ/xivjaTDqt6YIFxLmUhQsq
Kz9/OL+AXuTn1+bv/MIdcTry9lm+80F022MFbSoZSJsFSzC2x3bN9nX2U/y66AV2/RbuCYXvn2S0
WUFs2W3wj3KcZiioU+z2WIiZcJLJ4HiS+f+Z7cYmJSJ0sy1jHpSeDXlKojL9PWlJ/JiJ2NY3vT9D
gUtlQXacguGNyHydt/SPdRWxZdFimELq2JdAc5HnZc+6/W4pTA6FRuK8Csh+OqbGwTfefUFhvkx9
qpKL3wI1cQA99TlhmuzhBze1G2+DVylbDHOwzjXokO86buwsoNqPz2/QpNppsX2BHuCq3cdW/Nvr
uB+cQqL4fsjX5G5+0T9naIa81IMkTjwWqwzgpLeBca6OW3LZHCLjpXtzNIigQertMgVMGXG72b13
bamCwIUGHgNaQWetLutSpxEqtAk/77s7LvX4OvL9jYXVAzmPwB0IAsy7W5hUEsIF924JusV8aDYn
RYA8+IzhlfidMNWI1fzSn2rABnjcqVCIUDXlEgK02qAhBSHid7d0NyyDdlp1Do2hMXUI9XpnVwwm
yDCErbTfiWgtHImdB8Es88gBWn/0RJPQvoMHVM0IZP/u5j70Hj565P3uMvE642mrMU01RPygqu7X
MpEo6Wj5l5Stb966e6GJPJRzYFEuIicNPTxtUsv+RdMuU4qc23rtsgbIBd/gRNJAf3MNw58I+xep
UrsERqWVar4eqZ1XqbS8xobcO9Mj01q4t2e9oOl78yH4UjCJubkIHcjgj8LmMY8G8g8ySeNZX9MC
ttDeT+FyuT/IgGyy85aTz/FqXbTmX3DeyAvO1DVzswhJWWFUXYEoCpT6YicsRznGcSdhJcGhweM4
RoWZD8PFx4OK82BXTudsH5gNJ/+BiO4bpBKDUoT8PE6vYdWs81XmA9a2/HumRnNpaDbG8njKPsiw
SoXwq8W62VhmUbqZaAqyPhLlvH6dC92VkfBpTmYPWIJ4JU3bqm7V61KmYqvuEyOPQKrs29uVauXO
tQ6hiyxv8R0qz1cV6WMT9WEIDqUGwuwbQLEDu6bwW0MTsmNEc6btWHLGqVzjRrYVTcJX+y68lttB
pUUnco8EDKHAHD3AJI0i8nHqoQAl/mJPt6Eqty+8nIXZ/s5k3p6Yd1aKNXErqwP+Pt0k+Nupq0q/
Ln17GSs4Hg/o+ih7wvr9S3PXGRELmWFGSzQ22pY1esK0NMg8zTKgnMcaZ/9gEQkXTm191EBjQD0a
rNRfLxtpDPmgtYdTzMMbWVNgTA8D4a1JVo2n5Wgejx9hOnW5Yi19ujXk7VvJCOT/wuBCe6Qdnfzu
GYDvS0BITmer8/Lb4Z5R6X2oQX5EgVyz4jXCRlRVK7/9q9Tj/ROU4d7ZPzEEZ4ZBJKM66c/+OWAq
0iNNZgR0wZ1en4pW1gS/sj5Oe8G+COa1KNJdsDT4GBoUB3rOXrMuCWOCdrdV/r0g9rvQwFbSEiqI
jzD7BEtdE7D5FaQGAKH2NicPEKHw4XJHlLuUbCI0roLQuwu3g8llhR7gOQpubD1hf/v/FiAoVFYl
YhgCoAtOW51mS1iXIN8BcGpzUMK6Q/gzPS8q6vgRMqEfRijtIkjcqu/OCU5JsYeI62SeyNqlpR8m
fYa5C3ewwZxZa5tOIcGtsMdXTSe/KiCp62W+3tHI+jU3mPvBxsQDpKYg1cxZjwi2j5aafve1bTIg
vgdXuDajOd1HSYf88MfSYFoljaSyQBJGb/ZdkJxnC4eulqyLLgNUTYjMPDtwZYedWNKIHDmncJqs
1+Dy+j4neYIsXM7jQnRtr815If19sqPvENkYmMhSOduFHA3H+exWa9oOMQP4fjAjtt4dwgugSGt6
6YYMrCBPiT0aav11bXDiqp2MurmPy302A9Sg0OWI8q4eDCpCMFjAags/OqPtrLPDBQn0ysDHcwWV
2vBgwmyfKKTeA+84ozMpsMBVeVCUfQ9qo8Ze+HSzVKXRiW3JayXCclzuu07nlh8cLgz73gADIhY/
bG3GBiaGJNLMv4xV6b8hH1vqF9m9UyWLqagfXTXg0ZTZbvcUVYZfGzdLZsgQgBd0h+OoGY7J0n3G
1E6s5wkW5KI859CkJfJNONqTm6PLVHrIi2VAT24O3psO8H+bVdE6er8xK96hrDOqC3rhCpRVZbxp
OGVF/MV/5VnOb8itcp8LV58NaFqeefXtsZT2tiTGom2i/HqveBPfcCJ8Gil9QfwtQkPKTUBynnc7
Z0I5y6cLRHA0r960L7pk4zy0lmFeEUaEvYPpPxCunnB2DNQdLixZe6LP+uvVkLCV3SSatUAi9fD3
1JlDa5LkUie1S6CdAGvi+HLsI0+E5CL1ggcxReO5jiKRCE+J0jw22FOn25dIJNd/pkhdb8AwObGd
iaBJkBKxNiZlREAvGYT9SNr7UG4XXHKlei7DRnk3ST9wrDui518R5yEtLlIeCS5HlkJ5A2PW/y7E
WmxDMUoiXLkSRalZlw3GjdEMd1PwsszSUg0LDl4WyXM8d8wYvh3MQxnFfU9Kk10QZLK9Auf/WGr7
sNLwa5KqP6FyJEAX8GB7fM6eE+6YP05EFK1muefwzr+txxV3V/dT4vbsKI4/ULJiUfrUBfYDXec7
7bhKuO9YwEJjt1azfRvUy9tvceSA15g28uS+2C6Sgn6lnWxM2sADck3WRwEMq7DMnBy57HxIsN2U
eu/VmeZnki6xcOoMQfzF+ZoI7PJ0if4NniHc4Z0nadtMHArh0NK8mBI7hMW/mK2Jg0oXZokqwM/N
5f8fcrZV/QUTVT7CHmTv1Tk0l/xulMsdUi473sh/jVyIo3y80yJWas5DAWJ7ngJ54lsEZVLbtZiX
nhoZSgsG2wucE92gNnUkgpKqoZUcaI2wQ12mhLemc5+EfDjOopWEbdyciqsO/TZajLiG0wbfRIzC
zBdPEBd0G2hPDDhFwVUgPb3E1EbmYI471sZ3JNxsC3q+uaSxeg5Yo6LpC2geLVaiopI8vvBFqk81
EcAeLvnAWJwX1wQuNGDmhRa1ygulCKwrsH2kCusaW5KNSaI/QE91PjBYd4tlNNCultUGvliheTMv
j9QrG3jIqXJOL5NHWnK48n2BwcZwo1tur/NRYoDd9mj4ktJu2WRntLbF3/rBLGqjGUQUr1Uf9+Ly
EZaRkeL80Ck+YKYEAeXSAeHmWeYZ2D25++nfnICvyis9vUAUFxK54ew68AgQ3g2GS9i9doIEW1re
7eubJQexYTW8co9VLIQ8hneHOZnjJk3O+JBKnk1019aN298GhgVXWs0kH7CjXhfnQ639QrVrNG9x
jmZ6mdwpqEilK3+2kWWtnHfDtbSPcYQyl+YK4dy1qCwAG1BwUcMmMPYOUHCZoI7cI3aeokD1bEWp
l7vs9bhJjYgkA4YVbe124QXG1VeEkxY+xhWpalncl9YPJySleH2QL25ZhUACLWA9K7wK3KrbF4r8
h6kydwKIu0VtZ43E+jeCERlccTwuGQ1/6eU7rFRG2VIVTX/C6M9qP2aIgZ7rNK2+a+im9G+TKf78
fWdYQwnFfFnHSO0HII09zp33S1mQU094fZAT9phif8/grFFh/NXm9WvEYM0AeyhUJ1Y1hEBrrLjB
U4jNSyv2c1JhZwIRMDEZrFXXfOb93UzJsne3XH3eIejjJPOoC5RYQ1i32zRzluythvhsov9zSYGs
pUJT++mm6p9oJrPUUl3d2C7vZTlcUpu2YXC7HTA0t0bhvbZHuklm9T/sWCO5xXe0iKbdNkJFPg/8
046VaGI90NE34YdEgRneZB7E/e7WYxYIcInaY+/sBs5Y5/45jrWqJFyX2vTt5EU7LARpbrsKMicy
1CMsqJysvOl6gjaBjjVi3fBIRDHmEgPATWwssQvw7dCh0ywoeiC1dmU7FkmSf6Hd04dlnvgj5D/0
onXcK0UCpzRjX/aW66+4NyNIriWoJEn2Kc1wWzYFTarhUjlaiBEXPUjHYuVwW3a3dj/0YZHoA6aP
j1/2By756tmzij12vQiPw5qrWBYpDC3MUxb+D6uAS6taOxNc0mZBWCjsrjLfssyIAC/q5tPuvkHz
du2ZV87j0a5JkwpEDsAiHf7GkygunGq1g6OdPfD7Casfam6ecGMZSfCgzXIOUfqi3CTE49BlZA3I
GPZZIx1UlOtVd8vvpgk1V9VVsQTdyQWzXA0Kx9Jm54cX1vKhkTalqrYVBu41Bv7ehYQti/bRoY29
mzCautqRcrtsRiY3YJpJ62bwwnFduSCn/IO+ChyLELGlpkFfCnF0DWkqlse3/ZEeI8NOmF6xIY/7
TnJIPSCbmsO7t8dG8tOMD79xVs/6rH//SUajyQVssrscJ5/fKKscxXpbDg4DQRjc83MtkfVUB2s4
FdFrPPpFPletkcM1lWYJOntijBJaYvS62dQUxAC33Rsy3bCB/lEl4d8XOylcU0HD46Kc/uk7zoCd
FhVrbGP7uhJ7NEKJDniZ9wYnhjNO7OU69V0udu8/B/CS8fldVn30Qsk+r1+CjOfOwvcrN4g2CQ1r
9RlqtpWS+zL8qdrQOYZhvwWPVP0jf4ms33O/tk4xLrH+x3XdCU0TzvmuprG2CUI66j0g9saa70OW
p7I6UHKPZOu+7Tr7v8CffeaQGCmQ0mEaBJclV5I7WbUHHXQXUdOZWWshBhEaZfLS13b5/w7d6Xyb
c7UFPRklg0VpSbXrdNLl3+Q9jf3caqdsrr/0OShKF81Jv8DnhdVuyJpEkKy8hVHo7l36GHYmGT8e
iZuN9jCes1c11NXgFpGNuSGDqEBe66TQuwJwCIB9JHv9jfGp2pBgBgA7ikQj3VVxe825admMBcwO
5gdB8jhS/4DSQgHbutzxYYzr7hVGq6vxN11BoguCxCPxOtjGm5lrBwj3/pyKNFNNDj8dsDC0thaL
QuuMoq+Z9gErt13nlEmJQA3NQFFeFSt8WdXXBovbaJnDIMEFez7fffACJagZqHExoBQVuKYnsBhH
qmaLXbRQ7zSjAGtkJfa0Wq3T1DHjtnUr6NwVKdilB4DvvG9rjl8TD5qFxNxVz/54cj8USLq0ivon
X8iJST4UdAo8+P6I4yo3B6aaIJoQEsH1v2dan4nLG5PN/6uL+tckU13AyCnGQya6Y7We4i6MvjjV
hfyEWf8GEwp0aUXFICm/9rlGY84Z79b5GKOWQvfKIwRqLRdDVm9aw5RZB/oPG0pNEiUjwnxa0QyP
TbK28BMiavt+FfZ+2YqMi9GLTgGQvpvZbknp+zCsHbJ6EbQvl1u6iHz5RYS78JphwJ/h+dOl82ez
MkO1DY7Q7EV5atfzaZiQdVhDKtcav9oMKpk2kXD21FeabXN1WB6fYYa6buKyDb1NG+SrBG2Rd2GV
n/YRLQWEMqU6wGtAjQFU+Hb95ubl3JJu181xzQL+yGICh1VRlhgeiFsxAI7amprZ3wGMHe5LOYWO
DH2LcamQx6FQEyqxSpXL3O3tZkpfHC9LJKCqyr5M17KmyTYu2wu6QHE/1PgEEQLdA1iOtxbxI1NR
n/AoLweCP4Rsbjh8nilyzsQhGvEqYpwPnNgPW8IapCFKMQL+2l+2hTgTHhvM14anGCQyEGBQlQ4Q
eIeLwDCJUomqrAmpr/A3NZ3xud5RjIUt655UdqMMAb0KuQ4BxlJiHNkIkNf+WoSwmMAMLFeIGfN/
FU4H5OPdfV0JrD5gLNFKttkMeBhLWiMZrAULnXl9LBY7Q5B97wBsUd+ng/cSAB2w/KMdTnfmhttB
sfMCb68bf8hdmKy4/ynw3LwlNkap1614mZ/5zjLZuTIKtqvZKU9PjOWfFw2Lv0iZ8sdxPPBWGnBx
G7VLPfm5J1lb162/yFJAL4IKdSJanlUoAumLtoaCPWV4feuNtdV3g+qcdxHDRhUEcf3EMTQ02ITy
a1/HfAmRumMsNhAuAMRFQCj3BaW8JlzJPCwcpXJNttwUpp2BqC/VYFf/lVJo8ZiWrQtNfBEjxgaO
OzE3CNRWrStEUwm8i3niVvXkRRTEVR828oHae7sw8jxhWyfT2oaUuuRPNhPJe9eCGX8Ru9qYzLzM
CJW2xy4XX9qUnESnDdy/YkND2VF5vQMAkHfsOkpxDVWHcjX3zMDOY+/Ed/dsYSvVl/AdVmHcFJ6I
e143PluIle+0iHDu2N5XV3/2A3abIDHmqLaEziiF3DUm1eNqpOqBbzPIoRNRxCkmoJploDmdAgIv
M78GyVhlpfLAsXW0RHpLJE2xqDERomqOXwnjNoPBtNperPpy+ki0xAO4jCjwRndl5jX86uIaU6Xm
tIjU5PDhT0atTVfc4hGiKhRoSia/Bf1JosPX5Uf7jBIynTOEgM0AOkauwJ83SFMhom2QiRzXZDRm
qwc0RIHdaMRD1W/32/KhSiiK9mx5+BRUDmcPuM2cDnd+Z9h2YIGQRtXSC8aZG1o5udJhXExdrfT/
N7NwWW9P5sKaHt/Ucn//lHAa32SpsiVGp3N+I21lgUefMT6KZHroaBMUBklgrUq7TxIv/PwSDa+X
bUDJjzkEmF9cvsb7q7RbLAr1RS/IdeYzifg2+PERPkRhVGrfXZvKRRDGzj0yumklnFrHctHtEoH3
cq6P1q2ZCpP8lL8Tsoa7vU7F8ZlVSl4vheDZKjgmz7mFNzNJInxnrth/e1h2VByJV++macHavRR5
/gqHgvhl5uqoO9t1x9XzaTuc8SKgYMlQdy9eXoLCfmJvZJCs19BSfpk29eljpFrLrxs/nYtiN+9Y
x8SWzc0qh7bcToimb4+WdY0eefHFqB7gVDfdHXLmt7okB2/urJwhBUbeFK2afW/DuuhtKGOu+wcV
ExFV+Vpneaw3rSLJf10bNvsv2FPdYwLagxYGyJwpSsp9ygFQLB6n4CbYryj+7x2fJlXFIbgEAIMr
bNlI9yo9OWr05iHQC2btxqmFVaNIuK8CRLAXunIUxBVvU4Jb0QiGS9Vv/l+2Or0oNJhvak7I3jS1
LjfH57L1aQoo0yOFXsREO1QgfFghYjQ3+SCi6WQVuSIjucMj0h8vlUoGBG9w2j2maO953ATPtEwY
p13ih6KeGoOso99tkQ3mh2tQZc0lyGTdnYYjRujmfmrV8Xm3qugV6vOxCODf8KXQsXnf/BptN8Fe
4DMgUHhVHStSx1f9XQvQafCGVsTXrEOvRVWcPAOILzpXLfVKqTpbqw3iG/vURCd+OkXTOK3eYoUB
MewvAJjOd+3tETt4uP99Bl80hoGwfnufQRPUZTK4qAMO/+uEyOf3zY1xrgoHqatPGtHnQHBMQ3Pj
dFMyH5o/T/PBEu2/rtBApq1gblTITBHAxnSno9nWQLPfaWzaKo1hJW0bejiH9n40iunoS6lmH2IF
dYsYOKZqj6gaom0w2m/wZ9RRG7obFrytE0JmlV7UPo4YAP1CtPRIW5BbXPAHNg88bIGbmyd0ggsx
6jMcbRgD+EU16AFrM0qNpWvdYbCCFwoksLMmqiJtZljaoHmYUdbb/GbbT3b2xnC6eoHbt+ft9FWe
8ry0DNyAH7WSQvw4EwzvTV84q21FxIa/HUmWct7UyWpp1KJMlYBgT7KD//m9EZ/0vhOL7JgAHQ5x
HZdfGqY+8+2D+j0C2ouuA25jbhNgIwlja2gPgb0tI0Ltbq4uGbaVne20qvzwXSrBDHQwN2BA4R4I
mgFU3/rMN8Jix29XRrYB4skW8W4OR1ErPUtQYLm1zAv08JR5KXtbG1a5bkFABNNtqZbzh4Gf5+Zl
+CfXLMtq5GOSYkWq1HUC85a43lOaPXJCP4qAqg47EI0PRiOBT8RR9lW5+2vFP1zAbxVfz3/hxToZ
3Kh3Ouit0IAOsIIT3eqcMQSlBOX91I9uLv7C0hA9/NTrkvb77LjuoxI4sWaufWVonjFJJ44Qmzqt
zQxWLXI1bBI6BZlCT8tAob471EJzRX7F3VFoXc/+QAfOHmqrHALAN7CH5/mrI9Ns0CPbZDRh/Uzb
YciZxfMbrKmCSisIymkwbZW1pJ31oAr/fkuXowlEedKzEsISa/S1Nz/KUzDpvwjyMYEt3p6W6wi0
FbAg8ark8zM70pajw6f+ca/Fo/mmpym25uesB+HL/IFk++sHwqVpC1/oOrjngAGQSDWzvoW9JHbl
g4Ajq7HJVmlMla3O5JqTCCXKDjO3NY20qPWKRXVH5iLOiREIcZwM/0wr1G8TIM24lVhVA3kBPIqj
25Xh3qEDHZsTpQHcZOluQyE8Hglw7xgxrU1VR3vxeKaEDhKnWxjckJhKU3argpXcGxhFVb7sdaUF
4rkN8OKnDE/O+rXJjYVlNz4YNGRnQlr4r98UxzrgCSDV5LeXiA+//PoNfAJPRTTQOBPN8BHhT0pR
vNgcffnUU9kP+rPAZc5qeZ9gfJP2cHcM2kYn7fcRdQdDK9DaWSbt6PiN901ppCJg56f3H8E7+Bqt
aKBbpblRjN4LGM6WBiLrtGeO3eez40FtgcK9QuYhkkN2XJskgR59AJ+uE/4DlkOWZ+ODxp/ul/te
b0H3YItPS21kTvlznmx3oTQ6t24R5AEjkGieNdnNRWesKYk/dSoo4nmPKlbEke3v7M/Dw5s1FDTs
8KuQBfwuEGvmRml0D6aR9+0QHA0Medc0ZNFn9HYrJfqUadl04eUM4N/juViLYvH3bqKCD1jWFYTZ
jxKJPJiuoylVBaID4Q5KNjmiR+d5L0kv6u59XMDsD6uxSk3rgkh/DXwaTsx9+izZZNJyBSzmedRp
RhMTbdTvVkeQ0iesvF7Ez9RwsJhfOEj5BtHcGjpOItHuzSypPdZDXDB9rqjT0UZpIGif34u9cgVg
9VQyicRlcnuTi6vZ58mvMv+BhDmOlpA8XhIt3Kl+20HZDPI2fLH80eS/tJHP/ATfc06SJcZdJrqL
fVTEEyj0sFJvZIfoxnL9ykwsZjWQ1QXMKi1oqyOdc+j6xtro3E6Jcht+GldambhpMzQCZJvueUfh
L5mL9CY2lUBpXcSnmidNXhB+lVZ/c2Kce9OtL/fizzDN8HHfoihnzYDRUYe6j6tQoYVQ8iTZRtAJ
Oayhvi+UgXORn2X/nZ3YVmZQ4rcB9ASlQ3NUUfYZ7TVujR9Ng98lmwxpbMS9TPQpxm4bqZxFRkYs
fy2auRZJxO3kROFxvdvyGUMmny0V8tq++O9c3p7ou3g631q3UzDmH1VC5xj3FxjczOVf3LK8v5qe
pyoSzMhfmQ22SC8lOUUqu4nMalUCpKhn9iLJLZCh+NXY7DcGOIhl98iJSNuNKOAOtDD42zuitZIC
wbc5rXDnBzOtblGNG2C00UvhWXnTPBVmHVCqR5yMOhnrrWLPLyTYpbtu8yRzLqgyKYqIYEmCLth2
+Uz7YbzwDPtLC9OZbyn1ngNB/e3wiy5lQ+qqvM1iNR2myVFmXIsByLXstgEtD7XkP/q2x/NeYvYU
sPxvBXu6dV93oWfse5f1vbY9AR2mNVDRTTzVNN7UxiP8FOVX+YMmlzTSoE7aiiK4rze3rHaOPIQF
RlOlR9zsiHNy51juBG3Gk26qQG2Uai6DsdU03JLBWR9FnjXvPW1DYS+QgeEqXPKGJDBcW23kwKiG
f3WBP+o7q+yitvTI1BcmdnKs6yHaQxFZrH7zLJlAXo/XdmjyJiv7yENfrRRrjsxw6uS+dBage/E2
o6/8iOm749VrKAm8iQk3+1E7C1hznSdea0H+PADN1oEBY4SLhEEDWwXaf7aNfKNF9Ot0LC8GseeG
XmvzAGv/dirx/Glgp5+XOzYQJicaq0hfA17Nsony0cf2Xpxy78V/bbmTDWSxX3L1DCJ5mkMg+nMU
Bo/7VPcsvH0jUw8lpGKjeetT+cNGYauIqMwcjpNBLlae3SN/PjGRHIGykMjBJIB6Qq1aH+YVX+ws
BwTruj0w5J8Tmslfnw+EQv1wQBMQRnh3TRjRNunhg6Sj1mMboUVnI2WYunpM6MNGthUqfwacvSVc
vf80qmK/pkrNg7KcLITlJsU0cyd/UlGx55fQ/DtQ19NoHfVQe2PBTrvBwSERXFTl4/ujm5U7hmJ1
UzqsA3EZpvLGQqyXkR+qpos3vNPlLBsdz6gnAl0XXzbdzZ+zHW67lEpiaGT9M3nIo5clYMPJi8Ea
SQdSJmwxdbKFPT3BkneNsWHkLF9Enr+Fopa0tVro3iy/63BLwuQ/ahNubFD8xYtw2EEjORgY5Zkq
D40JXo/1VYzjHVzCSZP0DqV4OFkwb8rdvOk0ci1VpxOmC6aoxyzjZoPdqYw4/U0y+ptf1QhhsbDC
xRWOoPLIdx/dXuprVIs4agdtTjpTVUsUZ7jgGwRbZ7SThUJrSUZzczp5iYb3DmiACSJowd25pu/j
ZH4JCllIsHvc5SELCSPqD+OpBecmNhMwQUkSfylL876KtkM9OhuMj/8LN0gREyJq7frv7RE5moDl
uDqTQmtJtfNejqMUCf3XCjrA3htzCgIPaAGK6NJrS8kp3Hjv10WcqA5rilSbmO9i3DPdneA1gE7f
glNagucND1gpONfBl9Ic09EHMb6tHgLIZuPRUTP8PKfTYi3yNL55uSnbYq9vsw+TAXnuuxqunN1C
9k3+4OaL7SlgyDvSdtilllcoUO1patg1OHlFMmS/8PhT0EKhVt0TKL9PtagIKxEb77vDw3TGQ4QG
kC5ZpyHoSVmwF5fyQkRc3TuSNpzrlQbtvxkVEDDoEAIOoGVRF4cZSna20u7A8jeKlDn9ijVpXMwZ
tQyU4TUZFFgmhHYccrKQU3TcS7bQv5dxnG6E9jlCir3pxYmcIAMBCxpp2Vr77QMoP66+KNeOhTR1
I6uozSOw7dBlKb3UGrLDfrnr5wI7pHgSN+lzFWYaqwTLf42yuD11yKXvuN7y4KpD+Db4PtUWzGWI
PcPQ323b/vaUpl+ILSsEnQuBLxrKVacoH5hfPPqi4G8r+W17EKgcMNBFdwg2K+regvOLH9VFuVKt
tt9uJyB86lO3FWrrNJsSweXPQaWpUYVUNLFLB96kybipaOJPUXFrCAMfMl1KrNtBnPwAPnbAyCI5
BsGRPDX2x6Q6cjQEd6gMOB+i77dLlMUogsbYfzOsy8kLZGgmLE0U8Xj2D03mXYVB6yqORpb4FWFt
MdQHbbqWFldeYH90Iz/Pgjebs4MHG14oB1cLNJ639QHdBmXI1olMJ5u1q8WeMp1znkP1U40EUzIC
aLMhtDVoKmQbJVx6sunckY37lLT1tm+pe9OQorwJAbefMLbe6oIvVICqxvIUU4Ra2RUjI+e2m6D9
5nbsiTd4fUmWdpKasCb0hJyBW4LhDIU0g8bQfZZhKDf6feWo0DvGLmDYPusARJ+QUkSrpV1HAsQC
EkPpW4nowB1T+/vMRp9nGOKvAS18pJfSV3ga3bgiQ0G0wSwu3JSPkTgwOq0Nh0sR/PqrgxBgiQAA
TQl2Sm3JHz22ww7tdwInzytc6dDdvlBXQro9+bylBnZ5U2zC1OidR6z0isOizidmlOZtoNnbb0LW
qE0XMlwwdv7yRYrhJpSvvmue1PH8fXsX8W+sOO0RWM+HEkR2U8tHWew1ciDr+L7g7LuN/6hNa3y0
3hhmawBCt4FRPVUjikyLsnKPDyr9fXdiDSjVaCxBhf5rmeHyw0cJtlXM+GhoCYVvJAQuaZtUpr/A
xJ/G0hz2pDwz9w8eqYuJiBXLHmnxwru6/ut2EHA7pn+SphaFbIDhRg2wzREhWido5H+F6MErwTZD
DDdDxEuWy+vcG08mllyZ2b0kbS6T1akV+nEHM1sCT7D9ovwXmNHPPVslNMIPpjwIZY4SwrDbT2L1
5GhDD+RQKjm8TMSC6a3Di5fsoqeWImuCB9BSkahD5PKN2OLgpfGE+nTcPYUja8t9qGSyG0sKBp8n
NijAjBNswYURu3WLnZrO69gPrYn6FGDwYUSIwbkwXkn2TGI2IZ6Fyxcvh2YmMXyWyAUalMEk3mzD
odzzOgw8GVeKM0Err9UFGj+raj9Wbk0fXzuNim91i//QtblWjrugimnwKGftmj65UbAETY76qM4h
TeUvq3QlXpnfv9qn3zxQuTMfVMieRZBwF6ElhUzjn8kkg9bFdIcwqF/tBbi+PwJX9CG79Vg3LgSN
7heC1YveFU/S8G9ietVMykyENneZZNLGTktmQpA0NCCiUs3CDeV1QS2ADIO+M+Gk773Zb/afNVb8
9LWUENkpLfAODmOeIyQnQvLuyxgsIw2EzsVyDO4FItvG2eOnPX31wyW8gXUfP39xXUZdbadN0oR+
Gqhr2oHv3w1t/GiHHFRCFE9iIosPqjq/Grq7uUZzQgXG+9ag2j2jq6PrbV0q5YJjl9TxhY5ATDE6
CBUpJSuCkHhxxcbHvkgcVMykP86WsaC8Tt/e0oau9KOr6DTxlvkvX+kx/NPgrVrjuLPMsxwWOWrF
W9tNAgnoV+MD+gN0PT5KabOwNzMquaaUBo/YbPwZRwpUx0BwOqs5RE1QH3CHgeP/YfCBmdldEO+y
70lo6qLd0I6S10AxT91qfpIuASu2VBZRm/s28T7KTY3VJ8txWyOjCdKtAnAva6rzV9+oqecFKoXW
fMdCguHULRcyb3gsISVCWvdmV2pLQ9+nRKknT1mRB/jfLzR3qMFba2I6SP0D9rNit4IorWsdDGhB
O0Ln8zVoE5G220yLH7zh8JApoCig66ad8bari/i9BKgIqWSh5o4e0W2T01clsXJAvJ/aAA+F5/sZ
hQnHuM/pARh2wu3Lu50ma8KYXnPXycFdbXkxA3CT8Rjp4CbidjSJvRiz/aX0D1ijLCKq1Bjln8Y6
CfCzlgcSqFirAPy5UwduaYwg8BsBOBwdvdjLdWIE/pWDRO2XRJ+QtQcChXY3TEj6SPfQt2ORQjCP
EDRgAk4YSAf4dIZ4rLepdPe5SZ1iN6YmjKgAakSPeB2bGSOd5Ado/CRJ0lwGNrd9ZXhgjWWwicCY
Ojxk+5F82ia/8xVraW7Gr2oAWmXK9k+KdO4vUu2ypK4mlKe2p/RilAebA4UmYcJ9vYdeTxKBgM1w
atIB0KcXM8Uq8a5c6rrTFxtKMymW6Hi8Xc6fKGYOGfN45OQULofMnJvLoBwOuz0BXJi2wyuEwRVn
3oGqU//Z0/ZgthM6o5awyX99f1iQU20nA/fkW89UFHoE+8VPaml6REJfbAzFcNybZmDUxjDXlYPX
Xe1QwfoWrlXoY2xduoNDmazYwT+snSFzDs6L3gckeSysczU2Te/THIGySgmQZirQZMvQERLr7hbf
Ws/V5Q1KCoMXpWgh0bmM4k3IeLlsJ872n4kalpLOsxOA6DJU1HIvGlG1uGA0MEVXob2FKKIyJTgM
CASE48E2UdBNZQ5wW/Mxv/ZXR0Qf4Y7y7yrkmWcsLhYFtkPNqc83M9SsHu1Dw0+XsFS2Cqg43wES
/8ERNfeYQRKwyNdFccGst1dhACHpb6mVddq/ib5I+aJ8AnLdF9wcDvpHJp6HfFkA7u9KiQv7Zzg0
x5IyfDBA23C+2xVpWmQE4b0X74DDNnGIhm+q6zGqwHsQ9QOhuzIeOsv2TzIH0Kd273fxQ7ceOxca
T19SCzjE/BM3ADgoUIOOshDOui8yuE3q9dNXroyWDnq710Mhew8mBGftvtjUbQ2cAMyV5dq/nr4o
HV9luEtWADpW3no4jMBJ4cfnYRjWCM6tOYDGSQytBIf3og7rW9MR+04idr47kDYYKeYKGCPS/gY+
g463p2FUrg4TBOgKFB278RlzKQBU0alXYugNBFeZ7C0f4kK67YisZEiFyjzYiJOHyJ5AQNNl38hQ
ciTHvh/Jqvyy7gumXSZYMkxYj7FMjXs3nwolu2FxBwCZBKxaiFyXNgs8WXzKquZBbGUc5xuVZoYb
jEx8QWzxBwqOLlBbGS8NThydCn15xztqyPPdT19MI5Oj9EZMfTgz5moDkmb/sai8AowmNw3cbpoq
Jw2i8CDS5QHzGFwUXZZnvPjxqCCv879DZd3B5TLcAFOdRwR/eFHFxWdU583osTSw3E0qyV2EgLDQ
C9+GLljpT5Y36cuNGTmbPHli3prfGfSb7BTayzaMSUQ6TKjvYICRhTzyOpE1A1Fzcy1P8gksDRpv
JftmzecLpAiCMty/zkAManYnNc13QdhDrODSJrAekRyCFySUk8kIQOqRkyGpJuGv8RGmczqc6Zhb
ftiresyGfOQwuCdNd91RDmBt/0PfCydiBvSoBoIJvbQlHl8LzA6E/HEh9syXvzwxSpMHsQ1nv5jS
e8XmBn1M49z2lJcSTrxd+x2aXiLnqzSOoFtlnDGyAVG4R8TiDXgFqeSnqWUmN6IJ8/wmwCz/HJ+T
IEiN1YNVrGuUWLviV7dx4SmpLgAWiEibGPuBGPy7Yme9nJteVdQ6WawvsYcoFdQpp1fE2xoSSJ8M
iGaKUaeWsenrUbJdOQa2a+/nv1tqa/imICyIZ7+/2mCfxsY0OM/hgxAr76RRZe+uRoLNnGbqHwh3
98bD4I6zST87FIQBcD3Dn6ig3Z/CCAb3MrC3reJlIlOKVzIXyfvNa6gL9sVsLuwxzkc3pR7RgI87
AHkaV7jiyza943z80FjtuS8UO3rLTQIZOWwchmlUlkJoMRVu8U7voQqiZAYcWXp40rcZZjb4KToI
LjfOjm7bPYoMFS973uMbP7yEIOUIgyCMmaEWSl89E/TPcdLaRuo1bEczqSsNuimDwANb2xLuaGgi
D8KiQWfC8dI3bXfD9Zi5DnSBGSfSPV2XCl+TrNwE/v8c5xMxfx18yzrv1I2FsYjgKTP1u481HVxU
U2SGWw3Q4Ac7kFdFmm3d+7S83u9hwwKiogCweJNMCclxAeffGqeEs8HrSlQKwwr/WCgt577BreuP
ed4mNoQARYZOt1G5NDqmsilD7aWow2wFDbkwrp+UnX9Fa0KaznnddsKugbBG1zDPIsqRBpMeWH4E
8IR/DtPiwrTAA8g+eoAmvqM2KVteU9fDAOZ2wZxhzHvDnmYAbRR/2Mi72u4jaTHHXuOjWXLcafF5
2/9By6GbOA2V3LTl0f3bKcKRHw3NlkOVUjND75V6fgW2v84WLAirf6eu0/dtJ075NXRvbEi83RQ2
ZzFc3sRsHvcuXFrE5q15eiIqpvUlddYuajhsZSpiYvQbdCJZRicmdryVQvJDyMAm3FQ7+iAIO9iN
kuUu96+jmoh7XYN7tBhk7lwt/yqMBA6LzIGfyarDZ0MymA7/77C7O8MV8q9oulHkfl4fBKD2dilb
NIo1URKhcZm7IRL3TP8XJdXiN9A38JOntJa+x8yF84ebePWtgkXu7uH1mm43k+KNPtJObJrJBsp4
ko0usYQKq1i6QUyvA/LoUKRP1umDULuw5M3IHfikCXmj5cNIDZ6t5mhXjoz5BHD3GGHEsWuUk544
6aICO5uKhDET5sm47HCDPUHO2qlxGQmjWVwZo2hWPnpAdbonQdbMaDoy7LBoAbSYDdNq7HyOmOTE
55QguswIswDVeTpJPAkIPUeRZi1ft16hgGtQxvMZw84rWe+KZY8oLazvKAyhaCBd1oznU0qkH0tQ
BF9Zsu5QEsM+qLwnLdszySMf+4M7q6pF4BDRKQ4eB/w1LKH4C3hopzXDDaWGESVcJGpkDoiU+UGR
MtL5UgWpvDfwOktSBuq36l20BapRm6+wtSaX9D2XeTwg8Ck7dpa9IHaN8oDp+A3awbOwP0iOI9I3
oifyHEToY9NC1Z5f6ZG06URav67lB7/ghpjAAy1qAZhx6fKRr+xTRSNlQP98Fman1vigBsXeT9C+
NeXQwm2+h+SRF+WP9w7EhutwIbWjFw9JE0c71L0OzCJ9E1cIxz5jV440gzfHQ19Im2PABMXvfA7H
nq4ZWc8kccj2860ppuTLBb9m4RJvmAuuuDNW78wmkPWQHJ7CObQS2k6t1/GBoGypfhcM1uhzcgw5
n9azLAmfgWwFuokzoV8PafR+/0RJONgFTGmiZvggvcMMzzf/GVhEZh530ippfCVVeU4CUzF1gaot
Hys0daGze1ixnV8xoMZN808mV/du3Un89RVl2LJXN7t2414bIBPY8cVg/kz0bAN6K7d5++MpehW6
PRGDa9p/es9/usu4G5Tjijp3VLzyaZ+NMjHpkylRtHizHy3uDC0rNIR2S0ZMLUpu6xQg0zstdX4J
uekVEKNS2pH7Dk8KxYYvkHObRyyIcB0Qz4rku4YrW4A2W3I/RnzBObG0sBrzI0zTNoQlpEcD+Luy
6yQdciXNI9Cv7SisHnzXwAbl8gRbGLHK5ap9DSRPVbSbltRrhWyLJXn3R6xs44zcR2AqTxgZAlZQ
jkF7jlSXqh2U4W0lVCvEn8M/7a4Z2OKzWwI4B4RnlNhMAtKSwDH7cZRc3EwKmVgQnu6Wq2NpEp6B
r4aQtPqYqBYTbQl3vh2uWsLeMLSVwFNQ+wkDZRWZ+UTlRPH3aTwW9sVnlDcQ4A6k3NS2+eEIvgpk
dd7VUH0XinkAbPeY/y6FFRz1cNCjONBEnDVDnWi9kv6P2rW5fUJ9sMrfxlfa+rQ1uxJ2Peux1npl
A1vJyfniQAuaxBh9IITkAxq40OLYEE5kZCiT8+nfpz/yainTl+kXCXdP/6q7qt5iJRxz9Zlj7G2c
8jZ0R+kFDSNDiA7jS5LxqXsxzCajceHRT9HXZaVg3wclBxZXZb9YbML7z3uUvFnxCivEaA4KRq52
E4TPK/EtMB5KHd6Z+2pLjOEm+j51pb63sDc6GiHChXfkldr3cihmBJK+Fxuw6oRD5Q43Rp7/wAp7
1eH3e7b5QSJfoTbkU8BnTEI5Yv3CYqN7LSYORx5XJTpBa2yW2soj3PYPAfBB7/3xU3iVE8p4uIaO
NF1wSYwq4LtQlxI5bZXfWUVxrKHpTn4bwhgdrVzRSry1j3DDy823Yryg8RQGHg/jQmGysHtRd5PM
OGez7j3/sWI/2BBiew0688c9a6izXzfa1CiZIf9czWi3Dpxsa9rSSnVNzpgrwvEdScj+HdS4v9fL
H/9o9MJHWo5cOPMLPCc3Mu0LdvcekXZYY985bapd0fjl+QaZSkdQTssrN5cpimZ3Ytka5z5airx7
oQD8KMLUwfup4aFl23HHDII2HeEyj5C7k1e5GxNz3c1bCHnU2AySx+dEJHLXKULyjt5svfIUMla9
PzglMbVUJTJy5wSlPi4dUTXxLLpu0GcLc1FxTiapXsPp7oDbQcHMEIPpGOJhTOG6W7wu0UQyxQ6j
xbivQ4muvTjg+MKtrbZqNG9dEFsfT86kDPHudYw2MF8TjkLXFErz6wAmZYGFlDMwrhxWu0PJvQF5
fxyyuyTcEASpDYNKTFGBZJblsktuJuKbrItAwk4PfGITWEmZJXjHowUP7hv5gpQvBHJcBbY+18uq
RvWgrxWVLksUPpAt81eQtJpiFcMS43V7UkymrZFv/8gK7hJfrAxU9fzCUNVw950gAr8SLqwLgHU6
dAVFB3LU6QgBHyhQfAsRylXmA6eOif+ZTIo0twA22gEPunci8AAFwCstxLaZJGbNEGYmaunN71bh
KqCEFPr9horNKVR5aY2ecFkJYduylF69uKUwn4KsP5QyM5s/JW/aAazwkPgp1b6ZrbLll4L/hXGU
x4MfxWnWrjeyzGy7PntVtzOrHCDLsdf30dVxCEY093ephRInnn9/FD98ffoSGRxNGUTyijMMWUqy
+9hXoWNm18qE21/8/hJnKQaD+6XphR9AsDcEu/Oxbrj3m788LIF9mdOT5LLXS8ubE5fx1bJlBysB
yuX65zd+0YddhgHDLRNEfSC9bVgeV/zoS0QB/NxTftxCGKJMmYCpBG2kohLVscaJVgZThtMDgd6h
D9GQ3gWb0YN0hAhcN47JZ6V84jeD+HNN+gq4usVlLykYsrC5BIlVMPp33BBupDaRPmRKVDkM7/we
KF9CWKdWeVk8kgahh3KQ/SArTaEiBu83QdwyT8tGEs1Ex0odayuN97hBolYrWlG8SmLR+mJ3sEby
jmoCyh+wsd2DFHKO909W+AN/ZH3QtqkZUbjEbsakQUzH+oFCC4UPFaLha5QsV9FA727Phy0h/HVs
n6VXbOgJgX8wANTdGjGXT2Rc6zvotjvWJMEwhRi4vmKoDCsD3WEVAJwEFBO4F3zXlrvHEwjpAg0Y
rd1r9xaW8v2qpO/jezfQls1cej5ktAXttl1Ltd79OW9QO0zj1ZbWZwrakRqFKN4/FDGFeVVeG6gs
2R/4boLQ3WbRo3og668yay4qCqnKvT7b8BrwIbUhlW1Ky9xYJj45sju6bQqPFygXUPEGmZglu7Kw
gFMhjOg9dNlNyWrdXDjCJrU3Qr37DKFebHW591Ow5X/9voTKe1TYtTxymCB0eaQ7rWMfSq0gHUq1
NlBFL5tjMQuxjV4YaniIvVoHQciFNEljRnq64S5FRCVl8CvJZX2ieuZx9qwJzugytpTDLvGeEQLz
b0fFMCMVRkHrBNYc8J+p12kqb/P8ePmnY7yGv/QZ59dW5bJcNERjwGkS/Fh3Ih0LdyqbSqJjd6TF
Trn+aq5Oct1E6ln3TCMzuqr6eVFxq+r9zzKZLiJDD7VnzN7WESF7z34oX/s3xupTtLHooYXrjplp
3kLD33RQMdFnZWT91AXilvPP/XFYjFOHEbPBNEF65zTBv2CEdSiujOnLRBGWXkeyu+HgAt+5mAIK
xSFBUkm7D7GHwju2bx6SWTPCp40lV7yLOXF7GJ9BWfnj76byCHFAxlvyhxTTKBKbxFRSvPy7tXvJ
wWx9HSOBltuT0AgQoMZFBeRRyFIsa4L2XWPoytoODbo6jTJsoHYcPjoaIekN6HojeWFyjOmt1aqF
oddWIIckNC6aOqKCK9SJUhIoVIdjM5nVPpFFxJnXxD+ZChi7EfFDyQWiLk9SbLUdRqCShX12Pknf
v8iEDZNJ3qA9gAa9A+zxxSKcQc9Y7rq7WFBCnlK/gV/9KF+6CoL/YCB0P3JUaM2HphY03u3NTOWn
APY7fJt7cp8+IMC8eQohQiTcR2fEoDuh3o0IYzM0EBBeZa1U7Z+emBnBNK6wRYBqbGjJ8LrA6QhP
osnA5iVEDIjy5GQiPXhLWoXNs0/YdHm1hJcGgi4jVRvbpKP61PEbBZ5cDLYLNkPnw+2WwtOi7lQL
iRyy2yiHx7bGDIqs+Bide+xO0KE/VItE8vVfSbMrvbxTCtL9kDQ9kpyFKA10/RcP6Ri4SjAs1gn+
N0yJd6CdCL3DSfCBndCBJyUspbjq39isAjq5b61chx80cL9uQBHVwQaEZ+v4fWZW/aEwfecwsJHq
W/usLAtGd1GvEj9CLTUuJQmIkDpFXRbRlVRMazfFO+pMbsbu6wXW9dfhGDdb7qtcBtMM1zHt3G06
ZTaY9lthMwXqrp0fscb6OG2mR4AomVuNCIVAgV0dqGpMMuMhkrcaXDQQaj5PFbbbhrk7xLuerK6Q
wdLhrLyH2PGyTnzpF7pllPGmrI4ySOG2LAPufbSrQd7WNgzSHVdSrI8/zMvkbvC20gelYvDfCGbb
urgX9TAVnntIlqlnG8rHkxrV96DBFSbV5Ol6qCKZttFGsKejALRliUxeZO2zF9caMQG4dS/dP9BM
dPHbRPH47+yaRjA/QhgCaCvBsZafe/4PnTl9F8b5LDnoU06mEb11+4c0SN075Lf7L4ZU/DVk6ojM
hWQqCR0GIMa0Ro7x58AaYXLsNliAruAezKsrI5fGILS6mCGtMHKj0pkT65un4b6DJ5+WrG+jLBJ4
AuIg2RBLGI+5O2xqKiv1g9/gBZ4zIQQjzNbHF+ECUak9x3O3JRF1aBPDxZ87CuKCH23rtCoGz1ZB
fPDjDJ3b1Ismi8ufr8frbRTlwQx6OrJX9Ws3J9k7mLCWdBPNofIAHB8F6gqm96dcBB+DJLKq6rmI
ELNyOhRF68aMAkBq7MOTVfsdLpqm/JhdL98di4TRlYgoPdqckuoPXdN5I8XAJNZ/GYu7o051j1TQ
cej+fZEWny6zfKBtdyurMtv50tILFUbZQhoolbcj/WdaXCUOkYnzVQB2Z9RxT9Koh/H6hXlp+v+l
Td3zoQ9/NBtwqoUSn8wmcLv6J3zPrtEF6/gMDxf90HVkTFEbNOgD5mlG9U5kX6PUk0CQmGjuIVXC
SQkJjn6g1L4HR+gvNuxIfRSenkDOOm9RDWooszDDw03ZcuPN0CA1ZyUtAKtjzqO8R0CWtUrvYsjS
bDIcAHfkEq9XeBjs1Jucqz6vTsSSOmbCr+A6VPOwveNthI6hz+LYeiya78WCNxsj+ZVcq5UwKp7B
T+LY9xdOc2M9lPh9QXMGnYv+pm8sraQWZD2WTah6h5wMT3EYWzVE5pvfQEMbbl3HbEy+YBkl8F49
MTsLMOKftBynCHyR/s5yxiqKM676MPCagioVL7HlHASRA6SzpmTiIFOfZYaVzm73CJ3/xWsMCqOw
yc0ISn37iD2Z3P8L7R39tvBeGGnhYrCETfSwLKGSvZdpseVssopcWyRKCZBT3ubHbu/pAo8yo9OH
VJB7YFSHr59+DVnZU1PVkGeFb+oOhW+fvXL8hp8q5hZ2yr7ChjMA+Vanbnqp0E8pEV1zwjqsRAn4
Md/ge9g9NgxVn8L1guO/17BzA+fkkyBrdz3HyOqJkC4WHjpxF9CNq15OfjglefMPe+Xtt5cs4oBv
/X5MXClMMSm0et97pclJX3F+MpCCsm60kj1aRwhybfZq/WiGTksPe9G6ykJa99ffZfDDDXa57eWT
o1FG77uGqaV9ubs4rsxt8yxx92yVno8BlGE2RbGQYR5TQk4Vfymm/R5LIzF9YyvJgwR03XFwSG0R
rj/YsrjOAVGSYpdHpbZAihNewm63GGti+rVFYAZtrrsXOFuTa4LExmRGKxVvCamHIYF37xC2YHwU
jr+6x37Nu/YIhKuZq/QTnf/eGDeiJi+/hcEknVUQldV62ZV1Co/ADM2j0t5s7fBlu37V1pMkZ7GR
1cEetdS4Zu6DQZ0ZkkraXXx7lqcw0Y45L+oneRaJ6asYaLkCxUGM1KoR1oU2cFy5XOXYImNF2mRd
zC2NkpDST76LMZz3N93RsdJlhMO1jw1q4T6m0NldYcIUnnJv/RfIir1dBw0MBjR97hjkVTE+ciu9
+Y5yZHYW1iOJrcWG00VHHmQzso4lOUmkIYiB6GJWg6PAtkSmrB6cRtrB211BRV84dPxrPqzrwPYP
EJ0h1VioeoXrCIXRVBLnzjcUpIpZR4zhHAk6t4W2oy73batSOt4mkQwhJxZmrX8SQb6AINIDCdK1
wTPZ5r3Osw1Mv0wsUs20vOHNp7R+Ks0aNAfUvJGJa25cdA8ft2u3LI05qikClU5UmOmwfPXkeDSo
hFeD4aYfd2nZW5xBgaDS+D7ux8J+LECGCBiBQeyfcekEsXO6BeIRYcF+a6dsGtBr8gqU/tMBchJT
823JD5YUAk/o9+lUWY5Na1Z+lbRiRO7ue8Gnqi6iaYNvu3jbPE44QC2P3oKPHcdUGK6MSTF7ZdiG
PS2+lE4ZJv+1Iz5CDBN/rHoyD+LK6BfRIYFCiqDKKH68xTqe4DNKgE/MRmS2mDWXwX+bzJLaNXy7
AOmVgvfKfKVX3FK2WHNWcWc79/zn5ptBvrFKrfFIp0ZX+kIubQZKYUR0nYzGZflMw1gndmLgdMn9
rNI+0GuUs6+8BbhXPrdLXW13P76hFm3UUmhF/QeC3wIwVB5iAhRxZTXBBDjB54+YhB1mHOH/QJfJ
TdHLFfmIhd7NCX4VGEz8Og5e6UU2QCwDvSWB3T2V6ytNEzAcEdPoYHatOhK7u6rH/jZAmx0h2OTF
KY3KrEL8a2zm4xtJbUPdJjOX0XTQfOJOVNtPxUKZKPWPk+rlaRxU9vZyXM75jtV2zwzKqkGj0kH7
EQQ2+zZHuBmQp+d55Kw4OO1IL6rOe+G3rGij2igFd2XT3ImODlxfbNibcQ0XoXKLytnacOp8Kjsm
suISA9v7+NlJxRvQf8OI/Zc8rOhW5oO/j0gKaa7VShuqj4T+TwD4f0UEFbZ4Pzq/3RoifXMKd2Mq
g7INCtB/OPVeKFsV8F77vCh+1FgFqlZsDMkK7RAsvgYqHtzEtEuZRBYO5p+digt3CGsMvmU0C8DQ
UYTfMEYh8xs6DRlk63GYtKWcOmmL7ceUYC1k0KP1l9hCLY1/kYSPFe1ryjD46NzMr/CkUwofB3xf
Af3VggFFve/0S5y7MoL/uwKHKNwHx8HV6GBajBc+7XxRQSsCyxGxec2hW1qsKO5Ei2kpphgU+E2Q
A7Wnmiircr3B7ZSsd4Qg81yKfWWTEVnC8YNHeIDn+DWKLDZyrz13NC5WtNkUu/T/Pn7c2MT/2ke4
OxLasUIQYNUga6AApNWaByhcalo+dlXwurkeMJoeGWComyVzZd5Ak/XgMW36PqKfmmULLFqpfKcr
gfEJna+HuzcIC6V7K+h8EASZvdDziZ6Ed3eksPbh0h+YRqrBi43VA+YKN/BcI/rHbuSZogLL7vVN
CBqCgiXEoyWeujr7pM3ovfCv5NSaCEuBIHKLhvWbad3+ozCmDAYTACRShNs70wDM1wSoOkPt1fdK
IIQ32MGCi/VZA3ElMDrNmGvnPdRZerTamTAEtSd810SxV3J/gedfdnktaD6I4bfZqjg0QHGOm59i
9PFBgGy27Q0pKGE2CwNUD7FAxT22KTB1IX8aS+4i1zWJjEYiAcVkZAdDqMPu6W1PbfPO+W5uBNr+
ZCRhWE5FE2wzFvXkOkNvPiMAGp6l3mac9DeZmRS0k6G2yZrOO27aMCqlAjGePxtbL3fAuMwOTfOh
MNsLSvmV8+a9iOAq082SGJWvumVtai98kncVFUv4XljYxzpJH6B+gdC/X2G5yQCzfcdv4YrPiz4w
nPVbkt+HCTtoHllcSdrjbQgXmzFGA1bjUtv4HHb0XPx/siM+nX70uNT4ovZnbpVlLv1fEt9tAFgB
jbv9Vkd/nKVycyNE5yevO0pfkEjkhZKApD2JJNUn43E2TA5B/QlczLWB9yhjpR6ux2ZgqFNlWvt1
AzWtJHUJPqnFi3wpb9mJe6tqwkVG4ceBN/wLhUZTH38VWl/jX9UpN0c6gzrdmSaK9d+m5bK52YJ/
tujmossPi9zNaieenui3ZWnpMNSLr+X3GoVJye4amtI6TM5diJjoiQ/BndOGYq+h4/vty1kvBx2z
d3iO7EIgP+Ap9S7p2jzln7Koxh8SmtZd5vxTCIkNPVZvpSb9LMuV3wNBC3GHB25WRFS50Y3+yA9S
ZaLh8rAPpxiw7YUAtdWRfe1Z7i8jATRhECZGh5HeL3nlbIRJkVd/NjIh8xDgEOffD0Jfn9DwA/Jh
TK6JoopLpPczLwT0xW0wDzEZJWiIrLWtUfgluxpmQS7fhb0WfZXcLWAAkPVcC8bCnW24JzkkjJrJ
V9+AC2A1DuBAaflMh74cOyQyZ2MWI50cKle832LEJs6FEjMXh6Yq7rIDWj06nnwFDt4BWLqYTQU2
GRvq0bSlLbv0m5KJpVjsuI5mxgYqu7N1l6ru0m3+YFPQT/pgYdnsaNI9j9OaMex/01WSmEVCyxKg
o9Xq0JoniaCDo2bSkDtyLAAtrPug6NNUA6/E0RWwyPTidApze+xegpq4e3xcZE8UuWk+JODykm1O
AZK7FKC84WL9IJQDGQFtl8hm/VoSoDVuMr7jfE79cfxv9I1DsHB9ywklAEanJ1gRa8rMcvARfpbd
hQmJb+6aYnQCIO5K+iqmn0V6IeiQwJHhQvgiNQvKuPv2w9TMoCmZpTeIAbJ3g/FKhOQLC8auBZN7
gh3wxmBARkJcDhcj3IXGYCnj3iDj0ZD8dNQEHI8ZMdAVC9WjKvz2VRH5pTmoJTNs178R4ObYofB5
1iTHPVpp6pls4E8gyoL79dIXNTS7ANKqg392rmA+5H8SA6zovDJ011BdrTGlOwoUX7YtyzQsfxA8
LNAq9eKwj7rlktd4ZkPzmW/2pnNW2GeXD8/s8Ap0gfydM4ZesWGVb5Gg7NTXzpdc/Gzittx4TaDj
jPpsaKa0WAKa/qz5zFDmoIXWuuDUP3/Yf/65Ayh5mo8Q8rbSZvjlBM5HEYyLDadTZMt6X+R++Xw8
TxaMLMtUZRjjWC5cJDyuwnyCWTeGH386hO3ItoMTKsuCQSK2OHQxQDRauV3+Mtc7q5abARNMGOJl
ppDJc1vtyuwZ6q0pM8wvY10HQg4D0oAf6McmUFH5WsFryn/IYtJevrJlDC5oCNLH7Ctf0VuIutJN
9UprKa6Bwj/igQlckY49BAOlyX+FVRO11fJN/w+0AgVL7BgjQt/yqeS+PE2KYXMfBimzGTxKpSCc
R81OiyLOgZr+2C5JJhBJHVnonz/sf94KVZOOxX/SUOm98+/sbvY5Z3dhI8pcddR2BrNPpSCzCGpR
J0G6JHvVmvg8HULwZzsljAWvX2LiJmDrt0GrN2ZgsdLKMDL/N8HWJMRhlPhXBu5mBTOjvR6O0Tre
uu4HNgkXWuPPq9dzZu2kkgIsTwAn2PoW84dVrD/HdXAgVm7zwqz06waJabYi6bG/7SgwKEiDYEyQ
JIQClVG+kGRdJY5uAnZtzad9MqAVh4fZE532pn8iSoHS1wIhHdqhfOSzmoRnLeL56fWigRuDhT85
o+CX4PAZuU1gCILo7WbP6WJl+lfCBM66CkKbZugMKCHxaYmgZHcTIXooTDniIPEcAAzehFcukos2
IwQsen+KNuJi+J2vdS19YzsJpiYsgoad61czhq7TtN8d2KDy154CloE+FZ7GeDrWChbrX/3sceQS
nsvXUd90th6603ztVdR3gh/kO7Cmh9PpMzAjZ9G/q2oSbmiytjoA0DFZEbeBmT32SESISnKL+47X
+44+wk/Nci46r9uoVDSwQHom1NtTlc+RoUXcFAJzn+F6xDA9aYAm3Kn//rE+pTiK2KhR02mL8TAt
ryZ4awYnrq8gMEsNCjlvlQFm9zBmsVHvvWmUSLg+Rv5POrr7o8Wd77oORTqXB3e2CgrsF/Rluxlt
czdbs80qIkygDE+Bfojah6pwMn8NEz+B+akIN/8CkoPJYSd4/zVL20TxNp6Y9zVAHDP+HmSmebEo
9Q4m5kTfKMECvP4iD5I1s73B0g6P8ztQcnKG/OXdNG2dPzI/fxaSvwW0SOJeM5gNLh/sY/862agd
mYzFwuyxZBODcCC3YwhXO/Y9/suteRORviR+GaTdT6zh7LRLFHwIBdGlTQYtdhWiOxJqIKEZ2gos
rER8JZfEZwltAhAZ+CdqJs13TYIn/m3Y8OL3cQEpXMKaKI3XE4SWkLIFPuhQuWkqHvR61FgLCIql
1dRLO0etGMmXsqNhDcCn/SELrN1AHIcTD4FVd61Kjk+seKsn47wZ6C01JnUs3oyFaHkrj0v3JC4T
98vUFekpjNFGf8n1I7J1OY/2SWsTPuPBf3el1ptwufgJv/2cnj8/xYvG9NLRO9aHRJ9GhJB1JrsK
hTntGztYz/RyK4dr7NeAZseuy443YFddhOkbzo2ZyZwvaf7s4tsCoIpx78z0uphY04oX7RW1tSf8
vvgA4Bux76kXVMcAwIyGLeR8UC//qzuA65HbkRV1wlYopfJNIl+xnaa4mPOIE98gbh6a2QqmNjCs
aTLT5aGHlIY/bShHvJ65EBlI5wTZGWdHd3OtkDWW9npnqslHkRuiTGz6rL6HASbwWs+a2m2ky0i3
5Be9ce8rLZsIXqfU/LYA7BOE3FLD+y0CrW9w2KwyCpIqTv6ZCenRekiuMEM9fTuHMr0fe77R8vpy
F90gTXHEPUFyTXMrhINUApCN+qwG2e4mNhxo6SPiuudf6T8ClUIqBpIw/2zHz/rFv50fnXOxpy2b
oRMaiidyeKgaLhCm2CIv3b5BipqLNmbj+istEYWfm/Z1ckibfO5RN2OKUuzVccX/Jxis2L96mOvV
NzCaEa/P/raK80j5JFZC1LEi+bZiwBa8sq4KJKK7vNGW5kO1sGGpstHH/giFad3Uu+IjCOvChiHf
3mB9w5F1ugk4lXZWsW+Vg0B6PF6LL02S1tO/QA29orcx4hbL7m0jUKHOmhP0WMJ/i1jLYkdUc909
TMO3eil2F7kJmerBT8iQd0uUMVGHkdphgluOD/0+djdfa0VzI081YOnSZfoum8brlCS15z2fCGuJ
MjPV0l+Bc4ostR3Dn0ChYE+py3FpwlYeqfAmPKPRSU9JL9qEgpexy0R8LZdU9SMsaaPVTeTITwGn
BUJuw+ERtWhN9z74W5bTYD/L0aGBnNphI6JhWU4klmTqP5/5KFwmSt4nDkKdJjYlV6GeGccHpX5l
OTijwaAMbtEzRBzBLF6oalFqok7qNsv9PRGrQ2EeIic0Rf6jO8rs3MexgANSGa0OK8x8FPWT5LQy
9i07zcQSgLrLu4v4UJ+WYRIl8JqudBo0tkzFVtBnIhDK9ilZYJBE0roBcnp0b9Pr4ROLHJ6fJkCE
I1aEMK2GZcd9E+mMzaHF4CAzxJTYEbyup+eP06Ctphab06jg3L+Q1sMFsOiUrSaRfHBF+Sx3tbAr
U8+5yG/FyoY1OHGAtbWC+/6gY1avmM/Sxz+FfXqi387kzc3Zuj8VUtHL4dHROpO+OcCQ8hi45Ayc
fnp5szfKSHnTg+cMKiYvVOsJVljIOqIzcSdjpmCetpqM6AslzM/NYdBC2MaFEnTq4H/V1s/Zyy1p
04dyiLh0hfFFANn6Fhl87sCLMFEJT6gv/j0W4dR+ja02gnQInFnKy48kO71NuHpppkJs9v1SUjrF
sxOXtwJV3DwXEpNbptiifm55ylTz9wH9R9j6Twv5nanzKos/8kEIxjwC3yq1di3zKmszqHXXNh6j
0aVSgrNsqZC+5eI2GOZmremeXPjs0SuUq6drd0oqFuWLP6fJFNicwJv8H1gDtjA4yd8y+Lj0JKRJ
NOj4KC7uO0asejTVXlHJ2Lezpso2Fkq36FOosNu7j483Ezc0zlZONNUxB+7vrE2Aj80th8SAlO3l
Rl9VvwIXqQDFUz8ZsbvtSqh16yVMcr6wXAZS1Tpyrq8Jkpj8qStSyesrmUajPuSfmTQYHORJk/up
jI1NBjLzyraU9GfYYnHf9e8JhJTekvXhsKWAVNA/pigOKugyukmAGoxDYEeWK+nXkIIEJTyTSzSs
ZL3queTT+w+4MAtfoGgH3DZ32JDk7YSKihXJu6ZLKfa7HH3SQgAIPQZuv7yUSoiZN1TSfdeZX7L2
Rz2BX7en0vEt+1komgc9EHMpCNlwNQnnwr5/xH+13Jwj3e9Zk9i+rquvtJPgoSBwBM8UP94tAwtS
dTkkJMxATBq2Y7iPI9o4Z2QxoNQ8tb1BFvkOEQao34vkv8qJaTHiGwDN9gmA+hQBhtSMdwOGmTfg
eGgMNl0dkfp2EJOzegypSNAmcZpULSNNFYc+bbK2ofnJvo0cScTPZc3sKorBEyDSmxgavRXp+lOh
wGzsgVJfp3xf4o583rX2670avbEYSN6gTrTMRZYCn/4aCsq1FoteiiTOqFTDjuRgSDx7lP30m7DQ
oOhL6UpW92CtSmC5/x3/91+upSZ2Tk+It3QgMZ3kPGGkMjUrIMQo1ygPiyE6MmLUz3PPnBKw3TyW
ZnM2l128TIIQAR9O8H1+L99LR6M2SnnbfQNQDv8lzw1+MQJ7FwMLeG52Xl38o6wH+GjqEBtQ4orD
/3FctVpLKWa/FO+ZAbD4xAS9fMuU2lH07tpKObThUlV9OQF9RULv8dE+A8rfRbCUlrIRxEIZyR7i
VaLSckLxzYd07a5gHw7BRJjQNhmFII7s34RTda+IiVOHyWUSXx1vfYDI+jwy8/vT2fA4r7SfW/9S
GJV3Vhl1HyDtxdNJNM9RPd71XP9YEIw/46ArEn8YMZws0Ruww38UkA9btBmXdpTI5N2jbbEAxEuH
c6OOSRWtMg6vFwW5cpwsRIeC1lho0WX2qxYaaX+7tIBa/fgneuBcf6y3GbWCb0ZT5vIn/gt/zmXz
5u27uMsCDdzFelDRzQp+cJSxlK5koas3EBjt9csqTzQSe+HGryzcG2DqiQp6ZOofAz7A4Jfg1B9r
73/du86u1RObGbhZBS4KksQr+kJELfyQX82mkkFS/vMShuicUjv80ezBY9aHsD+mXtUZjQky8vea
4co4FNBe0FylSuoQM8FpYIpCjYXppmc6mc1wc/YsP26bol6ttZissNs533/CjPj4A09dCTAFpo4d
bK6AgyqQUAyCbAfZ2zM8sbxpgsYiSUEcLuRHS/SkoA6xA4QrQbJY6aAYOxU0uu3+ehKR4P/Y9FjO
iI9sGhTZcAGGrR0MUuc6bo8E2kOUfmwTIcYso1/VzfHNICqy7NTn3WwSutHOKJXj6LYterh9SGoU
ukFIX9896LIV674X/SpAYyWwqu1Ux63EOSJgIvgbpx6RmGjznc7k7fAZjgkO9xeK+G1em8VtI8t5
W3lGVDqaqGirOxcYWw2uo7zK8NEeKPrxtZ2LqgPuVl1S5q0larFp6kqzgRkEzUUIvB7InP2+kKXE
n0nLN2U0FF+3eW24vheKTjHIOmvSHD3EnFzTeEqCqocCd4tV+utK6cJN4a6pVnGf7y+wogLhLNP7
5xqWi6qec69Wig1WcZG8cAxzC28pMrV4H+rdkjIrHjAHzMoR15ULsgTOi+8EV4vAxPddoIuSYRoo
K5kXjzhIDqOHn2Tu3lfEYgsx2K91dhc5M2puhZi/QpoZvQ0vfYxjz0lFN1Q/eFdnrD1FPLWlXuxr
9zGM6gylZ7vLkQOYpNENWXcRxBct7qYz5MxbEvCXwwnBRgg0qwECXG1J1F7kBjA49wreCP/cnuK9
i/PhVvapx4EhaeeaUr4fI0CJoJ+NBrEJpZFBApwdb5fY+XKkYffnqnUQA2UAiquBKaz1SWuBKovI
jvPHSuIN10kkU7SkrwswFC1dwfEcqmKsOTOpZguGGAYefOTdmmbQ/vozhREbKLuVT5XzuWn1nIpj
avbtnULV/pdODfrEcFX9WryqcDPDBHSsucOPOBkgufyY7au2hEsuTuZuQ0dd1Gi9RnwnVTOnnQgg
ycWtLnSvvI06M8X3luO6ZsmlhTOvzyev/qrTEUq+yxOW+VHCxano5BwM1fVnDgXJ+ZywpeF8SWIt
ytqT9HGrb1EMS+B4qX1za4QzjrjgS9oLJz1LB0mBRJxDphUsnVpylu+pcw59oJPJ705YkS4VJ73K
1Fv8qrtAIEEdkJZ+D43oq1odr4SiODCTbb5oChcKWSloXPWGbdQZhKU3vZluaZIliSJoVh1g1aKm
IbVfBwdPxdXxICZwVMPmk/qCRLi77SC9eV4cFbXwpFp3bo80NsqfDf57LytcLySaGobKKCJeMYir
bfDnaUHh9fbQN2iRRhJ0h1j7JjY/dPB2AAa0z21hifsZnHiLkq4O8vGaYa1K5Iw16GRiETEWmM2c
jsRjTplrhhheAQzIL6dSMMU5bW7SBvnjPSIyQBGyoXE+DmYbgyvtWo60UA+46dKF7wDzKEaWQ+0m
ySumskSXl/tJy4bvDBbjNzd8Jdhxp9eehpxXYUWSf2fnDjf6+jugTWqnbj1sBonJdKTzC9DU2ddr
s8CsNMf8SvzsJgTiqzn2LVaABteIIsKZF53q7jhTP3HwEG0t1+aUgu2LdU1IfyiP5+GgFL3jySGx
4acnE3h8PxgOdpjDACXbSpSK+gwo32GopEcFmyZ8+ZfgVvVVoWIYiAPP+LR/4rlAW9Q7Q1fWx4PS
DoEUVtaU05qwEnjTJjNSefl7vqYQ6oGK7DOO3UpsCCpThtrT2D1ug7qG23HzAFso5V21TodOsrey
qfLjs4bxDZl/rcaYuzx39g8cUo9SMQgs9HB48dOYP7MR5LbwIsokEOJkSmuweACI39UghXdFcClP
Y17KCYoDm7raaZ7sIkJm54NRQGrYS3vhzOtja7QajK3iI88RkR/HfaUd6jt44rNJh7nXnXy5DtB1
OBb5Qh1lX/TpuYC5wHHsScoeejX3aruV8cR25ClgAoiWpl+hZsNXV4L/pEqm9+t7MdWK9k+kdGS4
/hTL7xi+spZuu2zUCgbnbtK7Q5tgWki0N/RNnqSSlEpnT41HF7dJ2C7GNjj1rFQUiQtH1xS/Qr7L
XIMXQTbGxbd3mEUHWlBPnCTDwAhrpjq+pj7ajgMnH1keewqByuC3LZ7EhZPpjFAS04YzUSE+QMcJ
J+9iE9pwKGjXYy5IWiXBdzkP9AOJw4+i1V70Zpzs2WyjJXkSXHK+udSDuKe9s/15hkUh474SZN3e
LNwk+iRM92nL2ikS6ZPHKAKI3drGgo0VaBDS/wMlY/uEp4BrdVlZBQUZ3ZPJr0tODVIlIdh9rm6p
GHX3yRwp6KyB6nmX28k+3ZCuPc3RqP61JOy1td7ExMmJBjdjuLowptA18ZP7KwQzl/zU41T5DLuJ
YA1/tUouD95JxRihkc2cysY6k+93IjUhbkUJH5aq27Hziy1v+G6r5vZEJO6n4EeYnTff5uiJqKXn
YPjIrSwC/4t3AZbwLfhCeVbKHQU+Z4Tvg2RrwHzuXEXzE56UGrpZuepUERKosoQdbjE3ovcCOMJU
XRckDkh66+HJbwbdQ6vvhIrBp7B+yeQIiWaeStRtaovxc8zE5OAmRO0ug+usuzmOaadGY/uhD3Pw
Qu8mA7Nvv39msDoDucaEMkKFV5YfQDkHV7mxBwtrE65v3HXVDWAB9TzEYOSmWR+7KvZzopOvd+sf
R6q2gwulZUZvxGaufyw2KYg+l9118POCf3vcfMNH6eczihHS0aSC/yIVJVDYqOgg9GT/1sHPyNp0
9dcPUnlSvq5/2/545Zryja6SiOkWP2uMxEVC3kWZPgxhFRz4tIOqksW62RSrVD00vle1lI60Ubnn
AfwGd2HA58Jp9LhgUCAyGQcJ4m4QGMirY69esuatNRbeRQwTeMKecrh56TH58Iv0MhhI20FnaaUq
pXPooEi1tj+taLkOmI00kmjyeWWLZ+sht36eP03DHxWjRxngTMPzzl8iQDtzeWVjDVJxWY3AP3xW
lnMN9glnPt69gaQVWQO117hzRgGWXWQTqUTwc3eQ2d6uIhweptzKWkiT/S9fZl0FHEOMpjElLWZI
0AHg40pB2UB97Q+qfQX/al3+Fq3Ue53jHVB7e1ZMayezjO0kTwuUdOQzCQXofyzyplbB2gXmj+Sp
7mCn/PtnD0SN2snE1CBU561DZQ9C22tNGWSx7BIR/dM4Sgo5N8H5t0Fxx7AjALzXzMWaYaZmAp5D
GCms1GEmmDnoWMGoHK2Q29btY3IlkyeRJD2WDq6z2NhViiBftyEA/Uyd82fc0rVsnf50tH6L4RLx
WIwOV9ilJ/CNvxHm73mYVjyoVi/8Q25NNZG0tng1wE5his63ccYs9a0IV1a24+9nQz7CqARJuhBl
c9LKb1GbOnPC/SlUSh4rduvH3nzKb0lMqib5QmFT3o6gwQAJe5t+zNs+8a9QGoasw7zB0CX7um/R
abwlWT/lbdKDEqPorNoZWaytysvus3SHW9bYK5RdYQybxYvFelwm9X87zQd4W84XHu636JdUV/Z2
W/2BKK0BoyhfoE0h/kwY2z2mI+qXANgdomFCrU1KOD4u7WO2tBeg74WKlQDtrBBs1wBY//uwVyn7
P9JN628fP7OvK8rSukZF4hJfvf2SVEKI4h5jG+OZLYY+UvASz1Xqy4LTqaOpVs22Sb/87d6K2IbK
G8wRc1/BDhmi9REvautzRLkWJ4e+Dt2VMkGSK8Fm9tEYvCAo8WGFUIuYG9DSDyKCQKrYkfa8QVpC
3ibEYCS4fI4YmMoeQf2pSu5C1uQn7TZwmIaYc1Rte7Zd5sYz6azL6Eeaab35TBC9QcADsOmy5sSH
/06TmltyRsGdxWbf17XztIy5+n+2wk72CP0paYhvEYQZRUiXzJQf4UWpal/wIguPxR12GlS5ZPG/
GYRbw0qin5MRIP8+iwSNqBH+Ta8MrbMakN3sADOjiFuh7rduT4qF6mzlb9ZfmoMPKEtGEvLkJN2S
VVi3Uwd3c9k8QZxXtLJfG+vtwjpxuIFcTEz7ZLds8R3F3qgYc1dkASPeAMhCeY/PRSzY6VZzGGtZ
gMeTUu7/fC8Nh9qekepmPa7UG3dPu4ja7Iw2Eg9itdNEFe9cKwwCkKD73kj+VBhqPvpDalHskW9g
CgAIDMD25RaSGPk32VsFMXcQReuFe94oJ8l9xD2iHNyK6emoUjpQX2JoAW8J3InZqobsWOYt+MfM
XS9E3OL8WQLbLMeZbUkrB6CxMJpgTJ6HdCSVFRTuuF+E/Qpa61qLkUTDhy1GLI72yglTHqnPixfE
bpg7IZsVQ9enZXSanI8068LtSc21cws2HDJvaCMQDB8VKutVzGLL6DtS/b3PKGNaEOlcxqgJl1Y/
0uuo06QrbEa8t4HHMHUpRstcxtXoFeKvGg4BOha1/kBOeQ4Nv8BHYtRdYOr+xz2FywJnoXPbqxrz
iGZJZji9iulRJXI5goloDmw7uTaU79vWwsAGy56WZPlIb3ZF/ebH0RXzWIDg+MhUSrezPeQ6ZpwR
6ytaoQB/gV9d+GBTbUpjPZp+yWoPQtDYsJluI6UiUTHu23yiSqZp/oW+4V0SlYBwLs1MQY5dxDGn
TyCK2lIugnrtESHKFWtIHBZ4ewWZOS809Ac/i7Q3ToGk8WtkE/L4ZOxQEe7LcWta9bwgjAVKQmIS
ij90XKbrVyDheyt2Akzdt6IuVl2CZzXCmaIU59pTTP8dHUIOBKWG1zUIWC45YNNApN/D0PXJXLzA
ghSIsRKydSg5wZa4TmmLHOIxxzD2DwYzhcKyyy9owSEXP3Go+e4MnPakxyKt1rADMX9WZNKJiUP6
UXy9gqtIP9DLP2FDHg+UKtYfOC1k6m8weuWSAfuNlp+4S776mDuoE8PEpTAE7Zq1CREGMaTvM7Ey
5qLpAfUHJ/hjCTlq8ImCaao6PGB7MEPs9mBkvm25KobAdagbm858tkCwMFqeDDL34D3+NWOcnxyg
gpH8P4NzKvrzWAb/6v5XeBwk9GEG60+I6dTMXqJX7IPIfOitnLWA+U4ROuRPv/kEN0HfBBi4S9Iq
s7FdC5ppj+KgbkqHywG7VEEI9sA8l/avddikGgGNe7/XYCixQv5LNRN8vZW8lEzl/jVJSAuDh5+L
2o+8YfUIgBwFnP6zdqeVjsHNeHAWZLsOejm2xJUF6KbLBrjmXPPvRBos5pIw0vp8li+SOdqMB5LU
O+MaA5SUqI3QUmRwfl7Af+3O13SQJSaMMZrysu2rE/wkpiruCF42z7mgABBXlOhaZ9AXudM331a+
XDRwFPIMOCSRDy1zYi2H+ond5wa7UYK3SCQsJ384hSRWlIyzMaK5UcgumWQLwU9mCpWGcnUQwdKv
z8NjEoXvh2Rt8PektXpRtrMrUWHymtbLAU0G+n6jYlXuVX+JfZjyEXWj3p9s9a5jaV1U7lomkLJT
HjDzOYdK7QmW7dIMOHXh1Gv9Wk8CoTFC00pN1Dw7wq7iBqfwMF06c+7vomjCAeERJTUQN+xXXkS3
LIiyi3cEjCMTT00QNewuHlVjXweqZWJkQssi1ux9gwbG2wZx1EStYQ89reGrGB5EWfHWJmLJGelE
NNaLQu72eGbtq5c77I8YC7k94+Zl4BNWp60hD9J7wooyZy7P3VkF0mlaVcNbsrCrCtWl4oun8tQk
2L+opPoawim7pfGnPQW+zkitxTKblqa4nztdKUzH4nIWPBo0IlFFhDKIBBfwR6xzmmtd4GdoxRPW
1xlVzrwSIHFyY6Akx6TvgdBNRsJ5dQgVoy0rfbjQQDFGPHKUZiqwIin/sBIpBi/VFETC657NBlX4
hyn7GjK3tYcgWeOy/oyYeatwwB5fM97FUuNSY9iDeMW3d7axx1ORt6Crk+tUlxhuIcqopj6X7C56
OwLvwPlv3vlewd94MaGg8xyoAg4+LSRC6HLi+SsVfsODneGkPhWnGXVtV+biNBMG3s2JTPEO0k7g
4B8mgsM/3FTiVgy45Pn1D9XYDJdXK0qpNRalMbiyF9VQl4g4oV5jEgc9GEoGc1N7ijEL4HqcZaRr
D2mNfXjHjj53pxehAaLrnHPZl5z5aRvHlCur05gUgm05XyzVEkurjSoB5n0mfRCi+3nuHU9XrQy3
BKFbcPL3gSB6vG54PTn0ptOoAUIXjN4VKwG2y53iIL8orKWBvlJ8IwE1OrapOMcn+momlMqHUHSj
HhnsHdjp2gGTDWBL6NgOu19WM390aHbG5A2FmIXXKeFcdcZJqA6AZu0/OWS3n1aWei+Lc7X+4TFl
BU5Pc7h9aAYJiBg9UYKPE242iwRNT2+Y5wvyXGHOXD0QuUE1Z4ScrS3yS+B1mndA+B65NkpsIcHV
1/oAc7CNIQO8380O5g8DG1nFO0Qnfy87EHLQmG8o2X7oWCOCa8580Zd6wlvEXD8xdQSOM8n0ZTHY
4rGt08Hmo1b5tfRYdgY7cS35vQNUP4iN64Jp4USDHQwkcupEah1diersjF1X9nE4YedtVNQ6bWbr
wZoJJ09ghS4kJLwnzkWx6swheTpmsh8GszvTpiEsc/PQdRi2sQ2gytd3SdnY3dvgyjwxwJROeFej
yIKG1SRdPvgrhnYGHl7zCe/YI5Pp9hXEEXmzXnSoT23HgWznjOWd1vJ43oetiYjKGgD1Kc3tP52a
wxXw9Vy18Oo7QFOQUd+ZesLTsnZVclybw9ZWMbXiIGsvdrWk/wATt8BuHqyOLVH9Ef10zu8TD8IM
CaemqVfV9D1R92G9z7hP57la3j6S07XnDHJEiYWl9diPmo0LM+GLJEpZdXqBIQLhm5J7CEt6GCCn
OTRfSeskb/puCKXCg0AZywGk6EbejW6BcJYI3cbEPiE4bMTqG+urSSIA7uXQNWPAKCBSZHYA/LxR
+Ia5n5yp7Stj6iaPPrP7IupkwhTOKAPIL5zvkTuOuC4ChGEKRAIOPH3t1unHNjmiHTT4uJX2YZGA
mfD0QMqK73+Cf7lyoyu42wxyGXjYjS0blMPsugIPCfO9K7VRhb/jV6t8CYzpfAAMUk/9jINOl2+t
D/lA+m+olWI3JurRoeQnC6VW6VQntDL7N6+MryHpqCfQ5UbWfT6vm5r8DAUm3lZmAmE7vlebbzkT
jqY3QxtVbcol5JXurROOy0dy2e71L70VkxtuWkvje8g/JbR1btpl95cC6HlHJjfjo1D0sC2BaVxV
CQqL8BEY7HOiqYqjsrK7efuxt6UtWxlvVEMDVYqQDozEF7ZppHY7y1lyOoO/y2VnVmXIOPQZyvRL
qll35ytDv75sMQ3e+JT5gEU48iEBM45jbWCxmr2hMLxiC7dPcajmmNdkv925wt1wOYtgOmL1yYNs
7BF7JMc/yTHocpgTNsKKurVot+XeIpbOeOukuOgNtVr1KpNh0QmTeJzZ+NA8a9FPv1EnAhnFaWdk
elBYoair3WFIgLpxGWjpRQLBXogmX6q/ghtdQ4Hx6YamiPDvfe5WeYGeVAfggWpK5nB2fdqsodbX
MawM1b6bmG6ASBWzynp8USf7wZi8l8bNalvX9VMXFX7UyMTepuc6K2Ua0osn3qXdGE+l6LSDT+ue
JDymEIEvE7LEcq5dnNCl1M5kwkN7rPuEVvhPPV5YoAP5YeCq+zGEvtaCxEu96kjTKyEy2/6Cp2Pr
bVZjWswTc0d4dgUO1R4mBSiRy7FP80SS4NIh/edmnkJ+68R13ToIGj1XJtcHu8fKkZCfe0Zoy+gn
RF2dHRce15k4vCLzxzNjPQ9anPESbIUjS7cctyqHdg9JKlQ1cPsAFGH8nGGO9zeOCW0VVn5C61tO
G/zwAB0sGFfbXfdy0mwHadbhsibq3FufF87I0Lnl1zRP7eGne6svbWfuvKjzvJI1u1GbJLSTHftn
hGcddJ+mYcB3yMVJaVhmzDhUlIMqfMQBDeC3SiP9XhYVeUzT7ldTCin6sx0hwJl6JhGCyrWdd5jA
zCVVkUBeNbYgijjKHojD4VZ34QJcmeyRVYIgDgzHLF/HFWE7rAK5nX/xT8wYDBerxaPYAsdrota2
YqIWRmY8BKdtPzvEDGt9dQyzeLC/euXBVg/r2xyRUOy8kIFtKXcOdzEmAnC6nVKOPSsRR1cC4WU3
Ni6gWHiUtvJAATLM0/mE8+syXC5dHUWrnA6bm5/6Gk0ttK9MknSoLAbdiZsDDjDbzac0gJG4PMCZ
+lXKsVJ7ur1WqzeDDmktfKsHsU+uXNmUhgerIAzEUbPDrObC95rGr1L3qnpdecxQXMGdxAqMWwkH
vQ56MlWPqVvV2Tm/bfLdFhwkbX+Qbh6859Y5oozCaFUFlT5RupqDmohGnvmLWI3IhBxsIIGGx+Sz
N0zi2jjZztvLf2Y73pY4egTmYuDTU+gr1rdbVLKeU3KRPpnj5XUC+sWdaXdowpCpP8YHbGIJbIGq
5v1OlUxVoxP8RJbOFHa9fpdEaFrZAp2gRWdSGprqw1qrkUU43vnBuPZwT8rQhNNTJxqZK4dPuhaf
MWhpLICd7x6b454ucHiYdKNDXyOBaNddESGjAx8yaf/Kj5L8QOHfSz/T2SulffUaFsCxsRU1r3hP
wefuZzzI9xX74f9mb83V28LtRe43FVlCsUcRqA/jMMgzr52kT2q5jeIjmsdd58M1G3STIFAZfDTX
39Q8cwwKQAs/UEEdmPtwXaom6UX5YNnYV03kuuFuUqaJYDOJksCzaZ905xjs7lhntPoMnF2jRqLT
wQ+gDlGH4Cro9ghF3c9iIlKy+y8qHMx/GsmtVuvo5UKcNBcRlEuOV2sxnUuzqZWD1PBruoOD6ip9
WiXskj8fxd9QC6q8AaEiQ9h+nh7oSUQLASewUr4fZfvQtFTngVBZ+7DEM2U/RcS7jbYHKjjGc0IJ
Cd0pyvFPdqRb0EcoSZQQzrC9cE5aueBOHQf7uVDCopSVOHBqeZvCSQDs9h7V+8BSjMNjqai9Aq0v
lRzAL/f3gpLJpgsIWdSccWiOcPKi2CvH+rCUr/vmEtgUC94q5zZg8NRwv5uLu34oA3VE7RvF9yJo
iREslNIF8Z6j7SVwTQ5i9K5TYrXrQuTIdmayMfmmH+LjvUoEdENJ/7oeCaPVP0WPirOOEweGSCef
MvJ2nGPJpHNvxwOL6UmkNvM9tVhRySg+vbcx9j/Np4nzn8PnJpRnaNYHT975i/2j7l/VyNqDkvvJ
l93yjDN21XuLxIOm3LhZ0BFdhFndUN/F2+FOXPYnZfhRT3dOrtQRfDEiKNAXMzZTTuodAtnFCcEi
THvhsnkOhlTENfCXkLb5hOn61xfMcHCyueK8jzCJAmTt6WjRRpgHea02NO61AhJNU41k6isCP+Fg
fB06F1I7g6IiCXCRIePaOtAiuY/+9LeA6qCgUY3fkVDztH6NyBauJUjiWGauP4er+oBRnOLc9Eu4
eRqa+r4ibF3nh5eRy+sPshysYQuHkO4L+/qwsTg7QNeWorRVUWx0idsEBqWNW6AMUfIDTVppdH4n
wZcSsVjJOaAPsp10vGiTzSPjHct1CzX/0vp2Lr6/HdxHXwSYAaCKAhFfRN8zgs9Q8PweJjLDCBLu
u5roCD1pzkd4Q+aNXLQou/QBq0BACobeiWngWJEFhHPGxsxFucspXLXDFHikEZdPCpyQmGuv2YFM
5O5GjfAPVW9RFnMe7Wxd6Y3UYjd6ta58bvgL94jsCdgTCiK4BoErP45I31NA2NgSS/uWRv6w41/9
jChWSXVIf8tGT9KBnGa0zNvGduqO54ykhT4Gr4M2MJpZ5/NvAiafR2wAwXwj4t1ViifHqFAYMq/I
+SFxs9Wodb/llTIUZvg3HI4jHhhAvXZIXqzL64jRLZhpuZZdRwqVmmdewOfgqEcXi3ynRYcpfoP/
+a+sqU4xuMbBK9knlMtnimDrKSf23rTVZq9AdPRT4HRFdEx5+v7LNSsEm9sfIviBdISl38uEjL0V
Y7/AxU0SLzV7qzB1L6fTyrE76Xkl8bF2alVVNdzXVv9HApohHL5WQcaB21co1Il95ssodIvRh4Fd
IrwW6cDpXzgsV2dopBZv3Q+Xcnqs0ubSxqaTVEbfZFLtvEvTJyEvYH5aKQL+Hu9eRR3lUzcjQQ/s
udBRbT+rQs/4MNQIwhf/LIHzQKXbRRUEwr456wcoCTOjPoJuCFnrQs+nBX8EaR37ZMdy7x9U4dCN
f9Xi1BdyRFVv6VkhgTmIN11cPGN5mkbEhzKUs+o/7iFLS0iwCH0vTao/8ttk7O1BB7pm8Z2h7eMT
4mA5RYE8tBnD3LZN/4NO+KiXKqfcph+89cwrR+hU8mUD4GOPUfxDTxWAfXxPm5I192GnJzwaiu7U
sTPlFJCVtRnCr08vQc1Yr5osTChMXFJ9+a16vWvryhCPNJ0sOBo2fjjJloTmXqNk0ncr6Jng+7wh
q2cS6LLB5GkfU05EARwGSQ1mIxRl5Y8LNbwXmpvfbWoodZc5Xq2bqzRsEjKd16XQAdNI2cSbkWjD
22pcCx8eNHDyn9csSGuyREzuryS1gpf4TBrTxEX8iGF/ZWaYOk6QDcm7RbbYt2O3ss/skr83cH7q
D5klN0SqiwlSB6YoXc113wgeTqS9UHnb0lodjEvvWII67p+N3hOWQzSuN/U4R6ZRaRRqiUiMk7p4
9Qf9Hj7+hGWuKQevwhciYIvcEX9MiQCDYX6t+EGIB9AOcB13TrlLMEtlmiFqAuiOoxwrvG3WuwAv
zYAOnP05+YamFlASIG1Mlf4lXO9wqBLmdmOE0ZtJZqykS9ajO4H9NVr6oqGz8RE7EeJLUzT9ANgT
OiES59BvMj/v5BIJwr9ePkXy59LST0L9g/FOqohPQ9B7fGKCsuWHpgqYiE6NRTMrehZYFu+Dsgnx
93M3LjWNeen1rLcyiWBwueIzj6wToV09Mssl5DcokCowFk64RwuJAIfRu8n6AfkZ1QGrszwmD72b
d3bAa377My30p26KP7uKv+29cB9Ds/06nwWXk14mF2y7AHuCV/gbk/KvDBNHMh/xQ59kJOYJd1yC
mZW1w3FjZiwALwFpJ/rOV6emKp983HB8FUDrwMsUJly+bR+pcGtb0Y1mm12IRs3Zw6VnFmRu0AJE
wFhPbSqbSegv57z9AdnyGzvqvHf7SBVWLIMCRqVgTakNSMIHz58jUxgwGG6+v8UiQAv5TAE69w+2
Wm+3AGvlKw55vNggiOjBP2AYGSw/0RkqTFL7Ubk7ETFMn1Qe9mvy8yJrVeCRhu7sZbYbzKtdUni1
QVe8eviLX63xcWUixcArnpXURrK3qpJonw1lLmuDL2PrLIBUtOsT+sob3tEBqjVmaOmw7IC593WY
L4txqz8naDgn3vrfgJxQlZZzM8V19rAZa/1oiin2LtIRxUiEaM5jVnnLaTj7tZ23ozcwvZlbRssp
EU3Q5AhlzFMx/HENE3vIVYNscsbsFmnCr0DLtI8D8AM22jRTzVb3iW1N0tqxQITXSKmaNDydZSbs
t4z0UqMjlYoNfGj9ketsLFZoqN1yJ8DtBhlyy72UTbIMPQblg9DJQqTuqWrENE217t03f/HX8qUD
1wB/5YvdyJVUe1sJy3kJakbFmEZ0uStK6InSmkGwHrOFjZLUCK4V5th1HQGqusBMCQV38cCZK5Bq
PQtarw7+4tMiGSmvYF4wCoVP1uB4PgbLzYcZ1vz0wbS72qfHjRLYRrMw3DNqkglaGHsKUZqjKORD
cKinfe8tH6WS32UxBH1DtDL3lVSLjHRWh3GQlY2UgGrshBdeivuLfl2j3bVfLaXOfoHsJX28EwxJ
GAJJ3ePozQzj06H+SnyDcsquRTk2xdAEPql3jJTGfXIa5Y4rxCKirgY2n7wB6NGUdW1U9HShQr1F
tgL1/YANV8pnkS99chFC0UtUqMT5EKKB1dsvbKSEkcZLwz5Z6LXNEYAd/3ubmWAboDvPN6siQKu/
9Aq9bwehxOJTFc9o8m+BMmvzJu1jSx7skf3941VufQnqJzSP8dbxAzQmt3l1zNd1x7GX6bXetlF4
eRaesRLSG3ZzdicvNH0yFM+VBpsnj/phXjdm9Rom5uSQVBh03A8jUBrz0Xr+W2HcOQ4kkVEHJXYM
tajabZ7azXWEhcbdQV5xCSbFvjO/zMamU7QMD2OS5/jm8B9zyWu5UKGzwtwFJlTc6oyJDQ8knUDc
fkOqsZ+dA5rl8Nr8jzY5c56WCTbWSO4V8ru3s6XoxEYKtCetbQ5it4poveMkE+iIVCTcRY4lf35G
L2QJb029Ul40lliSUj1Efm3VYKr7A+u3jVkydxIL2kSSVJU8Nx4e85qGg/0IANw5LDHC+9/4KekT
5rcFjYWCCHrEau+2G6ddEduxkSI2SOUzFKBctulX9K1Ipr6hYGijSzwemFi32agSqkN8d3yLu+Ac
5VEEVepII5zFUsYtG929Njy0RQo0tvgssLUPaZSB9FvAy4M4EBNHdmSnkHaZREdgBKULOyoYfzAm
4OQZw+m4sK4SmLzksEnUHpN9aZIwOOipTIPBdSeG3hc9PLKlpNpF/hlW4/Sxxt5zv2AWb3TMzbxQ
HHBX9gGFInSWFaU2y3Qje+IrYip7VWhIYJc/wf4vt7bOJbhVvPIeYo2xfbB+qu7Y20hxmNg2y1t1
AwjDcgtXjd/J3bXu8PNzjKjMSj620ssqaZhmWvxoZputZPuMQTRWxK2yBcvaGA/v+1YTdTnZnAu2
Jw9oVuFA21S2mHSp5hGR+VMh8vREIYni8EWFPYwyjTdmGW+woEcOg4mGfFbyyiJ0X3fBe7pWWxKg
qgwdDJN5VkB+GapNXONlFxGvF7sdL5mRkYTGfX9+giqxPGVJmL7MIkqCh+CVtyn2pWjNq4GAiPAh
IHoJUM4jnGfmlfJ74Dzq2YtS5twS+GCdMdnn4Gq71jdphe3uf+jvblZ7l34yGQ32ru80wX1jGgoE
BFE9LEFQMjaM2RpQFYkiLQFdXqaFWArRWQVxIswCJE1KpLo5N5Iq6J/T2F9NZ9oZLGnIMNDRaNhe
PWhBmHPsPPdZy4ToJreLapYI/h9rQcPwrYjXrraLj0tyPzHYuuCGxKjTjV4TR6Q6clhv1q4jaImC
iTW1i31Y34LHZ7EQ4Ibr8wozXihjqICPjFebAUuzTcVsPMg4Lo2oAvy50Ch3fGISxqqXGRnBdWvX
EOVIl9TCjV6/3ah/Exj9x1COwX7YVXD+ghmS5l0xUhsSD9Ftz2SAEQEb4LuEd679sbzbR2r6tTjb
vcvRC8qEBbnvLC/n1uNlqWGZqgu0pibPTo8a2QLDd2cmU9xqOSkkoDN/uDl68R7Nqh6qyX2ajWYa
4nSaWTJoUnYrT8LdUTF/O8TlS1qO4X4uEbm/XwuOnggYgz+jAvgOvNth9hvopkFaYtPFrK75WW8l
R5dCX3uSGEkn7IyA8m2syx1u1YVhWN0AB1UG6GHcKQNHNLjVromhGjVXfVA1HvFUQJO6TbcRbRwF
OVwMJSkPQAN6X7gBKrljCk9hv8HKlgms5GBE2hT3A4k46yOHzXjdIH0AtrvPJ4i5gSnhJjn3GSgs
Lhv0JelLZFaErH7qeyDf3UPleH/J0dvqw4pTm0oXw+2JiOtFyBwHb0QnzelnLyI3m5q70tqvgIEj
6TwE4k6iXXo7OtfwU10INIWXKk7CFwBmvEh5Impl3TrZsS8HufDf/qFjMR8mHj996IOeYtdpoImb
mGV4kdINf0ralxNYSZln1g1Cmoy/SJ/tHMB7aQo78VNmNM3rEgCZMVfz5zRHNs02e7Dl89aZTJgh
/vKTxOAZRaOXd12r6uflp6g02U7/Zng6uy0RJhUmWUA5uzEt8trsioeYvIZdQtGuNXpkBoZXw5sn
XLzmOqe/Ia99474cMZS3sC/p7mRHwh9TVonTx67Gy62hHtm7eBYctcY7yJX3Nfmrey1d66OOlLUl
l4ElH64849qSDYN4jFUtdmSq9lTmQIck7mYITV78kj0ncwV8fJe8Es3OzB0pepL4uodNl+Y28hh9
2dRE4a7fODXy9EneHXaGoO1D+hREAWKQIaHgesdw+SQ98JrsVS4t9dg0IVMauTMOFNYiVEMnF1lF
F9NjJy/RFFGK2JO2LHTnig6bWCTXwGThWwiU02pq+25fo6YSZPN4PgCqTqBbmUBIfXVz5yq5a2WA
GZoBspRRTA8vzI4nfyKZjN2geG1YUG079wiZuSBPAEy5GiWACRy0en7lPXOOZ4wi8z1h4DpVVtEA
cH9jTXivq41qJEnR5Rcnydu1AUlTc9SqOY30AWMNm9iw2fahanPInEZcqxVXiU07hcHSBxukAE4x
IGaGMHpt554gjUPTVLBTd6IHp7FpQDg+7DGs0/cBu2+u0LKpplSFI4zdN/tZB1iAATNt+LsIz2zw
lFMT99nnbzegiKnrP2FcNuw8EBglN8iMqsKSZuqL4XiUE4v1ae8g/tInLaljWhjvqj0Hyg8Sozpn
IRtJnTyrnMb2LDCCmCIIWZrdcrchTmOD9TN++Y2jPLfOVZDQYPf7Fcc3qGdoHgEPHsdK3rAlMA/E
o5ibKFuoLEj0tkWdDz2NlxgV0GZDjp28zszDRbdYVs7umpRPfOkvfhN4uT1HyczZ6+cz7XWVfO+b
WnOCFYae3s/x0gQZfXrLy73SiVt4GR0PkNebbgNcQLkY0ivWRiCvOPd2RJmagMQuHIohoJazXlfD
piAYrO3U/ZWYUlGEqvU/2S3Xpf4qzuBy2ImVHsThhrXMWUF4uVH6+yI0quwABJP8fpxRE2yZmFTi
RxWFEejbHM5V8dSqV+kQZ2C4WmLZRfTqijxp+DY/t2YtsKlRU48ZgdVtPqu0Y1bi2AM4jaEDoeKS
LrPaq+dmjZPLIWoYmXHE3mvRBCei4L6FCPiVT2SwhkTP3rtlmBAmdI4hK/Fc/1wKXKBB7NR7wQfH
PTI2vMDMsk9X9gh/uEvSDz0/5jb7CM/5TvLQ74UUmHIih/Nt5zJeopsTuZmMljM2xCEBe0lWZVD/
iZhXFw05i4N2A9dkAwXNvTwU6UbLca5Mrb1O4SHgOUOZCaaHb8azs/FA3iE2+3FDp2LdvfiSwY6T
sxyoUNVuTr/n9xZZQbDnTiXEqs+d5bUg7AMVp/cTSXboytgaATXAeWL+PDAqiQq1rdM1UdOa3OlB
lzn7F+7/Qs38F3TkHYkraCahg/oaNpiyOCe1I52YO2XkpsAVBFlheTOGuLe/KjAPnwCo8UezJrDu
fsuEQXFLoKYum8imsu4AhHiisE8MCOia0VWYfYLztLjN8fkZIYBuxZguxfynvBBWfPQ9BRV6dITV
JCavDOch5jOcQCkRkPk5ll7bnMbD9u8GPyxAQwlhA3VgWWYo0nFJFX4q4UvHMcxatbVrJY6GHoMP
KyuDTu6glIW0DUu/R3UIamITNvJOsgju+hOUNWJRJgwAyk+ggOEjhIqEfkPTZWAcQU7M+czJ4oqS
56PneXMOoBba7v9D4yPiU8rpkhshOAeR7BF7arcY6G4j0X7AKNVyiqFPHrTgFJWxZUDXFNURp42T
SUEKP9LzDCkHFGoidoHCW0ZQT7gU3gqIi2HRS+GxNtIyH8d6UxyDLvJvbpiHNU5qgCNYDltzVXm5
iBWtkV5uJkkWHwuPHr6AtVchon0TSgch99YRzliKirj9pKgTcm9R9HgOKmpepqADR5uujuao05e1
dbol7raT/BNGgL3Ex6975/8dx/QgwvrzJtm1a9D1+gnIJ10+bXzcqomo4rLEPSMX6vR8dRg2du4i
Pt4x86CYU7RupiWhUclGcMCmHqemqUO7UcC/4nJ5QT5mH7lFXHXqEwAxL2xK3TubRow3GwfNK/Rf
DQn8oXKZNs8ckTU/FZ7qHDTXTPW4Xemz9poJK1fGppOIbfgNhePEk34Aye/wWh9M8fD+lC5nCvO3
IKEqKfPaUqbDO6cxnvuTazpORyrva5bdKRzf6rU67P5JUdNtnMVYCoeEe5e1HkKxcaRGk5nY0+JA
WMw8JS9+4jby2egwAfJJRzP94TGpAdpb4nkGD51wlqtAL0ffNJ0LRqBjexCDgGQ9fgmK5Z3+Gpww
b9z+2ajGPuw2FThjAAV/aAmfbPB0VqtZR99swfPydV7zsqonRsh1XmWKmCGM5vsjyBfo03hh1W3j
AeJPmMM9slGFZFR9ObUbUbXWxiUtpJQ7vYGcvh/sTNoS+FXrbJdYjBouuHHOIugVJd5zLWx7bJUV
AoiQ9a46KS5omaRW01yu6bS/Gh7VAQK2w2hGKIKofkRJ3DFTXy5kGJM2LxcQa0wtJfgs4FPkb44R
NJ1Innmd6cBxtJ40Dns6nMA3RnGjzsuZjYDKWdgMSDNtuN2ZNPhQ377gLWOwWuM9raB8Jh5F1hH1
YzLy2W5kBFiQRORNOLfYZlDGMgWuTnll5RnUw5IGQqVJroPE6rQ7DZXo+O7yMEOdoL6fGeuiXux6
aho88eLjbkf3aqS7NHQCyakpX1omkpncrAkNKaw/mFxMuSce6ZlDAWAUNxKvyHY/3yhCzMSITY4O
ibnQioqS5EuRnqYcqAKw1+Mwgtdf3Gkkfqvi/Gnw1EbVQ8PcdaNJW8tNjf8ugaWiwt7Bf5XN63qK
+uFGXlJ7t+CZAC/YjGcv0IzNO9IYdR2x82q1xJRnAayd6OSeWS0pwfgyQM9k97EwZBL3Qu0YUh67
pln1UU6lsS5J/jfREuwHoiF7LCvUFha+YOpdAeFsi78GZCsszSpJSDPVq9qpRZcxDupIt6ERoOdS
8fWuZhVR6AuUdgP6qQfh3gHy69dbniJOizsSamjc0e1wqc4r7CBUec8h7mH+ogwyVWIgzc3K7hfK
rCttaP6QaO8pZrY7r3YfOcwabZjqPWxsMhGKHcNvtvcYeFcvCmtM8MOGgRjhYvKJ8any5xdWcJ82
CAag3YYRxAI5cgvOSKk/kuALNm2UW+TxlpaZ3yqu+2vfmnSsfq9Pc5Lo98GzlEN3RMd8i5AqcPeO
e9M/FO5eX3v4TyOcq63yjKxAe+F3aCYUXHaj50TqT3znEJOBmkM5sy6symcnvO4YQtWkveq4Zefv
Kz98WsfCirgedqgbqaSXK3d2JGeW1BNuWryidQ5YTWPlqgAPapuBVVnsDI/UtBquohYjES28Zmy7
lswNcGJn+Qgog4E01sovevbzjiFKj566HBGIgfiBKJAkFiOHXXhjO5FLXQeu+9EyZ72RO35oQKNH
snM2TbOL1BjNJlE2qZg/174o+as084dpX2PBKzmoxclOyxxdYIp/edZDwCSGETknYOxad4o8Yu6z
/CgxDwSUQykcAlnv536sq7enBEyfCUJrw6YOlMUJTmSqUqPJszZ4/A4zBSMC3rpi+0gMyj6Xm1BS
tCvg/B+uovgYCE+87gyFvepAls7bHyX4WED/F7AXd5BWhm6dP3XJFQoh8g7zguQpDxtwtkbvb8fM
aqrusKXxFJmnJxG9BXcN0MbEd+n3paaFiumAREK0RyWDFGtyBhK3Oc1MfN0nyQ1F/KhzScnQLm2s
TrVAXTO9EJxhiZzMb0ONS2l7a/X7oWQTC/vk+0eyEhoMwLPGS3S9RBasLZTmQblM4nXcJ0kSQS8O
8lEjk3LgKWNdQWdOIT0nRTY/FHscvHUuAJthh4Azv4wfvc1D9ny6VPZ9MTuj77hq7+cBZUOxeIhd
uELE7IFhJv2+lwSwTQSqkPo+Dli0ezrSNfwzvLXO2l97moypBFE9uwrTHmUwhaaNp+oeF0aDXl77
jkqcOqyuikjVQ97w6BvsKJyAAQkilH6SYwlZ6quwVfE/NFRnZXlxYsHZmPoVSA4TyMA3z6Qnoead
ineQ+KVxNyBxIgJpxqarOWbro0aXin86kmxUuH74oEAgsHxb7Iq6YjGsWcsBKihvnQtt2k3xmAt9
HA039JLnSQ/hNPMlE4livHyZQlDvhY8rH8cYDmxhmiZQNPMbbnDEi5MTtAUPW1gF17hMc4L3b/wk
8QdRcsP+V9JEWky7PZAjcMdOc6iCn7lXXqr/M8jn92t/cSzVAmunorFez0OT/GcMsU91vDUf5shp
FsHrFcxnIudRemCXwisHLc0tzLOHH2J1V+LzMcDHVTW8B8cZ9p1/xYMZWjStLgon/CyequhHT8wu
Ew9Wf4DsvBUEskTTF8ySIcpfhDq8bTzThmRYyVCLTfU+CxIVOCFWB2pBhRas9Li7eOQpoFppXCig
M8A3QZIxM4ygLxKfMj6fYRBd/5rfVz/v1cC9fYpnzLWU0uB56quDHsYwsWyToJtvORDBNfSwrZ7f
X7uEEEZVOj9tHRSP1DqDHBwxM+d+H7Knx0xk3P0va2CICAzrsscmfX4G2KB1aqKIcusvlySMzOZj
SqGDj5wGsUH7xGGLOWbTRzi9cd9bM3a5rXCwfd+ilENv3PurVb8qTDHsIhy4GdkBNzUqlteArKGE
fTrmWhCTN/TmtUNkBVQ2ER+qMnkQUNsywYo5e5zQ6Vp/G+o4SjGlRjnUKeDi5ll21/zORKBzjhyU
SWV04UEvNfcQT12MCjiEZEQqLvgeCEaBK9B/Mebj0GoQS601Y7F9wK9Jmy28SNZxWAHiSN97e0Xk
tev2f31l3d6m6/wMNkggu+kTLyikFTJq6luKHnx1PF8PlgQmqwPEaQAbvXtuvHdRo9+tsRFJgM9P
CCYoTfJ2mz58kkrXSHlpjfg8E9aSlpGo9f9zy1j8wZBjheBh16QGLs0v8IGBpxFNI8jcu72q7JR1
MjV5qOewXWyBHgZzd+IOj2BaZ81gLsZc3w8tTqZglLM7/XpvLfBlZG0WkcrmZhLgbT2aNaXvkACR
JR6UEOBSYBqsQt81IwvVwiOHYc443Gl3v2CKum5Q6v4GeUPiKLLB4hTrvRI1oppBDw3OGX6quve8
EKJV/pxUpNGNU0sJ2gkf7kcqX9K1SkEtZNCD90O71SyBeGJV+5Bw1Ax1qCVums9SzEUxIF1ITByX
YKE2uuxHSEJNbeEN7Jf2fBAV+RJziAyNBUvZh8wRvPlvm9GnMX0vUGKEWjpeJE3DAbSnJrVGxEtd
uBQDFn3aJU1dsYJoomZK3rjq6f8jjRrJRO2PiIi+jjwuMyYYtWspe/LivbFl2W21KbLELdVwHtJK
OXb7TeVD9gr7a2NGasLldeLT9maxxZm4mbalW4js2NOkXwlllh4W7AblGMZB5RrVVpVkMKUBCOkP
cEmNbidxYv2Yt0aVcbvg+krrftc7Mt07BXmglfm+ELYJdor56FCXZ41+PHIAHf6+aHejE23QzsT+
bUC8ZVDrhLn2CxcOCnyLEDm7b0w4Xd6bz6tLcCyZLht5hxct5uqHrblQgSYM6nY7oTMIxN6aUyvP
gzGcNhKXm6nQ5jq4JQ7JExXEWE4/ka8qZWNCKtrVQNNZqiwPF78Efw3lAuv55mtyyoFxIjt2MfQP
P3gM2AAO6ZGsUoJn6LxFnR4Rlf5nn9KkqgaVj0Lill90YVFx/l7u48t4zx6Ahiaxo5SdsukqhND9
fCcrG8YwCB9EmIorZu87DSoQY0hm7+QcUQeVKFtJkUcZLvCWsMhATcSjXL4WBTNnYVJ3jLF592Wq
t2jkse0uA93audMQKYOgaDs9LyKWasx+ggFN7OUudCU+eMJTmx+YKPKzrE+DYghOcMBnFJK2WK2k
uNzQHwtLR21yk9+VCp+rDIyztnKmeIPvZ1LSFW18f/P4qFSjTNMhDvyrQ3GsQpNuK20bowOwoZPv
YlQGqO1jxbTZHgqYd44l2w4HiTWdGNfQqNcFuojSk3WQhMsGQheU3DfqyJA8psOnyIdln9gnvUsC
fsZEAnUY/x9ptk8HPv9iFf4JpsF+ao23iREwG2zoSpAiLB3Iq/LFRP114JwXEF4hw5/SWb/Mem1L
sAnNd8fBHWfmKCDPrOVfxzipbuJF592Mi4BIvE28q2KQglZLqzHgoZZcHORc1jsJ1K01fV1h6wKQ
TZ7GLZ+/7GabJpaQSs53dC+yUw8hyaPUpUTUfN9xbi5PsBiWmcRAbM9F4Na3bJJFk7BkBmfafstQ
vCuxXJCVR7C/khehYhm+DHzfKd1g73hhnj/SxnZF2Gkj6tA1hKPkT3+CGpjHZ35Yvl8rKQUG+yH8
56QBnUdS7MS982MqteSuZmYTgmNrP+AD1exuvHlzWm40yGQLWxvQsnDeuF69iYLnKADeoT6jMLry
7mRdNNA/gSLD3+makg0GfZBuqPjjUHDyPiVqyOBAPx18iCM0EhKAWK91gqrRTrd0iSD1y0QIR4f+
PXuKtJ3TI0Xm7HMRFp1MiVTTIa9HXmcZi0tGSE/C++EY7vDBBTrfC9qT7FujwroM2uEBDhO5MJaW
y8gbHMYGICLPnWEditUnbR0FGLjeRSGfA/oUL0vFMlhybdb8fsWX9xY3+4SfRatGEQl8ugue3AQP
7bAl0ItpkxFcLTNkJn4B7CkTAwqQS9ixQUsg/1OdBtxKvsHjSMR+XMFVsEfIyTFklYKiwVyfVowN
j1pNY4rHhY8dOsuzyhWEp7rKDTk7r2mHoFBHDwJ5Obdai6fCSEBoUl5t7LVIuSI+k9jDEdSFuzK3
CFllSsytvroCy5w1HQJz7rmcdEZKVUAsAsvw5bSJctzhjwYy272XpUaGQVbwkbaEtjGAzYIom70T
dOx2oM1cwveEgASNtqGq9xP7SvcxsMJWOutdK7R8gExnoyUSiyHQzA9A1zEKcz7qKBRXvzgp0Mlz
5FmrQKztJcufueEyfK7RSBdFmMptEM1vg0Z3xui9ZWSZnV2XI8RaY4Y7/7mSEsdNcrIM3sCpHOfJ
u0B9WsmUa9KrqhzR+K4p5TGtsDLrKTa24leiCbr7UDevaDbaFs5fM0/Vob7BjItyFcrPhC3LIaSZ
FYvNtukNcUTjwpcLKDHTnYRFpxYM/taGn+2yWoPPtsMsOXuOnT4J9ZxS+ZV5i2C1/tbOosgQMxiB
pPiqn9zmYs8851v2GNc9liGu9rB132dwGz2FZaQz7cd+ozqfmnqhkRSVffj+gozJUjMav4d+nNWb
6DpTJDwNpu8oxfJOrImCvqdOEyxUa6x0GZPDTnn65vthro67LP8P2pjLn9x2YJJXLcXr6PSbnOuk
iTIWdseLih3Lzz7khVkvnjGPRIhoQRFplqqHE29tXEqlXfHTQ43jv8C313K4EXANMlzg+N4N/C9W
aCLSkTvPiRLj9B1g14WPUEQsYZMTjsmzER3sG9wwTua7WlSt0RrtXsnkQj2wIgPiYIx3KVBKE5FJ
3O7OuZltAtvfSabP6Yhwcwiu8K1hfpThLyLbU1uwTHtMQGabC5b2hmkAG++J+wD30+WDj61NaE+Y
OEi83T49KkGpu6QuD+BaDAJhG1+6k5/OVKTrkKejQw/8x8vyrn2ndtI4OPNKC6cLbfZbEK7HzSIQ
BKJ02UQZGZYHtfV2aDtuQbBtle0bEJc4rojS1KVNjksws9x1U5Dq5xp8vaBADZx3JN/rFfxWfhXQ
bX9vcZ6jM9z3qUb4K/WZs/YCheOOjb5eVm6CWq08p8J2YBLtMZNENmm8KyXVT4Ih3IyFoyMfWLLp
XPoirNwmeZUbIRBqc3E9BJXUM5ysioZXbCSlJ9fwpIn1JTl9dJsMEMkwLaY+vAqwrWrUFqZOVj6t
Hr7/9w/Pdx1G+6aNtFxedStUP32Hry9sZ6g9uei6PiOsV6RG8uBEHd1ayq+LQYOmd0AeDHM+QcFM
D6uYLQof0M2tDtqIOn3HsEyGzUspzmeSzIOMOTOu9R4F386A+WnzQgmVzkXS5EfsVSjorpLMTgcK
qJFGWi233QNjsX3HbA4JhuZiLAH8CUYPRsncxJj2Jr+kh5ZB+GX2//t/W/mel/6AVWXKNIntk2uB
AMu5gVAOfZrCIfEg76gTIDsZHU3kAlpjPop7AYAgrOSWdtvejvR9fV/1tCeLRCkrmpN9c+AIjv9b
ociIKhCiAL6OqCThd5acjMK7JYQSUoicHhFvvBindpesDx6hxrDkkvpFY2gfU+epH1DQxXh6f/sf
sCVim16IWe8qiDnjnrOiaLE6wbd6sOsiyHy5w+7ymbvnpMwxxvgo7/3YFG6S+F+CmMN0ddQ3j0V+
18HJv1pQUPvU4CyhNZCkxI91wDYtLJqDA8J93uj7tmTgD66GTCbkGGRy3kC8Id/JKmKLW5aVk6Xi
bZuJoVfLgR+o5GqIcddovD6QVzsuSAt4/sakKxo7Tup5DZR7otyO2vPrYgBYujfkXKFe8H0k4dkE
mSn4dIJkA9lQb/ZXHiovR4COWRvE6Paaz6ZAQ1fR8hnRbhp6dOU96+7meXNpCMXkXyD7KWO0Wvyi
zVKJvBkg7g/jbJcmhwFZvzmkLCtHbjBsGzpBWHDlJ/W8akGJLwzIMwlXfSdPlgU0f1yIfybcgihC
HGuS80S4jjga9T32wJqKu5tutJDp7JTMVIe2sRIJHDv2NSnPcSsaEsVNcnR6S2RitYODEI0hgxrQ
2lIMwZO0TR8Cf5wRc5ivxwudFiUUIz/N8mzRat+QvwLRq2OcAx9JDmEWXNNPETqNhxVJ3sqwlYcx
7T10zkvMt9ul9bFjDvstB3m7tGbQXm+pdueqjLPL849wSARjepXIkkUSkQSo8M76i7kfitz2DaHv
wCNk45Rf72GhJyop1XLiGHdk0D0AU8Mc9dEXDdUKnJU28Ba+YjBmlnG2dSTb2FY+8b5RV+t27BI4
WSsVOWwV0G003wz0i6ZVcUICTjf/JVBranejktplMn+MYBVftgrR9QCJw8qArkjoOszO43iA0h3L
LK6IqYQgDUgbtegpfOwR/YyFysy7GtGKPXw4uZR3mivzTLFphS+3+muu/a1FreWLYM9dBZl+/jjm
/lA+DR5lqQRvqiaBFEYBOAYxQ45hGpDD36c6pQQcXIMPl0KHATV0hJhGrwuFXylSwI/iNwFDlm3p
nLr5sT0BPBF3JkYowsqCNBfNvb8EdmaaV6F793F3QHB2YNMdgdhOd/kEBuM5ocq6XkjHrziI6jez
BmMKSJjpnZKiqEWG3tjNXPPLuemvsU2pml2aM6bdni344Ot7st7kPv6av+hZIQyUcyQ4SCCAIBFA
uDVZnTnrQXsRS85aRDt2U+YMgvWaopFgNuonkyUHpeJsUYVGw34SIHtseB3vLqTrPwzTFR9cfJqC
XdTwFG+GQz2xUAC7F3qEth3jTzKOA43PGlb8o7ftYNCQqe6Q/NIJ+ceDmODWaxA40ULhVUeHE7Mz
NTzKAARY+6IytsNmmX8RruypqEH9zgVbEl4iRGUU98qZZIcLkQw25sq/gpKZ6HIN+plfGpn0iwl2
l+7++m6347bbagtH9f4uXKj92Z3JGQ840SUsnT6zzZLNp7IQF76SyLhkMNTEeE9FqCCRJe5WRSxk
wpuBESOy2/RnOv/SQX48E3KIgv9hyLPtWNJuvNEOecZnLCB61kGr1AJGe3UQeEQZidm77S9JisHB
So/uT5nm9hxhET9KkwnItVyvjLlK/k/31ltM5sOT8uvr0JLYZA9+IDfcSrTcJVMtThjCOwEewfy4
eBJUSKfhU5UKBBj5nTYrVrpiHM7uaRruEFiXxrGngKxj0HS+GJZ+Wsqdzu0tB/A5/jQGWA3QQ40F
eXX81rNBPGbyCjj85Pewp4Do/0zB7GLQ+Ojp7pAl3YQYzTIBdVlNUmo3MYb1I8+7OvSvbsxZOdF6
U2e10xNEIB+qPAXB1caJ3KgPeRYGS82rJT/8OJux13h1X81Dn9v0nZZvmZoXJ+1Wchas62hnw2Av
5eRCvSka7gQdd/Vu3rZN8x7DJ0DAdjXhZ6RJozZUOZl+50xnM55dQImK/fF8rjJPj0hWT6vgQmal
qALsXa1VmQsKtV6Q1xhs1Dz4nxeyzES1XwcrwWI4y6CKIjdione7OJMIFy2wP5andyOPd1eGuO+F
IcJX7+w4yckTE+PPb5WOPlSs7fisSwweELaAe8XFm2W4Zbffq4UQ+4M2gLr+Hf7XlAkrSl4sez6E
FVBqmicT2ZKMx6lj1PEDpKsdQYRIrzwzH4NcuVVbLfBUli3llGVEAYJaoVK5Bp3DkO5HJp1ON4pP
BThNf32GiO7yYB2MX04xW7hnP/+R8l0NeWUgcbWFhwYtMR1lKaBPkQeViI9UzGaVGFAKzSqNQQ9b
7ILCJbehpBKXxfC7JRhtNPRuKiEoiBS0OL1ephjjMqZujfllojEEhp+31GYBjxMekvEkcifZAKCq
IAwvxEeW1SNjJVwXx6sobFxZjiO67RVD3MCoDD5A/3LxmqcAYnugq9DpnDHHg7WzIk5qhvgcp4D1
8EvRxgRnCtEQMbSznf+sl8W/BtsSt9p03dfMgJY7SlhPLn+3z5FXmqrumrmzaMbpnBYv9LDd3NNO
Q72c960CG8ll1ohjHxgtO1RLjjSVPH6pd2MaFFNBPzcCA9JgRMaMhEptRN7aEOGTUzX8Gg9QSTaP
FUS++hkzMgFbmdVcaHyqwv/c2GLxTMXB2xD0F55jhJ5OZXuuAerS5XWXxeikGmsOmaXt3gP4GQA1
VhsUzRcZc3dizovwdni/JgNZoRA9ntEx7SKnZG6MbxDjQqxCBfvStwFVijS6zAEs+VuGYpWQVRGr
XIqygZJWlBm3wP8Vx2FfBjj1FbjewovpoP7LmS74F1LyqOKYTrg1QX49rCxuA4jb4bDl8Po8pA4U
qsLcIUEO13FcZMUv8TQotmNe2Q7+iPLuc2Gm1pGOMngUHRRE7H14oXVD9X35gH894IYIfYJS5Wx5
xU+RRybv2Ig2TO+1p1jxbGzSC6+mtHM9WWaol4yGf3s8GU2239S7Xf7lk2zgB8xHctLpHvrxwgao
zAkxR6iVzUAlc6lXuy5nB9Lfvd9Vidr3lUP08dSJZQGApnVAgewuWybVfqfPy97FoYTqDZeQW1V7
z8fCvrFrunw8NUM0rlIXXGL9eOEVdyaAmiuy2MxGz8822AwJynwt8qQuppqmTgomz9+SiDJHGiDa
DJq1ov6DA43jVWvMR+WaH7r0CyrFSaqQWr+Ji6SnAMRpavyN9C4AkuwbJJWgRIm0yI2dRGrLcINY
uh9VmrnHwNkOShE/ssv+3K6h9MpcrbOEmV8yoFRHXklrI4EsVOZlO0Ts0YG6as+hbduyfWe6c4Dq
fgr7ssmhr3Tt40Fh6u0XxO8QjJ6VsUYGVgN19L4emo7KTEVvYBmdhlXxCX0uIEcRVRIKGWXp3mLJ
Vdvi/nrDY2X7if0XCM9lXVlRGiGX9XbipqOiB5buEeFi6czQ0rtIPJJ8Cb+2ABz0DalLGRV+J24T
5aqQfdxrtfiYf22nNVGCAlT/NxHGvI+mS9/mXE6bUmNxGCQuLuCAHL/pr4Qc5mPYDP0lnb62hrma
DFioHnb8mjIqYQY5uKcuPUje2yGlXb52DauSLqaXYQzTf4zcY9st02bSErX/+ZFnNNdQqzsroeFN
u/du/zhU9lL0sNBq3ieKnbtSDz31PUcSED4Un1yh6tmZ39pBMQfJ5tdRJP70+YQqoF15uE56mYls
AdtyIYtK73pU2jI5ik45UvPVZF9/RkjqglSKmoP2usfsQtwwOobPd+vVVN3MANuN+e21QNabPjSb
w8LG3P111sw0lz0vFUyIarV7EmAm3BfKRqfi/tTl8o9T7vbSlngSbgjACZxsckXLppJJeP2ZeXzX
vEUJuyDMKxp+FnAcXg+rrK8kspJkzTnl4mW+v4xXYIuSJXy+wghnzxlcfWLVJH6W8ddiMLZQo65r
evWwdf9PKg97XGLYXrH/QUQfNmY7S0+rkKInZGO+Rejk7llGlZWg4uN0jMiBUPVde9YqVGxUcGYo
L3ZMVf4Ma/BNdJstFxotum51oYv4bPTZRzAWte6fpstqMOiQD6a0m6ydA70JweBvU6bRt07+SqaE
5MchIpagXoD7hJGhKQtgBtkeg8BECq5b7ckTQrS3mknZ202tDDaBvpEqgptkgRd2iCeEyyHgcWGo
laPcHJcPDnJAkIytyfyR6B8pc4C45G0dzDfE01ndCN9KDUI8tKIZJ7bbg1Qsz34c21heQ24849nh
pdd3/UNZyjSbDVMltRWrF9Kxk1sPiZOF21eX9Zyfr406qjf+mPKlAK6v8dVNkGmUDhDFdLMYhHhC
BcrlCoAe1viAVB6A/Q7odml4vGCaGqAZbbn7lT+ZgT1kQy7geEqrzuOVgTNMexJNFSPaW+nTaKk3
dXhQXYVWYz42tNOkq/InEUJMxQ6SCTqCIv3No4ZLwjQcX43R+ep+A8w/KxgBc4RsaRRp+VAOF2Rk
C0r6ji4TcamNYLOOPmhQNJHV0D6jUGBNBmg30eZ4ObgIPdKc39cjIPt47F+6u4VHUPNz+5Lv70Ly
WFTzxYBvJy6w8JbSu/c2PA1LRe1lTJ9iOaoSrnP/G/EDNBx1Qmb/bBqTHVszkPUYp9axVJi7UIor
mp7bBjTt/Bs6356SPWdMtbL6AYcXao1ZUa9u5kdktAgCLR+tSFFXTqXtp/gi5t/SiV/dPq6QU4x1
4XpGMFxQWlqXiXm6YkOS9igb956mAaAtwlzoKOedUK+31ASUDDJaVAb/rW9vmoCKHjKKJ1hwyqBw
UHR/UN2oU2PGeuOpmH6N2ZV74gEZVU/13IjyUIYVvMLy8KIcEIw+dqf4PLySaK9ilwB9wIaqXeC6
rm7HbTZ4uQd/1kldZu3fIU2Wz+IFmtAqgFjENm5w3kVcfD25YF8sDsbCkAh3wh1gN6UZ3L6HNIa1
FtzO8h/vKIjQfoVIQ/45pwtN6R4nPtTK3qWvBTFGa3cH2JJhdOYWYekmGSc7X6C07LJUmPIfvS3m
NxDlCtdkIOMdKNJdAd86r+k/NF9EcFKixUoVTI2iHaiYzpDYXkfGbYE6CR2TCK6fSUlSz64YNbK0
+j93z+jgcZVrnVzfuxpANf4d8clyl9ayoM6qYEHrydhFlF8V5mmomAc10XGvV1xFLgzC4QQXcDL8
+XE/4Ql6VVLdbHi08vYtSgJmE8zhK4tANOBm6ZtcpfEl21vw/Q7G3JFhT1/08rXKkypUnBVnbAp+
vINYGISY1mskiorfVRe65mbKpccueY4Ji6q/FJd2n2obf4aZTZxnXgbbT5rqZLONeoKAetY145O5
j1/Fp3QpEnZ2Rp9by1KlboKrEqqXOCf/K+BRnbUvbuiZxNGUDiBdRonKnm70INeqqy6Jgv2E8zOy
JG0CWgRflHJvDcs9FHZivU4qUQmRhPMQofRgkj7GWPRekm2bnZXho6nNkbY9qrNW6nuAUJM/iC4h
a93JFu9YPYp+/rPBJ/wUmomiE0TCHH/Wiclvz5Fg/mTRGE7NgIowftJCebkC5TPIgCv64zn43bNq
OpKmujVbaUYQ5ael1ajxwGk4Et0+CNInHUoTCRFL3p+gXxoVQswqE25ozDEKR6wlSe4SvC32Re8K
JOVxf8wGKnzin8DYqHOWgMFEaUzvGQgxTcEZg4v5xZwdocFFAuxEKGZribqfbIFmLOVJAtjLTnSX
63QbJfN0DECjwNodWVF4rVG5LnmH8qduF84omQ4je8u0ap0YRMfkEHQIyT8x/F2EhbOH8mcIEoxb
LEr4Dj9R5ztLNUe6DbYht2GGAPfYnzPRWYLN7kILsiKm3hxgW0cSeByw0fIPkUBtA2+Tb2s+DhMP
czTlLvfrEXZ6qidFMpk85A8pMSjR+GcZj8hkOaPoWKhgiiq4z9C+/ywKq8utPBnE/1k5Z0ymV5sS
93WlvjfhM0xI9+OE2Vhi87gKcxcN1UuB3WMxQX7p5OYLHKd6MSLCApQuF3/lM4V3RsfJS6436ZC5
r00vRerIXsYg63RXtgBb3g+FS8973Q+Ho+PmM8MurJ2j+iUDT+CvdPlPK7hJmfexitrtp+zk+EP+
wya+k+DfFFFLGbUHjVxZj16hIPsiVXUTDXqnlH8WEUNQ9DplS152D2f9Wit3QD0CrMrPnScfHVbE
6xSxlnT8Fn71wtXoERyAnBFFNdH5wRA+2HCWT+NRdsah3JLmdI27/rmNgth1UPC//T6lyJdKFT1F
kTJOdsVG0H0YAR4rC7aOkfJuPt86JIvxtCvDFnrWGioeIOETyxMxV4qq/9pdGdBf9E0g9iHMxGh1
XJQ/RfhuiVMsra3C1ISnTnNtmGnmTFX13CzZyLvl1m62odKvEvmJ723xA7bJCpSjw7fWWd0IlHA0
qME8F6jN6E48qXgmMAxKBB5IvhEklo+Hl29yKIH68poGavEsGojgVKTuvUP5Mb8iaF8RuL93Qd5u
MsujeqY2q4hd2vJ9NhD4sB8FLa/tatozfvoUFQaNAROfmM0iK9DEz78KqPj3Hoy489d1f5rxHnW+
uB20BySxzVvqY3UOe1n57NQiENLOAU40rKPJVOua6ZRSrGKwpaLr5dF1zNmM/x1WqC17Z2Ic9Ylr
jFs761bE8/ScCkNsA2o7AQ/2MmHiBV/R+diipRIX5DkE0Wt7xwTR3KcEG8F1g2RLH94rJDvOxx8Q
qeOASmG5aKSIdAwFjnwNAMYSg/oOojQPvgV1cQcPC40ek/vuEWhLtGE5EfM/L5XkjSS5GNOjilLn
aCuC/Puh1OayrV/adtwH/5mPoN5Q5tRIwpNBu0x56QSH/fpisPrzEoQ3J7Bas0R1HULnE4nP/h4j
Te+9+MIXcifjeLuu/kyuQxYS6lDGTUxSGbKKUP9sWaJ4UzsUn+BmI4vCpJOzJGXBGVWIeeaor5Ia
k3qZMAdsOViu85UvRh8ZRg/HjaEkPVD1f3vgbNnBURpMUYaPJ0WQ91BG2rLgdlg6kLA5seoIzdq2
MZmlHG2vn2aK8GP0jhTXqvB5pDIUT4b1Xcrx7cZ4SXonM1gNfQX1p79ES1/Yfan7bJkxA6LD52eW
uvLjAVBCDB6NkRRFXOSZ3/GGo2DfsCccEjSdE+N/4NTBrykHLK6ZQL6byorpTPq1mnsOe8jhJhix
depAeafYilsW13xtQGVP1r5CxDbEb2gNB9V3bXetu+hxg/U37SQ40dnIxEKf7VrsS0xFpUPWSBR1
2QxxtROjylRlQd1KsV0Kh722Ns9HMTQmZd+71fyo6+bxkSRIzVwRLFherrKlBDvrd2xsDhhdKV9U
Ve3Cw+sWYrz4XJdjB9h6GTbLSRAe3jL5h3Y0w4kk+sm78Sl1A8jGnggqS879D54TI+uxjWTR3DDO
VgIklaW+Dn2N6muV9ciQfMWTMJ1W38QckMJzaktWBcC6YzBCqutECBL2nmxvzN+y2JnbG2fxTiTG
nXLWeF3Sx7W8KjgxWiBoTZO3DjXSchZ41nHgyFhycZnHIh51uGlW5uCbiDl5iRCAmYxFx6PC6/AC
NTYHZfOXJWcq8VowEagXIerdePC3HtETwSEOBTCcyLhibPslkc+TKIyS+r76QC1Z8kv62ZTFKBb4
64XJQ7QDWQF07fZh0dzgQfcZh8txa06viPZm3CYK+nR5YHSf9O+VUNpafI9eaIsZgvZrZQK1K9Vj
5OnYbL3FVUEBQsI57bereuOJTx9SKaDbBmeF2Kc/2m14NmAawujRw/Wtgwi+vs4giKtWcL32IkVR
YMnMVpv7yC8xD8/WEbxzS+M5O5twCQ6Ld58T0I7IC+w9CzglrKBo43//B7xH1SjFVKq6vGRg5a8o
fmzRWB2+Elp8wPTZqcb5Ld387IMq0RmwxrDsIQu5/EmXR6hApyeeCCxgUDwEQ877RhbqJujbLN2C
JE2SEkEusbM2kQWp0D/SfG/tUfPHqUD6MTb/x8M5+H0ArEoXSwnwtQ59EeVAE4wiA2k/+a6BKQXo
a9Wn3/wGIl3kR985/qFbTQb73MGiMNl5C04y3lkyeYpJCYAq5+/O2RLnsYXkAtNKfIbZ9P/EwTSj
U8MBMadWkz2t7owxuVl63VA9IEWE6exZ34FsRUbnjXX2S6ozQHNUGURV+QKgbty6b4FI6QNZ+wHK
TW32p6Iz2V6yp7BQl0pgw7hl3LtWbHVS0KhaoU9Q25sXfsTHRjwFTS2Fp9FSdM6PiS6kB30SgXf8
H6/CHBRIP5CYIhH3r/muv9ZOcqa01jl8V4NKsYyWTdWJ8KlZiJ60FlX9MSY6BhCQE2vXP1sBJSpV
xBObtCC91yNdYVO8fVWu7bG/wX7Iib1srKqP7U+Z67RMKzLalFrGoHmR7mT1gUhVpBdrfx0Uyopn
9P6T6ZSnxuWUgEQk3TEmAgqGmSR7RyONa4K4L7s8xLET5iyGLSRHShMS3hVvAC6jU2iXtKDGr1IY
4hil0w2UCrxcjqRZvTZUpZr4PHNO3bvYczI3hlwI2GUNuV5h/7aOCYcJnIbunDc66792MTrx+RVH
02/qsLVB/TGYjezEHjUCRP6TSlT5aUN7PlsT4TCiKkYCOQn4QBF1I8ni57wkCf4k2iOQEHypYkei
PNmiC/IFVm2rpZwwKz6RO/ymKk4zi3VTgWf8WXyldrMDdL+6BVlhs8m9OpZlOb/zlcIUqX04webO
l3JWJ6GRsf2iaWD/iQimpGllhJCPZ/C+etScubHWCqdX57E1JxCHlYF46rdLyq7Vtr02eOHQqWhD
leFdDmpHay9/TErBlq1ZgwptcKL4Dq75Ik9MYUPt2wLAQRMQMqmoLCIZgE/GVoK6zbK5aWjkKvgh
OXQlsruETEv6/OldCX6/GlygT5cw6wcUFkipQUNj2Ns/puOSj+AhSUiny3PjFcFOq/KmYu2jKiZS
lealMxA7jpLJUxRi7fzkm2hUixQmCObR6NSsqbVaGWX0mP2TP4NPUvmIPyRn6vmRTuQWU5DX9bgZ
bgkXzZQx+DOcu6Yrw3r51nsx6uh2W0B0m/+B3GUVyhZIRmrfCfPXEdSbvgEgVS5sWZ/P88EF54pf
xLzKpcAP0WWAW0j3/Adkl0Kf7zYHJRrwiFixlf5H8B9oH/5O56Dt1uneanqsCjx1mqzRebYKV+pN
CifcrvsP7WtYOMIgvtBfWBIl2kpAdJB2cot6gsitCH+C7nmmLA7ylXrt2xDXUxVNpVrhsz/9jWmi
9OkKtCDapddEHp3j7QkRyPionjdzCbL9Ifl0CovPey9AnhfksAtssYWHuTZS3r603L8fqOwiMrgc
7JerW6TvwpuPmW14+2vN6Bjn7/2BvARjF8rcITsgWc+0iCCA6Nvo2gkDNV7WRZBC6p5uOfxHPuti
qRL1Ogs9YQixiibq08nApmeng4ChN5Grbl/YcudgDm7lSqCHzdaUvXTLvYKWTzCGpcnmAnWAdAOy
htxZQl0Q07LhL/Y+EvoFY7QfhNC18Z023hkz0tzz1iz6JYKf1LOjMNSK0G4PKy0RPcpf/Fjf6ctS
1UGSH734d60OFqVcD6ERe7+phvG0296fEK41tPjvmfEzh0ppZgdq2mk/zS79IE+MpiRbHv1ot/h8
YZxnB0rZ7x8zktQCBY94ugd57bEZNRAlFJEj3ltWopKXTx3dG2pOjj/+VkzZQe5jL0Yk+YX2vZH5
145BFYYbGLARNCV/uBHXkERc3LGMZGCrCX84p3EbRPShmCmzp/pLcdecb6j/zOeYNSY0wKARH+pQ
58hvoqRxCMWmHqpzY0RjDa1dy2mr5kY6GyVgROHDdEc8yf0aBhvsG5tNiakAHEdHMFPuVpSp8BMO
/3oOzf9TYVlbFSG9ypPBgLEcJ/WJjbnXThzsNpF/1ALtsNYGlR95o0lGyx16xkzBgR9zhOd7TW76
XQ/WB42m3IxRCQnDRqJGgZ5Ma+BU2VIl6WCPW9YmrFDtts3jd5hvfRajxXhRZtuTF+VdNOM8Dcre
ToXb4pZ/0gpDoorOlPCZQIEIJk0lW//Htqv49bwen0hQRtgdHAh3ywY85ixaONyJ6vpXnp61LcRJ
0iOx/kd1SDIoLGXuQ0nPSqqTH5DdtVZUvl/2zz3MJqSK0tj7PHxCWLmSLbB7r22bnpzbQEAZLMCJ
WYN+w+YNfwTfjdWI2EhCvoJwP0NEWjsEva7WVTnbDfT7vruNRLK/UwLjGCzYXLRKGBE0UqickX9l
Q03suNAsOCTGeGXTfFuAC+VrfHQezuRkIgWux5/eBEi36G6pnfcrgRIRQm3wgN4PrCmT9fuhbr5z
1TSzrsxLhnRxitV7WchIw5y1WsK9I0fjJo2sXUyZCqNuw0hXO9fyfA1OBbjS8KpgSW96hOM1A0/l
+YNP/jLjSxtQxdEizhqFzv61U/dUWWmzfFCBQwtDVIUqr21MWSil/V9QjPBHNSJCXhbHg1Z75MvT
1UDvoXkXdU3D1UowZd/BDJUcNKh4RxaW1BuMwb7GyJVWkTiGR7CEyrW5DcdBjhSyNDlyPOYt1e76
514OPMKKB2dhVx0cj3mmp5qWSwxxmgvY9P/9zfUxdbTRy2U9+C/XOPF+R0QYl0Zdlb0KFyDShfVB
Y0TyiLEUpxM6qEzH6cPqhi7+zJL/1lVt9o0TZ1W41OQW9X46/AOTVODDGY9W+tJ6lQtiRjsv+uEY
qQY5ppqxGke6GqQyA3Wn1rLl0bXf8XRyjdBkF+Npk3A9Ga05JrdMmx1MZFGu/zWX9P5Ip9NYHsaZ
5cJFc2SOlg29glrJLzk5+A58bZiy0qkDorel8RD18GmI2bWf0ZXE+ZbSlwAWit9vHg8Y7azCW4yb
sV0SPFzic5UVUidutdA/fmu29yHAJKqKdZx09rmEyTlq+Iib8gZI09MtXgjZ555X6fiRgmT0suTS
+mDXex/2F5s4p2EG1GkRzbHUkoeD4PaValiDXq9+oKw6BOB33o1hwS9Y8kc5zJBSpKlBD4LIB3+2
RFnyIuo37lEHFh/6FnTU0+UtJJEN4U5IOARjsT9EjyBCByYCOb86DywMv8Qw/fFp28FCMDB5CrUO
YUXEIlCexEL/poIDShiIFdmPZeLs3sRtCi1O0uEeWdd6Nry5nCPPlltrisNok+YMy3KF2MX05vVc
ihOu5xRnIZm7W8fZ6LL5a+bcJReDAhMIyTe2bLN8tH2a9WuTwvJqvAM68eGRFshozBrkH8VL+NDd
iKNoVKd8+zh+3LL8XbT7KHWwgp57rgct5PWZn+6QE+zrpj3RbicfIWo99o7agMzqoGGw7Ff/Q4so
frbxLjMn48C0K8tZi8JVPHmALssw3Eq2U9A7ZqA9JRyOJz2BAYJTF1QzhyTmW0FCYIiIvfTBmLpN
2R3YelY1sAozmGqMvONvCUCozg/l5/v66r4OHgSl+R+/bvG4Q0KGex+/7lqb2YdK+jsPXshH1TSt
7o+FoHB0Gj45GKH0eBSF7CDbrUgFFGgsNu4dmEvh4zwHczioEjdw1JHkUX7TNaRWroE+vMrTre5L
RUoWWOlAppZX6ZpZYbhFDfVZq1NShaifhjHbqRSIhHa34GwmalyGr0xhkMEhKt6OgsWAAE602jdG
JHUEEAh+vakJqE2ribddj+y5QTZFfMVTuMPGlBuIM64x8FVm01WUZDH4KA5/8muNsJt20yZl3rjS
AfSsmMDpbZCE+9xjl1cYuSjcwh/91ZbeG9GFMWN6BOFQvaZMVjtiosoG/zKPBL6evejDV5mtxDvm
IFIiJSe+3/0UIm0AdugQG5vvq/SIIY4CHg8V7eY9lHUg8QGQ865f8/daxMl18sjZOpW/HFbLT7mg
4U0k/wDLq1yJLmgNYdbnzagOUCv9zY6cV5wFazvajj7Amy9W842mmSeWFXrj+S/KsX+KY980LG+W
FHz2LlkJu6kS1l20dvTjT26w2zRqIdZeFt1B2urMmeO1aUsw5K+tXuD9Ix97wz7E2C9DvVTJMUwa
k1LlLuNKqdge8QJxz80N0ocNpfOJsFLHOQfH4ZU9TK9WW39Wg7kimrX3azEoOvy7/qPle1nW85Pq
zByfRtwqN369z2k1hwWx5Qh+hLA8b5uS4bZT6gDfGrAZLKRs1HxDwFyRkSBjzNENzotl2az46RJ5
APUN6MX6BHTWKfpY86ZIuzQ+mScHa33TOrnUY9ptWjEgT2joLyy+Kpu+brkGXLvr5iyNrNx9Yz3E
fp34VmsfDXkcit57dshFau4kO9xtpfSI7XvBkAybbBVNyaD5r0IL9Fm36x3m1bEscY+jGAH1JEpA
mX6EWxrhgfgWRrGu4tDLsB1xvXjqXpuOqnR/FavzLxVTwsSTl3dFZ7Fbk1BmDKPqQdx1ynmTsT+j
/TxyCVEhzzmP1mhIslThaphrJgGSpOyg2HCP2x1PQKcd0GyMWTVVAeaHw4stSPwRxmo71dcNTviQ
j/ts7OZPU6t+Qs4ce9sHmcCFJ/7hnW/BkI8ditYoLDiJIMHV9QP3nB7CDFPAotghptmQMfvBl1jK
fG5V0qElnVN/lZtXbYB7bCD2YOTwbgZWmUDwuBA5IieIQKoG67RxxcjAog0aHyi9vOZcDc60tdal
9iR9+FTWucajyel9w9r7mFwEfymBT5kbWzBeXIy+QRC910waIv9KIAMxE8pWNHpq6HZUcE5ee9V+
wza1vqFNQnonyEjbIY3To+aMnv0pBFTIkLV6jtEeM0cEsvm2eo2jNJQbiNNigoT4/5Oc/LR5kqmx
ktyprYAuNkry5rZvZ9ew2M9UgaMyGrHfXYcVVNCvfrfV8YRquukQ35zhIWqSMWBNmDuvehclbDfj
BWGkouYPqREGHcPfzG0u+V0BHv2r2vJ/kPpmfo5q5l49e7bJEZARvOedydXS1y5vgP8s6AEN5+yS
Q8m3mhNrAUldXont9o83GA8tvn9Hh1Bhy8lH9sXt1m9cz5zgn6qur3luWa83ScwTzh29I8cN6U98
gUlJsifQbiBA03nuTeGCkU/NATXgnje9BBO4kA9QYQpHtN7K5LQNlIqT+Vk9z9LTqIno9deYAAkC
6MrUpzJe+ryfFQd/T5qtlyBch5WBGT3KDoPlF8ux63R3OAYjZdfSMU7weDQSdTeTIimU+8Lnzil8
4jIVBV5GcZSm6pG8ysJ5Q9LtZSVwWQCfNQNRu2OcnrI5R8u8CuODiNkUw17JbevmvLcPIbJChCOx
7CLz0plPRE8dImzDH9YKdDTFhTY1iNUdLUCvTLRz46fl4iLO5tBlGVjpczlcRtjrdhRr83Tu/Cvh
gQYo3tJEx/Gt0y/tIabLa7IFA6hllXd3PB4xOLk8X7tjajnm9gTDbrA5M4czy41SY9kFPkmtaGsk
7+Tp9Wmv64VeIcGMIiZrtPBoP6ZcLA1pDIjjTYWdC+i8qdDpYTzpI/ANEHPCpOpJpMYwiFH1IdZy
MClKNBnKeSSg5MDw+/oGjzSMZoGrPVkSCc8l0Y35nOp0bAjyOUNSZ4y9b/GvNaHVcKJakaVfXrXV
ITe9oxmRHfYR2A9H6GgFtOVhxjh4webriffn5UCbJkCx1nCk7ixWkKoub1RfcE8NXKGb9wlAAGMS
Hv7l9M7yt+pC/NXmNbrQt884w4DAqlJ/02HaDrAg9av7g5CZ8YQIpQeTPAGEzfLoia4LPQhXWPxa
YWZgKdSkk6pNvo1lYZzsqVZSSQlbBGrGxqIa1ILj7EV7I/2rW0ol+lfw6aG6C/bfRUc2rOGMC8+G
MQiWkOIO8Lbo46ZszgyI+T/cZCIvazHuBLJM4QPw6opCwywcbGQkeI+SmFeXnkNLpIlfG1c6ZgU/
FInHVNzNJ68n7a9bOSLjyPHEYijx4m8mzuu2Rsniqg8RJUkWxxp1Dsp239mYo8QAQlZdzg1jwTmv
xcjXblyTsd3vMRRZK3xkYbx2D8WFYNfteqSToFX9oNxBWKp5g0hLm1J9f5CaycF4lYAaI5pyCN4u
Bq2COOjHk2YHZwch5nBDNXas8QBCE3QbdU3p/IJgKjfFJchpxrExyf3qAnIg4Ndt1fTDOLWWcLHL
CoJT8D10hVhZYUZFpQjaD4Ucmktptsj/6OCpkQIn4FNvBO7EEmjqPMdOVKDF9YSLAR2vITQBQPor
yprs4kGMtpEOGctwMw/YfxbLM/mXWY/G+JuDoq/6EwRaV9VC4/P7m1ZDkNB0Mvr3ldYkBY0MQOBw
nAMLJ3IbPS8w3i2FwBYYMWofvegn3QD4gm8raXs0hlihB/Nf6XIQ8wvlc+eQtlEr01J7Kc6vLRVK
uqxipI9arXiIGl3DZNYjhDRLoJ6R0cduXNIBwwy/udA1hujEXDStPAUDN37mH3xWZ/CBgLRo+H47
4MxHCbdzwf/2VETx9gyzmzE3LO3HhS61E5La08H2pFqLtOiqzI4kfUXAfQy0EFJXEPIHcsv09oDx
J0CFpV2diAfPR0XdU8Axun+uJ4E4MS/WvcpaNaAskchw0jH06BLNq/tkdxgJb95XC9Bne/mrxgxl
HYhkDdNthOt6UXZA4OLfcRtTkBBxL7Ewrrn5nqFKkDvT80put6On0kJA0x0Am4CJPvvjy9jlg5Hq
7KWwK98TPQOoLKx08F6rasUBlm51UHSqMUEeld22Du4zLFgX+/8uSZnA9XKkc6yTe/SRZQOoXu3M
3cs5ndCZrcK4xkM0Pp96LvIUGEAqCX54yIZShG3BJ8hAWld5dN+CD8LA8QnsPyIlT4uiMpthcLQR
9q3rnE1uC7PpFmgG5RgnyPmx7iPcg5kq3aJoQbNpOSo/6VSruU4S/c0r6E4V3i1VS8i7Nl7zk/BE
KVR8Sg8omi7OQ/XLqMQ1qjJ/bAXqWEuOCrHqJVE8Oh1AiYYdpVJInlUaRt7jE9ve+dQjoWH9B5jY
NNAddmElyah+wUIQlbuQIra77zfrNqM5Nlrk77iS7+BovIKdY96A7D5DRLnDBDQCsPnw6ZJlO3cf
YbO2Zw2o+EWnwOIbGXy7du38M1LzlzmkJFp3KqlPKOx5iuNTrvdOd/WnqagKCbu75u3wXNc4AJuw
cF45mhgAKp18KiD51IVTxApX90XkPGF834S35+sFiGN4V4fqBGZGF0QdS+GFmkk2Fm4IV+yQQLMf
GB5WIiLmLUYx0mqAzy8wELx6iaw+Q9oXW6Ek/2zOjJBnlWvF8aOey18mu0vOOOmkaGDVCM+4jNHV
TmO+9mHJ+/tHGveDtPRwqwW5OvgEC+WECZi8gCFKvSWect1H5LiONGEp5s2McaCQto0FB58Duz/n
kpWj7uAbaAX2tkANUDMlRj1xoplT9xzmGQUzwkDgcmPjldhwq/NX4+3kPIhP/DNbP7oIVCR0Zjdb
GePw1JTdxlWCtA+/WYZdS0bfkEhFwmvbm4VrRIKs/ewfoj2/3+SoPFOfPFSyb2fYSaUNKq3f8Twb
Oc0a2zH666T+0NEjm6eXbg5IRUyu+u3UzTP5EMC3bkjzTpmd3WrxNJZ+cWVdCaoMB+ds5IdEFQVR
TSGYBb+Rac364vUI5mJzi10NyH4se2uqXRGkw80JgPM9dLCUBpJ7Z1z28HOcrpgTGFh6Ye0F7W13
2BNy1qOgOKN9TTxHLy065Kp2ABLoLqRwt8Cuyv2XHDavYk4kkp2PedVNNBi57p0QP/tWPCxeMrIN
c2sOOxpQkQe6sWbm6DFWpzaD8YBZE5TwNjfO1G+3uKOME4A5Pt1ouR8KAVRyUsFkEavO376TgOrJ
skeGXMagy7+aQ37AlGlLwj8aU1Q64ewO+LbUbCtGGfzNmOlLmtlXRwNhZSOYGV0ckJAizYJbXK85
32BK79ZlnbXK35cSJlEjFp4Sm5ofgfiluZ8ETufpUg0nt2ZTXoFW8wouT/I3eN1ZsO3OZTT/fiu0
7zR5Y4zurVA6zIZpTRgfHVxEV/roQJ0mZ20mmv4PTf3HGUw5Zr4a1jFyLTbp+wYT8ktEBItcP0h/
ckvgVfZQyuSdU0xe6d1MuPopR3JDq5iDVflbcsQmmdZwP3PAJiAA18vsMzo4KeMhAWBihskPQQk4
uN3dNnNOp5gsvzCvgunRUCYIx3rElkfsENI1/pGzyTpVtnR8Nvhrpa+CgKLiehhPO9VONR/JejW6
UpCEXZ3l4fl71dgqsxvDNJnrcX4mLIi4+FJylyn1s2oAgwxNztwYQ7x/uI/y6+UJG4NTe87cKFcZ
fYfV/VrBPOezSP+Pf6nvCwpML5oA890wfe5ULbemTP/NNoROvqLXUxOu/y5f0BMk28I8Uu0BRTD5
5QXwuNmZKkzYhYR+vjm36dWjyzre3nYeeHizrfYRz3IsAY0UfvRNeAOD7qvKKbKW83q4m13SzrqO
COp+TC5yMcb2VuZgGaFISuqbFlsttY6EIqB0oPUTtBjH2RaU/g2sHFCh1vLylKfH6YZjuT+/wSIB
kWmeLelY4rr4/v2jxHyo6BqeEO5YotF2BgPzUxpQizJn+kNT/Tf0Iv7RK9d2HoMX5Gohh/q2BMRo
vJMGzN3l5+hjofM7o3j/OOIw8zEYWlu9C3tmis06UbrqRZoHIMVh87V7cPi9SrbeVzHHn4OJrXDE
2h7fMaABo42s5HAZHelE/UlZ0xNyaNl/cCEtW+XLyJlNzXlYvCn6JHdq1ouigiG1jPp4NNUpUeUO
YQT7heiMvr3sXgLZ8Ar5zlOB5cvTytnE3yjW9jU768JFwjNqUAL/uFr/Xb8W9YyDGwN7ItYTjYy2
MFlsPoiKkYxoJM7semowf7n1qiXiCR8aNeV7prGwyClBRcp6UDJ2sTx55D0Ytk/A5YFl6JoxzjiQ
wtTLi67lQJZtN1dSpwk+sRlSxnznXyFYAqt5R7OYcTP53QvQFihMc4Q3zm9tA3W9B7PUfQLuKVRi
quBmC/zeFtiiLjTdEVNSmdFYzztVtPKIgFVxAnweBmMmCD8TMUfdYNKFcKD5LuC/hPY976CQAobq
CY58lgLxCuZ6dEteXznWoNjUXUSZ8et4n387Ttaz+yFl8p0usp4TFc9dbmWZKW7YIvDQxdVk9lpU
GgNqUlThn01z8JzLY4zf0wpSd/q/FhzvYsR2P2wEyo7W8ug+DvVCJkZWP8a6bjw/+ARlHRSE1h+F
unOfcxLSO+lUf+hewN5+YPes56R2+F0VJ5AJ4AjPEnWx5K/cpnHSZs+kg09K5IucdIYMMzH0811D
/WVylMvoO54C9NlWdetJzOuPXv+A6nDuD1JfdXF1IGxY/hBHj+8v0uqIs7sNwPEvuCPuf5SrCvVM
WNXUcc7WPYHz5cc9A6ReI2vNzpsxyTMNpoMckrSdl/vUAXjvqwIdHOFM+p3iFV1bsWldWvmd+ctR
9N9jA6w3xXtqMpqTSglADllMeoaaoHwMjsTTM75H5+vrukKHAZtQq9xmnNw8yeLJJcFRb43KJ157
jFnNF3ZN6XtMgtA9WdiX1DRGMYdr743UEHb0G7HZuETHlglR54sgRk4ow2oxO5PP2aOArYvxc/Cw
G6Xh/97US96709KI+jysP1kr/YSoAxrpEFvyGdLiVZztDEL4Zk8iTPbn/fVCqJ7h650UjkZO4xHx
pT2qweEmuJST8v2HY6NLSsyfscz9xVW5CAh77kv9zX0Tpf+eEBKyMdgmE/xd7TOvQ2USNSyFwDFW
pkZ5tBPT/dZmaHx0fE9fCw2SbOz9UaYwXbTRCoP+C3lqXg+mUtbKbcw2R6Jp9arcYvUjPKG3eJZo
mhq0GMNabMp48pGSMtZtOPy+zR7/3Hrf5UXmAzHkTFScXWq0+4OJkZXn47MqwlfuZwsvJMfPJIsR
ciZVl7mjgO1JOAAvQO/o5youutOI2VzPv75KFFAoHWk71P+dO9+uMnChYPSJtN9Uaw38Aq+BVfeI
nzEJu6fi8Z93T4QJ+3AYXQhrh+bbOirlrnEjPEBA8RS9QWNvI0JY1fUaGcqTML4Eqh2SJH4BnXwr
u822KpAUWaabrvIGU0F6CLcElrVCyVWji44uPSJnRgIj6ms2wb2R0OuET7b03GBwIDgLl9dOTvuN
kiQKHbPM6VDmdAUc7nV116VWq0IN4YHGGRVFkxuEiHmqF1UoTpQJWBC14572FXLRVOOL9ntvy0QM
BNpcmOqGd2/j5LUu00V2WJ8paxG/A/auWX1rmIc/niIYSyT8ZHszi9BGcauZbWpXLIPyRygYRapM
WkablnzS2DpCa+UVTh6aCTMWJ6bdH2O/ANYujlqep/vdwufgolSlcEv7ICIIWuQrEzKzDGdOARoG
EsBoeF3LzSYelb8/iVHMq4E88UhTPjDKYUXhQMc4QHP0SaoXiVzCX7LKwXVp03geYAFCwwI22Tst
53wBQqtUZwKPgcUolz1jln/uckFiPt/bU6ekaAEghQeB/PXlpDI9GokReK0qvaWeMs2fNXF1PUVT
/jQ+VIIm8NuqhgbbO0FQiYU/sEgtp1mI7dN8GphVa235vBy+OIWKh/CYo4qLb/jHs1ARruNaCUFe
Xs5sPSZwThxkcLWVax7LiAiMcQtwbvk6M67q3TjJg57/MZnAG12Zo6CSi0R96d30rYgDyHpEB/bx
mwckEa1fAYAhpH7l65MGJHpdzwdvyc90i4UjX5EAW8F12Xkd/p3Pk+K+SyNHwudFKlrpMNkfwvFj
fFdHyh0ahUcU2VL6QXrxvE+aSnDc9ALYwN1lzUHISz/8lc9Z9A/0jgWL+ccBU7KJNF5PaP/dHTvK
z1YcGvbT5xly+wvMAl58HTkGlP12DxhR8ikW0/jYlS2ZJTewg8Q8Gk99kC7OMxHPOD7ymr28hLvc
Y05KcZhfzfSQB7waEqNTb26xVmHxGRo/wiTYA/tlBJ6a9m2mtiqXbMYQd6WvTFH571Z0/aCyFMDx
aXS/4mg4LYHcCaV2nySmLpXRNp5PJO25Fh6m8ttj9kTqbo+FaZCINeomEixz53L3OdF3r1dcBU8u
/gJCZsMqLVfYsbGreVW3n/JPcklh8ZxDC0XPLL2oYa6CnMTY3bNXUdARSFHyTPk+PIMOjjK7lnHF
3DoZHHtF+iQ0cuU8xVsIeYaf7h+f0wQJkd6Wd08fHuE7btcVWL+4OzeDqZLxwtLH61Bk/uTQxgsk
kb3athJbZ/gnLzdHUqnA+gw+gmIeFEsQYMFOK6ykWCSbK7CBWeYhDiwE5adj3MoouFzkBTybSC8U
r+mbPKMdfrFxop7hyhhqUgD1IqWIAv9m0whPiADlCyqvyC54tCTx4WJaYxkTTFH5TTXFaPz72ToY
AW1K4IFkwZ/Z3ihrqsLvJFm3kxw6+r3213uk7ESwOqzORO2a/zJF/fbKG4hc64Z9C6Ng1SFgWa1T
O3vfSXMPO2ddXLNAPHOCXrpj7/Y+hVAkpoby9Pj+Mo1u1dk1pDV+Lmz2YyogwfAIRkSYmVQ4lqv6
i84ysq/kSLVLIEHWOnMCdDKxgDsYclLTnIzQg8P6QR1beuiy9e0xVsdZqDbfNi4ugOhu6O1C8IWW
9/fCy/2P+t4GOZAz77cmbVredR12iDy7haFzcBwzFlLu1bW23UzFFHhF3Ag7Mt80pvCDHLkheqxO
mTFzkvBUhWbfURu+Iqt2urawU3jVmrkE2E8TatAkK/qXU3U6InvllOoDnpFRVDqXyvkWDFx/NR1/
KdDh/7TVRzVk298idWeGGypLdP7Kj6uzIU0JMU2PfOLkGr/i5SsWWCV2FX/uTbanJ8sZeJtQbIQI
NnNHF4xyXKa3E18SxkadxMIgGxgSx0TmwZCg3/XCQR1CA8uixmlqdiO+XqvnU1yrOTMCHgf5TTwC
UV2jJNzRYkHM8CZcr9aLkQLA9MN4ZGOfLguo2efoxrb2shaAllFwsGr4BZdzWi6uPKikTYm9U3df
V3/KJafj5MXUgaTWJ5CEILax8hadlDJnW8bXYn40VGyexqrsRQw9+Vt5MF7zWaXE4iu4ecLr9LLk
u0Mlx+4Bi5iYG2YhIa/Wa4TAa/OgAzWazViB8pAF5DswBoubsVpwUVAeM5IwUusYBqvtbdzHhpgN
PuY41IorgN+dPr8K1c0qNMtuh5H5nCYP2dbTmhFCwsa7eTY41hvxkP9Cx21rpcLHq0R+0CreQrjI
RKMnMmwufg2b5XTCuXTD8qXUP3T5ihGeO9WDskFAUPJCNbiQcvkL3wLW2hX1wTYejVyFPBmJ1Us2
inj0iZmYfv9VaztCaV4Heh7/bS1V6ymhl1rZAAPRZRreWHDoamnIVLNAeh/kB6KcPGQ6SG84ybFT
4Wfueuc9r3mzprLIuZsmOgj/6mX83QyIHYQDX+udgNcM2AlQ7m6dSM15rgfEf/tJSQAZb/58Zlr0
zhtPYxIyZybxWE5S6PxHTTcwNOOQFBU6x+ORP7sfxT/9H6H8rNX37sWENV4qt8eaMd22muWiuS5E
+VydCrH0fktGQ5lDV0fIkGQG8+15S89sC3oWZA0ypCD+d7CCdZtiDbhK3W1jqbTIpvlolKmynf6e
yy5VG/GydKK71DlsHwR2c0ABlnAA9I+YIDESgXnMUwPhKGyLR8BF4XEYCWBDpHUinKn6YlNgDyjX
FHoKymX9O0bY9n5Bg48vvjs4ib07mBBrSn82WvXpYe/2DrpkRwn3BTcAnwggZGkgxKv49RE79/Hf
u5YL+RWN9eiOWHfyzqG2XJreNEiAaYhnOIvd8dFJzfyXmLQkJPODQTPTWxYUyJy8/8aPOKpt2KFA
esAW5cSB4F4BXsOR0fjo1nvf1wVfDSIE4X+2b2mSMZ6eNBYes4HBca6bOMX9+bNzJ8MxaSaGwhwS
8BgCqrLDRGqLLOWOm0tS1kwzZEawhVNmt+b/+TVcGEFP5zUYZ3KC0d1zW3I8YNEG6h5gzVsw3ysd
SoKYW6c8xPk1J83NMABS1b1XrT0pUyD3SMOvhTeaLUgZYFi0nY35b/+zU+xVHK91Sb5pGx3gY5P4
QUA6DPiRPa09h+ZPBwnT/aMk72Gud1p7A653XD0Q4ZvLFzMpJOOpnphvdU8pXjBqraGUSJPLk0uQ
5QBtlt/QrwGqpkebVYOopuofh2lbve37ooEp0p9F/pIzQK9R7b5RodENchr0C91WjBjFSG0oZZvQ
IfnnpYkkfIWQwPgi2G1WzQQWeGEVKafqhPWNsmBUWexKBM9HfmlF9IMz1ka1hRcNDweVTsG3kgtU
L63RGI+oz0879aPu8dbRymVONsbZ+RsF3LGDvctz/m2tvJCkCNiwUApNCB9bCOvgWkjYrKq5kYUj
+s/bppr5sgoAlNDCRP0mnRg5fJ6Dt02ySIXLpxMIoe/Rml/Yq+HcthauFfgg7mMVl6L7a9uMUHQE
S9efm/LUBnk3w9DvnnQi1bzPl2rOm7Dtj1CdnAP8kxNFXMUO03qWbWL4yoHm5Zu7qwjzdYb0zFBD
YXeFeCqpwr4Etlyy0mDrIckFZBobl7ML9Arc9yb3JCg/seu61xRGDIEm3J0kK3PCjxAWOc5mO4dO
W9F59EF1Ydx760yGcKZj7edLC1uSAYB1RXcSMamMW73UACGvSyklJjV/z+xVZx2qYZs9vPr3dOgz
WSz8xlY/FhEfNYCKRsWiAxZr8gm5hJdXr453ojIDzvVmm6cH8IKZaPAAAvovlkbMuqZ++AwdodGk
4fpXu2/3gi2ZxVRfCIGstw2CoxaG+h9vSOMbnfMp7QWYhwB97gD5V1pLKxh98zstsrljm8lNio3J
kHnHl94aAG0U/4CAVUvLYMRbfZ4NjLoXOTdaNvZQzI80kc7qmoL4btAawzEsMWpSXEOktfONfyTC
/m9z5miJJ0FwyRNsa2NCEz+wEmY6us8HKznLoXJ0VHsznn86P4OJdrgcfCA0yW6Z86JIG3oIhEYr
7zvZAiFcDFJEwX7Ivpl2AsPyzp9qlNwh/FqjGdRNaNTVeK147To1npp2/BduY8tpDqYYIFnDvk0l
2wzkX0SxfEhZABNF6T46xnF9eauc9xZ/LaNbbajaXmKYs8FKAGlVzqp9eIl69hbDcqVnuPW9zIii
iW1oJ/MYA2wvjKhgbDa/i53YZHpzQQUQbSI9kg/lpmVBrGozzzFZkPH0yy4PbjDR5lTbGGpmplU5
NaOvIZw3c47Io3FSkA3jdZG3S0uidFYpPwSiYsEZgObd5IWfvj6t9ojHOLeWduZKkcndWqv4+57W
O2M41MgZd4BBj/E4LtMCDciDDtHax3QmWuoyrHwVI1zHv/rDMq2Sum8W2uO0tRDPHz1V/wlMWCUs
KpqrmbGjETc2Ouw0fAlUof7A7zaMT4jZU64FNNhzjVPwttCFeylCE8J4IGsfW5BPynpsLB995nBD
HNIeVAHFYtkBo+moIQ6aak5IjFV6kwo15tfzo9aSrAOva1KdCjQ5iC2HdPPa5DapBrPvs8yCXBLJ
9J5w3SlG5ud3RQnXrnhAvDZ5Gv6VFefcxAHHEJJBgXX/zF5S/EQ4IGfSMtmj72T95fqKX4V/Fy+H
papAJQyHP6KcI5AGz1d90mMhEnJITgfv0itIZHbROxxMug2R2j2yz3cd76/N3B0TBa0B6XCieA9K
5GeBg7QQ6si4O/nSn2lk8dmbkFr1nXU/U7z/K9qgx/7zLvvLMPpJMB01LH2UR9P8ewMmOQfk8XDe
v9jgpVp3FAz09yFAybaiwnwLaOEo2iYjES09VbDJaP87ZUAGs1jw9xiGOkKONa6gjgs9hfiw5VyZ
dKC/D4VeEmAausNv7/m7O3o11yrAPCnEoDjwvMdJrXmpEv8ye4zS0RjoTsRgHCsZzaNAyCtrBsz3
+tLu0rVGVQkQ0i6o82FQy6LbumDg+5eDXLUJWJ1m9REbOc8K0RqjmEmJ2oHitFPfYZ7meVjRNKNC
hRQrhpiCSzPstJtE5eZVsfEnBGjMY8snLEko4f3k1gClnBLFw3zii4tW4WZW6y8EQj3hovzlk4Eb
mG4Ja+UQ+u1xOaIBwoUOWkLKmSZ5Zbl6wUQ4A+EqeeHNqPgqebbc24iUiIkfyPo0zHglgwR0M1Ni
1xOH2CuQ+98apDtGEosApSlaP9Uydow/9pE3sveGYVjD431NQ0zMTsoLe5n7UKoPGwFmDeOvooME
GgQoBUCmiV1/C8C8WAKj9BDz/FJcDWtRwhBdTfz/BBw8d6TFKZ3RT3FS7x0NpdFUnuYGpy2YfrkA
8xtWbLACm1iYN7cvuZ2zlWCZT7esxF5F2Yhyurxc7g1VsNGQl+qIuftNJT/0ykhAVCVmE5LL6KCl
8udXzBK5JdHzc7eLsKq3507ckytn+dsCuZQGEHxu9azO+gM8Yj/bklMN6ykJkwKSnPnCgXtcVQ7Q
ztrjHK3OplqJU+A0QgE8wvE6ot34e+9FcXqK9U/MltlqP/c70DuGvKf1CGbecg0tBbff3HyGsYrQ
1B0FD9It/XP6XQVU55ejwkHyJRYj3iT9WPLfM0+LgWgcOaEw1BVJt9/IdHMO3t/5KmNEcZ9+Y0Nf
S2eUKSjakbp5smZqgXBEKj21rYifkXe16uoUkfQDLTSu+yocHr4NARTh0nIBTztmnKNKlapZuHAP
eU42sB1MzDyLJkbi9GIjxpcdUrMvAhClFrmjlGlgmCLhrqIgMStc/MbDuXVBI1ZYiibIY1EiJ7Vf
2UoR+nemeBxByQxxaTBB8GI9Rytjp3KwXeLm5P9WXuiASmd6VwLlfkLfl4chM6iwc/PSqaG6v1jW
3A4GjSd1WYzK6rLkSaHbRTe6EZIXW/ra+TF5LZAssTm67skJpvejJF6F3xoL3Mrl0djGixpuhvNd
HtUa9md66GEOylQX+ki32DbSYGzpBUSCB6iJuj31O8Yp+pOTt4sWIBHY++cwCG4XlQzEDPBvEGT2
fY0DJ5AUpxJJCSwFtT7kN/wFZ0UxPUY6GAe1sx5NJlVVmnuQUpsi+0IX3Pg3bE5IYOLSa1Y92kAf
lE+FN18QSVfPrIfo0Y0YJF5OCR70rflGklyYiBShsfu7VBL9CC975P1Mbup8cypYtc0DPgUpjVHx
wPkxxatETIl8ywLwZJCoh5cYdotN6seiDc29xETkW7IlE1IoAYAoJesBBrRbSjMpNouH06RgW4Dd
6OVliGWQBgrA+p/fVPdp2AXd4WVFPsqppGCyJD5y9iGDAsPCffKUuOFiVJygmIbZrHPJ8hYz7fyt
eqxlnK70E9TmLk6Xgb8iGzU4ZOPBeE/LA2hJ1dvs1gRaJhLTTzNi9QDKkVaKywmBmuRa7umQQ9H/
9ZKjJJyZWkQmHaMJ5TTotcgmfWfqIZOciybOJ12kT5H/52ndc7KByxG//3hN9Xidm8/LNzXeyUtK
ScdwTMFbgTn1Ufd0aTeUQ9rGkVe+KKqe/ZEonJC8bwizBLlEWzkME+dVvXxJ323tDkkPh2Z7nvtP
AIcmI3C+ZgVxa1WehdQXnr7zvNqCLag2F++vGBC2KaUZ5wky4DuGuBa8YwFarnNyV8IErwdbUrZ8
EIwTxQeSPmfd4saIg7twnVpuFzXfljsXGJExkfeHzxX0iyN/YN9Pp7tpkvEee24tpnm3C189tOX0
HlDqqODA06jruaETatchm+ts6lmy1GQJkgw4BYGHl9R0EJfhLkPsHXsS65B1fn8tA6WDnSOO65Du
8H/+ZLl+t9u0YPmJRdbLHprqVwUp24U6TfEi8FiWjUjz//HeO/EBeTDLC2pZnGf4xhZ4EP4Iu5+z
qvw/B3wQ8WB6rGPIbu5gLx/lNgcYuqbbUvdDTS+aDqhBnkpxELA/ZHZdxJ1w+g3Cig3BmMCuR9lb
ZLXc/+e2QWWRf+sSBtcPo5SWWxF29UWFzwOppIRLxlgtvt/2sLWK8Y19J9usQEUSmMVky2Rm0HL0
/ilE4zUq+K+b4xqovz92rh+l+fXkGW7Rl/I82zmZHNbbqfKSfe0ysyCB97tTv/oUkosPHYOAcoMD
nb533k/A/g+LBHFL4OLSX7VuD+QWVSgtQ6sdkQYj1xUaZ2ug5i+YuBZL8ZMJlfQkcGwlh+4ndMCj
krAz+KFagXPwhwodTqLiU9PPoMDCBLLXqKTBvVsIFKLWkn0lh9mjGQRtLdqfMYgoq61jBRwXqKXJ
ZfNHv2MobTycU+5cFbbYwurdRP5nR0wK0VUfWp6Fd3nAJNVKSibGcZHW+P6QcXa+WLv1aWtCDFsa
RvgrPorWdMlIC0d+0d0Gg1RXsQ5wxjyrVZvYXpmjOWoMzyqOZA5UtipVJRzAJVI9D5qXVxw0Hik/
S+tzqJ/AxKgsbj759Uuhqa57drtegi5ysidmwLw9S9smhyrq1eiLUlBFeiYwzSIQpoLah0DaaY0/
oSxKIFMkzpRjQW8UOLTquamJDRjh6ye6c4G/j5m9UqOeIL+LlZ+6SvtYwbiu4XhxxHfOAgtABsOK
MmT2COak16c7Nx4yWiGt6bl07aox7hi8saMiON3TphxDVrPGbDbiMuk5sIkELqhoI1NBTn7xhmFe
prhs1Zwumjypqba4CTtsfJd7ih2XLdBzEXweBHS/E0Xh/38rTrc0uJCrjGkuz0PbrUqO+YlMnAkH
CK751xAHeAgmGhMFZZK68LMRRflbKlJhqbRTnj1Lq6KI4tabsr374w3bM6EHTopGXBDBkoXVr9xs
MNKaCJmTn0qR77s6LmBIE2KDXx5iB4LYNK/Xt4aNnphM6voteUe6sKCDURCfphZaDDV87o07ycKJ
G8VTeWkLOvnToCIs3I4GYQF4Vpb5nKHyslyB+qtBfnK/pNnymHmtNVzcDY6qj8g4vnx8AFIUnqck
0wTmtNawOQe5SqjPYroogmugKdFk83xXmSdOoPdFNSgJ5f1GTWvxWsjORvP0En7Eb9ARNYj4Nn6/
ObK9s1pyo1zi6k4ogw/QXTxEiNA+TH6heBLXSjt5+9GXSlo/UrkYKAgftEL7D59LvrPFUTcy0eeW
J0lhG4DQwpeHN9Q2WhrWEVRPRj3+v4LxGJ7+pVS8JeR5UvMmPQ66eXrRZdSDgIGKQnb2KaE0CYxV
BGBlFUZlH5hGxvw+VWzYViBPpFjTjVB8Ajmt0WJskhY39s2enVIiLYyH4Uf7DDDLY5atTUUzdeIU
GrV7Pexvx4lJlf3UU6se0nY/XoLj8WLyOI7Xmg4qIfMQHYp+kypLsfKeRXAqd5eNbCPaEFob+sqH
2XBhIX9U2GQrI3p3OcCh1cBl61Npdy7Dtctilt6QYBKwLPAfaRhg7G9j950fCEWAmvIYD23bJarf
prV0vOUIAzTV/CigMrT3w+df4x4hIVFCEorMraehNYeNP7aQw/P+WBrmtH1wNOxP3mWoEd3j7jKh
+5+XYy/ZooDQKTDFHeisZpW4Fl6LrVqT+yIfAEhvx0WAE4zAE60XDaOPAig8hXSzaD60ZzTGyjvA
7keBvS6f5wqSBCVB75L+pO7nqyT6sLYdir7jSiQFYSpF5JTCxJ+nUxZidOfvVx1jzDQE9ZpeYHKm
R15MoKJYXB2fVfRuDIgwz+nxhC7J9r3bt2tndxCaaUDxXfeXxC7I2N1PAn5eTilVeiyVvwqenEIL
qJyikQC0FYQ33JQ4j688wY6dphaxh/dGQ37qO98c+I0E2ODFyeXXS9oV28Au/OGSyO97lX1vP8oG
FQSgavTHx3SvLNBmIUrINFYxh77Weh0vWywDGYFalNr4j2tuTxwqEcsXkF+S7/uzxf/tQoljsW6K
XL1a8hCLOxA+61UpM66DJjqCBvbnmssbU0FURM0UTrQnba8XUuLJVcCRmT8IyS8MiXoaL/tJHPvq
k92g4c4Brho9txE83/c4p8NPRpLDSFIzJwVCuSHpZ9Pig1R2L/kzqI3SHeQ60ZzZgJfnF5vH7dn4
8Aw58BaKS4SHLwVjE8ep0lFZNwba8Xck4M+sg094d9Wc9hfPdQtoRYUDe7x/2Lj7vSw/qbpYjKbx
qoX6tAtnrSespBiZR6yCoUEmGNBWoHPaCY9BzbLbANKQdoBZZkbbaQWf3tiwDbhd/wDY5J3y8PT3
TxfcmnqCagGP0TY6sTwTaexIGI5jyNIZ/rYAs9M3EQLkfisEqmYabhpuoF4EFXEMotWoGkp+EQRD
49XoAqfJ7D7jthg2dKi7jqxLqQyuTrUNNJhy+M7lks5iQWvjGuTFCk2wwrBqrUOaWk8Y/gj4NgQw
yFemMT7YoEp+/WtuemIPcO2ZxjkbG6nWGyTVlhvpNH46Pz1XhCec2uSllVJyXL5B0/xLY8uXlq9e
KIaK+GU3wlnbCmpu8LzQ8zPfketCH7Rj7s/J5/9LBS3zT9VU2fINOrtsPkN9tebsWU0LXhMk9X+R
F/n62Ejay4umJUPJcl/b5YB7TwylKtkRtkTBzDTI9z+sYIuFiqA+57sj1PFyGy9/Dt+uB3qUnBQl
Mxhu6eHUxau1YJVlTd/Q2JVU+ogpDDV0LcfSL3jPZEu+7KQRFXX31Q5YpA50+YlpnfIyqyaRDy3T
haV8gM9Y9S9tbTJgOE/+pbDmlxLWtW8QNRGXH1JKa9Fz/be8BbBtK8MtMNbOdgZc5yoKlzF62y+t
eBJHdLprtjlIWaPbetOtU1BFhCutllfT+fELo5ZYymqB04rodvTGjqnZwA08/MgGbfSP5P8HSupT
3kVVbYtcJ+N1GtR3B3O5+Vw7qDHiKhtpsD+R/gddx9DH/VfgfEFMKqiCkCA0SZWMsOiwQC90NUcZ
1fMUT3KYqk2BFyY7rY5O+a2P/G2IaJaoEEI4TblWtBQjK2EnQJY20WuWuGWL4bE9AClMAl9aVvTH
/owWNrqdkGp4aTp3oVqTxVSBan98Ar0eMODGbz7EkqXXaZC10sST7qnROUu4slFm8hoI/5++WU6F
7o7P2KQ0t3Qc+2DdyaR7SJXe7KvYidF3FTiZNyaDVXk1nY9ASZ68nAy/P/SIMlL0BnWe1bW5JXbQ
AhpkbJLDbpJVkskniHkl+YJeWwnAmwD770lbGAkvXTRbEmjAFwq3EUTjwAtsjmDMpEt0XvFIQnCU
c1mQEsY1EMOSqofQIdjvkWxx2WeujobKtn05IDMyrFdvBTmlrtBsRLJ9eK/hmeFwhuxq0AjmdVCT
P20UN904zj98TEthUIdOfmKkwNhI3aHkN1743z6Ut8CGfrbU4iKq2Hr/bctIhog/tFYgJ9sUTKaG
/bMiuCFQTCJhLaFRvD1o7dBjL5pciyICUAoHU6YkI1Cy9FkZfmsnZ6ChOZFXXf+ThmaF1hRlAB+e
D/kaGesvwxC4Jt5hXySJjC/Av8C5ww8p+wdsibzhJ38fcTjJ0CI3XuVAwEFJhwQcxyHhnq1I57R7
Z6o8QxPGdZTwn4SsHOqUbfJjNw662frQFnMHTkK6GzvrmE4Qwqe+Dfz/fXA+Q24JbBXpAxYXcNzu
3e5tdRJd47/a56oTZNLV+hLt2IpLmg/t3Z81KA9dfUrrrXqwIve+8HyHIRL62bb/oUyssMHVqxeY
Cj6GOBG1sCZj5nimi3cVUm3ljIcRK0/wYXWu1atNgElY0BRUs1P2r+o1o+bbrsXvoqWgyNvRj5+Y
6giviBvaPk65JHCJu+/cPksoDyUK94SszH98oKXzzPkt4YYL2zW6rRAsFZo6Dj2jw0YH0O5jw018
GIfEPkF5GrfVYgGHsxjyVm+oDWIiY/3X06yzpigZLF9yYd7KlW9xM7sbcaydSEWIuHO0z6uodznh
Cp0FTBij9yCkCb5uc9qS7vJ1JKGR4kjvRl8uqg8MChIymqiaRyln5hwJndA+r55TU6RcvIyHJRef
j0gRTL9RptD7rHTiiMyXtGEwX5RZCvnRyVL4xaFpuZbOL/IR0n7CNC99nW8vaTWh7SkmFp16ZtNV
rympdaxKgXnVJEU+ytWqEy8HLPKEAwhWOxpjWVh4q6ALZA8u1oNdnF+jM8HBLjdCtyaupte2EygD
8zMVtyXWDmNeaYMbDLZZyoVAKc5j482oesAb98xizwy89Bx+RNPCltSWSjdhmlOXw5v7EB1SFOiz
RfSVcy8E+Vy2wL9Tmitc/S5IjaDoyCHaIB/10vBXab9/epF4c7mrpa3MCGebsXdrGogITeMQApTb
bDcqXMvVgkUCoyRSeLENOiGq7XFt/3PTNn1VwNVCvSVoWIoZKgJrN0mYk2EO7y2O+pLx2ESKK/IN
vZ6ws76xEZr7Aq8t5hOWhf597Dutne4r4re0jePjWtCqdOauRCnwMgCGdn/PAgSDXCglmi4fhxOE
3LQxzzUYwguZH9CmuMtGdMJa+UIXGI29xcWrtJ8T89Ng92POX1pl+EaT1fOabpX919T/3VdO8RXu
Ns3okoYilYb2kQOdg6vJr6qr7DjjPco8BPgHpfT98A+PYALicUuoGWchMTEPCsDnejGDZi4Nw7jG
5a3W9rHdX+J2np3So7s5kCYZUqlJhCr/jtYfYlJQkKr9b/Dx8Hs9ZU4I2u8x7XP2mFQvT/MM3v5y
zmM+puvan1gEVN95aUfEpDI8ASOD/2tEPHx2cGzey8Ff/rkzbcA22VDVME/kTgtEQYOFSh1rzQQH
rBZj6cnyt/Eg+kM1m71/6dCgyiufU+AeQxllLk6gqE9+oFQ/WO3UpTaU3s1BmHsaSzs6drGocFzO
lnYOEZnLDK3SrI3/4aBs2GLDA78GQD1DXbcnpB03flQ+CFX/teWy1g0BUst5hlV0SlKwQye/aT/e
i6+fI3tw4P4qw2uK7OLzAwt4/m3+AAlA24x/dVnGKyznn54L4RjtmacbM107ZUW3Z8mthQxLJE+p
TrgmwCoPfMQEeyowxuXeSYkxxlbdc61lNdwJBQgIXhkVaaFndAamRTZO00Szdb3ffc5mlWvhLPE0
SNSLTleZU1JdBt2KQOrA42uL3QSVLd8G+MYRo6cdXmod0n+4IFI5Q0E6Szj0MRFNLYNEz1d0nXxx
SKvZ+lDywXwxprJCT2Gr2QtJgFEDVv0aJVc0GR4s+JyPHECa5KoipnjV4G1EbidrZErH5YGiymH7
uP3N3DHwJZ58aKhYuyfuatePWWE4zTf4p5dfZkTE4X1CKOba+2z6nbF7ryJS+p6VXm0t25rckJHl
B4w2yfeG5ep3gsfmIkBpLlyGlAIqOqh96zjT+C4XnusLNGK6PXRf9rSs++m3LNNjLpCSUWpl9C/Y
LVTBznBy4khmZSWOB9YjTNLLcuFdrenrGEmdnTwJ8R/ZS2Ku8MhHuDNUFqrBozrVE/TuDdzBp4OV
0Wmjuiasxa9Dq+2fv1YlHFdwiOFntlZ9LiNXrNdJbwlMb/V0+viL73N0U53xKflK1prx2rl5Smxd
pA2kVM2r3gH5RZtIuyn5By54vu/Jo0Y/s8ld0G/LY7i0YdttYEI80nHfNFjVg1JhtjNyYD3JwW0u
mS0vj49ghZJvOmUDEwXT3rOJzKviVlzjZj7YERY+xlxUdWtix10GsiG/DyjjSoYzck2/XMs4E4mP
xv2HniJLuBdJB1SEHrp2JlPPVg2oLRnjoASx73V5s2UI1D3wchqWBm7PZhu6Gi5kdjVicgSxcds/
eJsrvtwxhEZ32xFNUqcPMimInkfb2XfFnv+thxAc1UbYgGjgqNIJrbNbSqh5C0eASDEdOC6C5Kod
k0URJZbKLKU1QnMQc1AXopTeSqezDlEWrTVpYQtpVWw1qpul0L6eVakJacu7tilan9xTuBssrpBU
skWH/JkH7G9Z0jkhAXEB1AoxRHQPS/dWzQU4D0wiBy4PAMqGfYSY4MuoaytdUp+1nqg+O93kxW3T
eQUHbgAeGSvgl2rhkbl3mT5ZU4xYgGFtuLDtTrVxmJ/2x08WE+cXDEZMkayIMfUrI/g30SSb9T6I
qrUKJpf+AwrGftLv8Ga3s2k+bSQGiIUyWi85zIJMF00wz5wvvjSK747JuRd3ohymn6gLwa76sQxN
YJ2g7OwTnj+/USAkF6APre5QX2Ds1n3G8TfAMXeNgDQSbBBP1bij8HxYRVBsR89Z7NC+yP3EpXqC
h/zznt7ZveraTCkSyOIhNyv1QQ1tqFQjpOkmcWZJab7EsY9KNlQib78sv8gmhPa/biNitVqmVwqX
TfMuHy9mx1sld6xVNVUS7XYYQpQOWc1fuTexFDTvF8wBV7ppu4T4ubTblsqRvtqsm33sGJPrKwNH
HKbSP6QKCDDNMj9q3p6tP6xcMSpTRmN5zGPgW4ISBQnf2Drd8xniWxdjzng86PJMog1T2bs0YdPV
lvnhrKkrumBQ+Hx3xYDzBMdqnbj4JlgVbNbuYTCjiIVf/grJAAZFEdGzfWnGHNVx7wRyhfBVhbaD
McqkaQ+iK6TurnYmUYUqlOjaTVcPDbSoOer7Ll8tbuviFQL8JtzZ62MR0cVTmzo/cNIaB+/zVu3a
CI3QLD8pItlZ766s6Njj2pjrio1qRWFegv/cWxciu/ZOj79g1vUnWeWqGitDJcMtwM/ClGWnbt/O
MGSI/22feAyyvvSwIuAgGtaS+PrIlfCDj4Zr9p60zYEKuA71kcRXjlbPFSFryrK7A6iGX4oN8Qxb
OJB+NlAHibBIUjs5h7mS4x5tmHHOow17dFDSyj5nTbNBGhOHhvrs5N+5sNjCDf8MeFaysRlf1siP
3lwNOhBLaQb1s4FNDDgPG6GVLHjtmkNAsL9/NIenUOth6K/VwYU4/Kdww1zZSVQUEj9cqFMOZFyw
f6cTJGPzyd9jXGhIXxw8ORK8lAvX/qEl+DHcrWj2zxyNdpxZ/rIV7PWWNpjUI8Qf000jNyP5rwRx
pbgmhW2bOHuPhObddW7uRWsCtLO8G4yJHY8J9jS64Uy0KD5gyqinhIqnI24HCtpsEJlgBY2tUK9W
plz3Qdi294UbUEJpqLgzqK1Bw4ZRwbd0fBdFFGl4HQf02FBlN/uIt8SfObcRrSZ2VZGpIdQl1Ogy
haJjEJI7HViQpS5xFsB5GqWEGBU3HlgGDMmCnvoleUgDXPKH5c8wVRHaQiBjBL3GIjaEFw81ntmM
mUK5mFUnse0SG6Imb6saCIj25DrQVRBShX+t816mumT69H1D8aqPKBQlzYwxUYAKHnjctuDK9c3K
qPfQ8TMDmCLJ9hQBnBMyfPHnRZoHjNa98I4AR5134delfmJm+iFH3P/syWz1ANvypUS2KFKvJW11
XB05cM5v5m3NttAYWi6GHgEePJ3JfYmAIwAO/ZhWvzEzRWf5vIpdcxDsOkB7949rgw9+5X+ZLo6u
kr5gCNA76j02RL1v+gAPpTqzrUqhkMBmXpM7dgVuBv/SL00bU6gJCRZRvnkGUIWdV5Czx9xlZORc
HLQXvYTObO9eaYVverszIw4jwL0DM13zj92eHc/81V/2Zplu4xRpSREubbZUBfwX5DbgpEaOHsmH
y8f875wh4nLC/niPpa5mFLPq/XNxocAwfRveleaf+irTVnGedSfdsgMtB3LZ3ZevoPi7R+uc5ohq
g2+ex1+YtsJCkFBTgXAmeO3AlSPJtjRCfz0qBuqSyoT9gbr4k0JRyYHE2RsoW1OzZP/gJcVEsPoo
BXVCbQEvpJktCN5HHX4+/2kq6UT8JS/JQJT6OzcLYB3YSjdZXo/T4zGoltgI6VJRW7xx229CZg9y
63QE5+oqGUlLvtgt2e8G1tuE3KAYinGjJ/nsWQO2ZgCKPpbL1bi8izJVRTH7x5s9z1tKjD1ymqty
8POLz6CWf6tgzSqzEJqO21vz0UfIsh7m+GfV5ZPPhT3s3v683CZrsv2Ao8FsFegz4lS7ndxtqX/0
UH5BteHpf0ojsb5nGJ36V09SXdaKgqrlXXtPGbUGo7UOUUnIVBwcVJqQ4iXAJ4L45zasCFQdfJaM
xUjqqf1gelQ7GRpnpAutuyMK0+ZozDkzfvgr8LIa46dv8w5N8Hml+rCimmPYrk+sqiwxYcfn0gcD
LEIM4yJWGoI+qKjIDguJtxVpw/U5dc5jCbwI71leXZmiPDnpr1Mdl3B4Scxqskx0X4Hv9DMl8qVY
dy1pNJLIzbFpU8nPbb7LcHPployUIKbpL0fQ++31eb1ElwtNE140oeAkqC5Inpe0uko3H+oFjnGX
jVQo+BEKi1Cu2O9mfUsfRrQYWK24bln5h6NMXjarc8v1p6sm9UFLMrldnPpIkMUIfT2/LjP2vbLi
bNNAWM+ZMgAPr6bCu722xf3e96iIB94hWK3qBekcbqy0j7dCWNDJdU65HU2pkmrVAtDyRo9yiRjx
TIE49uisbjTe0+uDyTKl3cgumVH3ftqoZfc7uLKvsNJ8zehsaMt9LZaHeQKp/5fI/jSuaIJu/9vC
a8cQy5Oj40lR6k68Bg1vXIk3wnJiGpd7JP4k/wJh5bhMy/8+jhgjIq2jMsvMdN+nvNUc2uF6Upib
fYfyCR4746F8ylaeOmnOqAs8vWU1BUcSKTxMZUdhGHZeC2QOSX7t7a96XXfIjy+Ir/VTKH3zp3oO
9NHmVDKlayUO82oKD1AhOoz5S+HuH701tYweLQqIT3U8IIuSCYkGnCvDRbUrET9t05Tynf1gG/Xw
F/i2Bkt4Y9NQGHK81IBcdzqIHeWZZKLnXOBmr2Rs4aaBazbv7UTIpprRds+68ply1prcJ/+OSwI8
mgWxZEk8jEEBBdoY/XCCT+FERzgIRhvXkI+mINL0ToIKefkQNWCjjKn7o/Wobwt2XvjACrKIIfQN
AUUXEOcE8BNP5Qx1hLBHhodeXsGNjz5cVUHGwRj6DKAt3PAjaEL0DDwJiXmmxMd6WJ76lbeAoBC+
TYQUuN4kMEeYAsk4ej6EVx5UE/TKe7GjcRXkJe9F+DLU/UXGxeWx/HduFswbZNcHf8NdkptdGuqx
a+pdKhBxo8Hzj3RZF50/bSobIfeIE+KPZr5C/+7mW/A+m93IPFw7YHfNckc5oR9Rczw21SiOVCIk
/4w/O+Igt97TSnJfu2UO+aOOJLoEjsM/v/QJOO6RZcOS2s/GPMdkRGwYBbMzfNijpozNMRd42sLM
u4WJvzHO+6susBODEFmbrK1dJ5xRDFFiQDL08/2u9Nm4MLZgsm2Yu6KVz73D+ulKjnq5w7g5Z+kp
1jHOIcoXjKy9I08kKsOys82CNmx9of+dvhkUY+Tm5FeFS4SpgLXXuxXmjGAoOez/mH6BSxHFVZuY
4n/tUEkdad5AMa82jBNOYTtnGS4wpL7DtKCHgL3on71fZ5k1D7EGnG0oON20BQJOimfsegJ3PcQl
YFyu2HXGBiUdzmHJ8d+S7nl4KnPCQFomAj76BR3oxEx9mqz+E1yCsvp55hLQOxMNjz46VscpaEcI
fcWmD7+myBKNvNk9dF1cMlZUiREeLnt5JsYH2z9htJKqGNxnjLOVsVIVLa+ihpcm+ZqXxVnujjR2
Lq6yV89smou1XyJTKXvmCFOa8AZXWvFACwp8wds51BukaktNL2j/QbquDDe32Ai/KRVQNnMDhC31
/DH5h5aUAMFSBan3ke1ni9ggWGcco2tsxgkEF35FawRqYM6AAjz9ie/DTwbzR8+aE6nZCm2fKyO5
hG5iYrOtbIpqK8BTsPGQ/W19JEOcyeJaDxOHw1daFQE8ghQk4qRKLlOw/rQ9oTmoUHlQT71/Yzbu
peHcUWknKRCq5PbDqQ541G2yZ7FXmfRBqCHJdW6IfBx/QqZxC0lzMhiOJJFBmHnUW1msGDH1bi6A
zZ83w3Ln2TwCwre/u4wUPMvpuY7xdVu9ch6xCoa6lFP4+CGrcIuaUWezWDBg1kiidERM8uNYshAf
T/KLHHTh62gr1k0gOEHQmmqR9MBb1mDj2FihJdCIHsS01vTE5FjOpf5cKGTVIH3dzsjBLljXIHua
V7mYyAipUBiFkHtrMO8YtWuSwcdpg0xdCCLgkuP32aQTkZ7B6wblhNtFHfY/Zzu3rzdBjRyabpXZ
/51bD/Ox01SaWghdXzodPYvQ1/C7ITj6BzS1JxpgAHaI9rovWQhcxEB1q9rOjHt+9GpwCHZ1zw/8
IWN8vXbOGzY2eCrBNMLg9aXBQpX60mnUOCCK5TgcNsCk9X+2cl5/do+2SE4w+tDI+9jM9RUOlmCm
1L1Mzm++/kndEk0zaY+/XDwBbZHw8FTRwC01em4EVf5/QToXFGOBxG+RNmLXUmxGPgr+zERONHhu
PmX5nqgVMt9qbgfKazS4cDoFJn1077TEOIB05AjnHE8BrGDu9Ec8gCVUrmwV9vE476EWr4PaI+on
UrO0twyf3/sY97wPtoXNheI8xsNzi14dg5WMHZjqHHGNtMesD4/HjXQdmRRPKcJ3LXjzpar63dXr
MS9Wfkqo+Dxt+XOrXK8eyQUFeuRymQSKpkxliWuCbRRQlKU9TUr7tDR3nr6eZAIm0W3uKqcD3Azt
/E9CBUIWKR2U/Yfzg7A0GCgngQ2MJCb5kdFtaq7LM1F9+Nu4e2EICkiasW4SuZSZffmXhP1xm7i2
uzEV8G0QF/4xoMeRJQiVbGvdQvCuFWPCqsCh+Od2qqVVY+LUylf7AMX87/F8xUFd29oztQhmMRtc
2+2i7grGUsnFezrrikQ9rLEdeo5/JRZAW9y1gAtNwSP/Hkeuk4sD/qUrALofFWAHcZnWMxs59P6m
e495Ia8l4qSUpAaJPtbjYgsO72sYf6G+MGbmBRAwLW+XLbeOcRoYMS+47c3/1XAyUbSSR2pirRqN
kY0WSy5hsACR6BR13GYMjXIaP2tLMnUXqpF8dlBGH9/FRtp16fJTHlkR1ghlbAWdspghcS2XpmOe
l5+TfXJkWQ0T23TWulpinC441atMAdGnEnSer3B9ajRylhJX3T1/cNzKfpPdLopXSot9Z3CV/N+C
k+yrwfnXdSbM29noEp8Y1O1OtG7W1RrU+X6Vk5kRobpFaFa19/RZ9mI4BFWiQBDxZoWhfourAyA9
kLXR0KC2S6joCaH0lRDc6t0o+jd1PGJzPye1hfJVYa5BjAfZUz11WqJgD1kHJjg8nVS3fXRM22CX
c9gBxrYmeeQ9JzuEH/k8N2DiqM2vuXmBTl/QsIXqyx5wNj+b6/Zmze7NuPYazXeODNbz2MmIGIAq
wtdEf1lJVWj7boP/FS+HtuEHIyJ8NwQaEvsaVz9Rp7u2YAn3AQtgseT6usHIoFtrvSoqkoacrhTX
4rld8espcAJq9GjcG5auHBZ5W9BGV+dD3QzswVF10Xypx6LGpqGlZ98Uwbheq3Fue4LKxq7rlAty
s3+5hO0C2q8du1LRDZoCOZsq6P4YPLcy19vGUXemf8nc79/IRqVbNbEUQTamQEQLjqAu4pIYFTdi
L0H/VhbwbeeOXMyGKJFpbLMzPsQRBjRdYSk7nEk4CRndJpG5CwCEwFA7xeJs7pph9sTbXRLMnUIs
wSSuZV1gacjJviwODs8/Y2QfLO/BmDN4ik9gSO2F9ynUPE0t/LA5ObIbZgxHnDIDc76xdVEIRtyV
mx5CqxdnksTy6SQtylJze7WCYS2IQi2WUF6HrS2UmEZpBYEmpWxxajExTxDOCIrwu3KOrStQGko5
gWarQLaHY9nFX8uSYkIYkOGYVJUn2S0iOzEOMngziZqWNSnZTfdaxSjz9Be6eK1eSSSZZdXg7qzF
3ai2dr2QvDO6XqmJ5hj76D8g13tQ/8AU4y9u3OyYRtud1abcaWJpQryRiekUO9nw951J37sl2jaj
hBpZ8BvRu8c6NlDFcksHqCdQaD++kET/KLSf4h5s4HIXAXodgAOKENpmKEW2BOT8DnGHRIit4dWW
D5+bbrsUCUohjBrKyXrlm3u0PUSXO2jMWEMNBrLja+OKTb+9AgwdL3lq9QclOkbVM6S+joXrBgiZ
fjTu/F8Xn9O/WZ0oRY+RpHlhI6/hObJuTMaGAm2j2+5qWEQ/hqYW+Fv9blbPRiGhbHa8XnjPaIUp
afuAyaMe4Yls/JLFXmcAKR76/lxHS8M9gOoYgzhLTd3Lm8/PxYS7Mwys+HCpZMoSP1AI3TGfqyzO
H6yvok8FC9dpbVvS6CWQB8/dLaIZ5BOtPUWScpJuyv2IxqjRMNa0sbnRt8I4Yv8a2Td6tCu1n57e
VIpDoqACZNE1owOiWzXu0bV4mdiAFPQTKoDx1l24idsVSkmuxdRU2ANDj/NyJEOIBQwyK6cTOxDW
pQT18pmfwJ2z4d3vvEJkbg7hiQm+KLiSJK72FZKuOfkPxcSq3LE6Ysw2Pgzv+lnw9V7aQZgFwL8R
4m9O39nczEYg/ihrMg3At0aM2J6S4HqUAeHkZsgfmr5OUiVK94X4MYg2agkjFFKeaS015yv3UpMC
/zNt3kxcjqXUVJejDv9oPj3+ieS9/E7e+PuLi+01s7NO93gWJpnJ2UR0pSaEBDeKmrWY1q+t4EPb
dPE0ovqVrsgoZR3WNXlphecyQ6VfDW95a2UgYC2H+TXIynt1yON1Vs551/bG6faxKc7U9JlF69Ch
jtEedhwMZE0XVWhUquOyDiowo8GLcGytteVDhnoSGGKhKxfBV+O7G2P38cMN6JLd1L91JWL0Pzvm
2dJfMZdmXaSumga1jO/KFfZPUNBiaaN9OyPqmQY8Kg1jBMmRyxbES8P84D1RIIBx4J3f0qAayc+L
GLOOJvkDlHpLVTn2Rj9KIYO5pp4KdxX5I7jVmgKClDmAhhpBzlvCeFaM+fjZvp9cc30ojkE+II/W
Z4AvpzzndMSy698+Do/aJnBO1/7zvch/EhI14U9OOADmOk5CYHlPDbdtuNpKR+8uuxWZllqcxTyv
w4GJ89hA5LdARBmodUxQRU5F5m9wTzWCQB2UG68ZSdgWGYiY/TBCaBVnzV1Oi1gKz9rg7jpKSjoI
4/LpEoxYLZH6PfTYpF7GjCr7t7NMGu2n/Kdb/ffhVHdibiF661zf+WmMxv49dKavWobkaFXkMtFz
3lHT6EstJLtzDsk9vwtf7oL7dPD6/rT980HUFJCCMIibLX+exfB7kmWSkXI+APqcpUNSdQa2QdW1
TCGhPnDzpdzpJS21ef/c3Y3WGBpfEk3L6C8L5UDX3Afjzi3WVDW4bTDGlEXbXa34G9ajk0V/sXfZ
u/A5MyYtzUDimL56hUsucNA9PzfM6XkX9lwUJ0EtzyEFVWWA8v4tOf8ExlHysCpSDl1TrqVsiASC
dmhrlLjtziZeCEUOGSZEYbXRkY7Ndx9mU/e2YoRVPXuOciAh0nYbPeoMsMBqLhf9GaFlSFH+EPad
1iCSj1J4T3r/LwISbbJFxNie+/OlXM+K1SOaQ2lpHozt2nrvWfCBTrBwO4O6i67oo3hZuLL4xLR8
WxTyg3KOMwc/WufQP5UvzlGtCzTmuvPb32eBnw8K7oKBP4Cw1+ExGYxwlxbgxMO87qKF7gwkqJGn
zYxm1SzR5EW/gVpm17BQn5KOiz2FybYLDTwNhdKPhyzCdiZsfbS9VkeYTOsuA4hDCCx8iJ2QbBh5
WBJ5K2U48Cn8Fl7yj4CAFf/I39bY0dfB/Wc8hUe66I6YowOwOG0yWPNWarMF6I0oEm+J2H9zpS7K
SbcPQfvX9dsy7kAAi21dfufdUikZQA1/7DeKy4mBJsAm86uoRfFM2Zbqe+yPyAETR7nvGlJq0Mok
j9g6BcrC8KscGZnox/uqN9puEboUZWUgEI7VKd3aZuHmrT0iegkh+on3eRqthDjylCSfXEBEm2bu
rh6L4fXllhfmB23Q7jZPMnSGuMy9siHVBm03OjMw0XvMHyd7eNAFbPJEWT7pIDqgnZJFJrQWnOnF
obNOZ+tVaRnIAReuBRuOfCQ8eynfAoE1J5zXqdRMOdvlm0bVBdas2a4u/hwI+1MIDvfDukWKNmVN
Ejg+lGOmwbye8CiSbVWdGelpeZNNeej+w1hCGa5WFpqh9iawl7azR86HgfsSig9X8sdIVpmWQDgK
UUEHlmySy6iTOklotlI3qrJh2P95TDAoOfYClIJ3Evk+PNpyZKlLjoHbei60OQmEJ2w9IZxowq2e
WE/4kTVklAHM2o+DCodkJ6VVh4Hg35XwnPXCEv1whOU2a2+oacWVdITcW+ffNcgQ2lDyJOEygAWH
05LAZj/etdiO502nG0oPA5I91ZooXnuDwEV0nJJ6ipy31nZ8plTI3dVhbYVCBA0eE5IYHP1AiIQ8
HxX+VsnVxP4RqnvEGPsM20dD5C9ajwYeBLqsJdtCtlmvkEuw4PIpTXvjynTZscMuX63iwMzTZPj4
gthXAH/NhguO+FDX+YoxNDpWZ+X0RPUgFCAF+++UyGhbRcd3T4GHhQ8GCZMa50TJunqToQhJy228
XGdyzUY3Z+YT4IEItcyyCAYtTzcKq53x+qA4Riox8lyOGg8qa3Kob4NuMp39rYwkRyfJWZ9qKWEJ
LGa5TXCtaEYP9GVK5qSZVWIyDQ2u0b/PnJvZJ6r2HNox87LRZg2uZyaTURrakDlTBZ/MAUz4MMWR
OsoGYnew1ZV6ig2DOJjdhMpCEJ0XE4s7Z02/WnRX/C6Xyp20ckwp8uTOQe9+QGk5d/O0/GHEWDrx
ttKlrO+ecdW5lzYayZfPTsQz0A0VhuVKZKROx5VBNTTVySk/5BaXtflf35BZwMfbkpV6fMRylVq2
lVd2ZIAhm2OB6z8l6GIs/SnOUfyRkMYSmILLebWccUC7yLrYFxAA/2swV+FRqusqXymq1PxU3dLv
m99WZGiCZESU4CLSyohXftUvPwucwN2vOdl8CGiPvetx2sVO9Z3bxI3QHutXWoE/yrPNhC9j7L8v
McGtzBn/+TbrYNm9xzpjHxfJDaVx6m9vUsrmfjnQ1QncVycMmzQ+Nqwh+irv2dmHtS+N2Yj9HqdC
122ZL0zWcNyzfMaDSLY70L5uxmxJO532wEGH5BEV7jkweu/3YzVkUAp6cf3XFn9sqH2fzmYXF6+i
J2Hu0g/GGSLu+wdFOrYfoH4+aQdZTwIa+VKiyrwtFXLTGDvEXJhDnnMvq3IU7bFMWrRS+Xx26Xjg
6F7oo6XHvaHGZEwODE9BrEHJdCt6+BlkcCYV2lvwIFjXY8QqKSCuA3D+fSutKrKabGaQTSZ16W/b
TAUwdzL87iEF0vvHnOTHD4pzqtItiC4QTXOasiyMfxV6IR/MKIgJoynnflCWZujsIoURmkkuxNJ/
VqgNoySq3tak3yogIhu9qrpzJYwlmglOP+blVmclslo+QvKlgHvP0uPy4yP8CrioHYQv19iYnKDr
CkXIGKboHGl9vhMW3SfxNnBbwwACsN3C+0wqMPTarC/hJlwE2pAa9o5ooT6D/gWP4wdt1cWIPNLo
6/cPyjXKEkw906/UNhL9y/+3cNhha6CbGYixrTjJNfDd5zdggvhaKBFhDyDCLfKkrER4R5/+LL+6
AE66vG5DVEdfDujYzXGvVV2Av3gx3ZaVyMCOEsoXI82Bc5gInixNt2v2vXe6QtZGGa/UM4iUes3j
WU3myFMisByK4Dtiklz7TC55e4OySJZIDKmXL5cBZ3wUnYsQJR1P+sqXvhl3t+A0B7xc1P+WYkEM
+adXjC4Q0Q2mJBclV1QUl6upOTH/COppGGVhyjDj07ZzIXlLUIwaYVc5kz66tKTLBLFTVyKIXyxm
+TnDJTl3Up9+5gvBIf+uQUiw/llclOpgFGIVBUfZ3XFubLf5d3cawUvl22VE9Q22Js4qcg2bN/Gf
AXKZOJACNN44oSvfrdqSM7xKdSig97Q5rNFc8fpu+X07BzMKp3fd+6MPg6bNmDh4zrN3cL4pJxDj
DaxfWyLihfE8iIhLMGGB0NUOWZHmS9nLbz91GZ583VMM6Ztj3hcip59PSgkSvLZOCTAtQ35nE172
S+8R1iJvO4T/agaT/JRfAg0FsCx5vaoBfDcnWigz0VZCZV2wtchg3WqBOAQWV4dAosENFiKiLwBq
KhP9K7hKIxW13BFG82he5Ds42ILdO8k3mb/7Q/ynMdGabsTXzFbev6wR1ctcEVNIodQyFwHv6X5y
3jpFVd9Lw1kb3Dt7JH4+QiOBzFR/ZPpvrzHGYAkfIzMFY4cys5em42TmvWPKwPzbVp6JtOh4fJ5M
mRNLDQlNMYZaVh1A4j1RodkjGETKz8LNF1pR8KXoh+xwJhtjx8K1i6pzO2LOauaSDm/Y+F4hpvE+
xiG0WdsmbqvCuK/TMBeyn+L8BIsZv3P7OZciceXjHLROXVbIXks7TDmYHDYiJrNkkvhGOCofTFeU
zLi/3e8wd51ZRbE6PLKXgU+sw//xe89HFvjfIIqSF7Ye2/RgLfjkMZOxt3VxIdmM3QRSnUsx8bEF
MAGoWsoJEzAPnglF6XH+a1PID/IPYPr8rfJGXO/fIl4reMBSnlzynwb6End6Iz/dtd8FeykoNcOD
NZO7Dh3z9SAT2/a6U82dS6b42QSIzhRPaCXh3yNpIWWtn9+9D9f39D5POvG1aqTPbDXgeQjGJHow
BSSykqHtUvU0foK+MoNr8thir/4z+qNUgXEj6WAgUkQRs/gkdpWcQt6YkLSuSvfKHHuLE+VPThtV
AapDbycAXCG6Iy/AvoNoV09WzMobxAt6HRffwbdgn4LLCQcunNiPe4+PFKD+j2YW98ccXuikZw+n
TNr5wRHt7C/7+8JrtN6takYD6OCZ5mvdeb+ltAx8elWFD6AckdEzfu6z0cag5j1ts3AthqjVYD76
8TBOhx8L4TtjEen/RLcPpFRdtEyrCggpuU79YNyGlKrOZAeLC7rPOX1ncpYjNTG437eKyEjkW21O
AZxBaQXnMR5JiA8OdmrkAzJ1bYFvSHmW4FLpHgkjR7uLgM5RWtByTwELwpDzKRT0E39Y3luodTng
GzYS5A/voWJp1h1Op83WTjjjwb5L7DYj/gC66rSLhz0tZ/vUzt202rYcvLbRU1b82m/mn68WWPTw
ukjb11QQp92a7HfcCfylfFOuJT5svGhIPHR3rU3IQgnSyUC8jnSRlxoO4CumZ7q5u2vWlzlbX9fm
LcpC8zwIpD28aYXO8yp/GT07ouzQlnjpfIJelRQig3lwFaJGcK1gVQo0Blx8rv0qZkmyc6OXENQ0
uRrTh7fOX9jPN/gaEQ2WZwG+FTaC6wRIY7j2TLCuDeqIdzzXoPo8NhbXiB1CrzpccQPBGbTSfX1G
1YW+TFmvr1Q/W3j1dBadKrp6KwRkVqIao5gjQsVd4/LxQCQBrHdH7DR7y/1xK1Nj1iA7AzBTonSu
0Q92UFrIjP2F9hi2L6JV5aG//DhQOhdvRddymLpsi6odtZCcFVqefNUxcMwabfHrfmQ0ucrT4mEg
VDFGvUwws/rK6CqehVKV2fLnsHXRucZrEll3ehatZNeCu41e6XASKakNgBIBXcsqe4eRqMoJY7Bo
fXunZ+fI/E6OBb0jDy/dB3RdK2y19CUqh3wthNUkufYy7AcIoBRzJxOArF9/HVgL7wShKKzXYsBB
zMFDfn9UwnH/gzkQ15pNQJruYxpjmeGCTqckt5wQ9ZXxYmtU91r/dFrfxGu8dRwLGYSHqm+N4Zs4
NJ1HKD2P+KlZ8dvlWdy8Osgp0RvtL/HWZ0VZ0G3tC8HrQCJ7xNhhl81TQilOi6u21xO99rjP5dP8
LHZx0UvlV7xMJp7StLvNBbgTFDeWWXyIYV3wP1xC0eRkhB02xalNShSQfuqbC337oS5JEMZDMkIT
qx7TwoTNW6j7q72kaHBtCdC7k2tCt5JXj9BoQ3tgMMgpSw3PX4HEsBBgBONkc8XTXFg4fm0Y05vN
QkMh22bCRuQa/f8wh6hcVqsgQsQ+d0wSSD75sK1bUdjJTKIgkfNzZNEDf2v/FprhFXyhoVQa8RHe
CLAceF233qi1ETF/SOWaC/gnocstkCX3vdENr0XpowbFWNUegxvBLQdIiMQOLdEU8NazT5jWmQmF
lB8H8i9JkKvcZblecFg+vMwsSv7yxAW3tH0pOMg0BRzgF/H/Q47hroQjnmV8kIrLu7y+miMuRUt+
3GE+qZl8HQQj17FE+FfC42+Spo3mvkEJi9kjHI3h9DUTPgDxsskaxhpOCy9U9DmCF0J/PTOxhh1h
7BicztL5WQE57+nL2xaEV8BCzV+lIB1Lq8IyTrjlt5ysgZaYy4m2GRT0oO/16uNk1plfYH/dbX0v
AcgdAyR/5Z3g9SNSPXKl2DXB5m5lWjA9IlO4wG8pQj3sk2RJcqkAQVZEw2j4FhcLhhQnCIdwrKeh
aZqSsPftcnz3YHEzfIW6VVOcf7VgYzbT9LwJEKelKUiGZ4jio0AbOcCn4iSI3lAHd5lRvwcBF+2Q
xKmOZrg6cao5sYqEtCtl30mGDkOUj1L/COOXnRpI7nw/f4dxdanpbmuRCNvGceghiujEtZC+eU+5
zUV7wYJ4+s2yMTTInEbesh/UCWoPa8u/eNxdGvUv7AW30+8RSVBNIBqYkMh50g8hl6NvmMM0WhmW
hKSw+yN7OHLFZOgjSVv0AdzRVO3HwKlTDDejdObP3QsGqs2BiC3kARB7315gsXtS39NArSVAkupu
hfdEuMgwplekaMT6EXI6PzAV96PlTtosgPado1p6+TrtT0tybi9qaB01zv7WHAdzU+eUuV4G0aro
o8vdmEn34NJNrgsPV/FeB4JxjdfUYBd0VkfSqly94GTXnDgQiCDqBAvDBsufo+GrFy61m+/fs8mm
tfaxwLj4tTwm1uy6Uni6maV+pvdm9nT8Qx4dHNyrwvrFC8oRFMxuddnnOQpePyzQoUaf+GO2j9QC
IX2xcx8FXkfy/Lm4FL5J78h5sHXfuw9Kx7iZ83I9R3aSbgZCSo5wkEUjlxAbB4Hc5fte58VRgwTX
ALPXws/wRDNoK3v49nSq6U0WaUXrdtbMPYbc2rjPRayHpksXfO5PuMNNrQLj86z4xqlg4n7HY2q7
vnvLi50Mb94if000nh4BcfAUCaGZIZJ0VcRKae0Y5areXcotNnS+mt21KuH7U6Nho/6drPxH1uQB
1FrbTR6ozZOzBDv9PyVz7m9/9a0DcACK/HhUPsz+XcMsJEjuGk6YAEtf4dNf71GOc25w74FFaiAa
2Wbcq9fnjY6HVkI/ZPgkTy5fR7D3YhQXHZaIqgwZD6dAWzmcj0D3gvVgwHT541gJun4T8NRARUit
LWP0D+0XJQdUR5tffhn22//kHbZuNgWRS75FoodT2iirH2Fiadh9SOqdRkPGCdx8jNOIYf91XFxD
lasbxmbf0Y64c1IIwTumIx1P1UOwvbZTH4QQt80liREbtneAPyEeE7YMT2j9d0aexJ8Ye/Hc+mft
HN22yncQbEpqLzRubxfiLGkiVNSrPkM0roKhUcL6AI67KUbfX+N4WSWJuO+a+eVKzZJCSkSV/xpH
GwAC/lXCHVKJoXMRMWf3t4yQNQYcdO1JeXefFAprTs8ctOa4JP4gj/XG1dMLZG3aT76kn5FhUQcn
/saKqgam49dREUw0xFwL8t6gI1hAeDB5REk89ZnEOYjwIBPh4oEo1ou5J4aocVZ0i6mwDm8XZVnk
5P4s47hSOMPpnIbvcA9y83ozN1yoSWsaTlH8B1twlR18aZ1nbNN0BWUJtVzp65fwrJJAIyghy0o3
q0m7hRbiBBR5uIDO9jDMcZ5Rx1VJj2slnoZKrlJryUohEl81j27uYR4rdbbboONyU4kFl0pbcSha
Lwha/DErBNk/N1OQnRqD06lxUugcloMEA7eAi5JLnOWa96k2ZYXWwurbLPlw4piX53xgMhfI8WOl
CGG85gDPnIYMOKgC1SlxTgXpICz/M/EGLKL0BoB7Z16km008cqR6T/ecVei5DS2LUf2NwQk6rqCD
rk8TLqxtKtjULhhYc9htGgde8dzfTh4Fsj9xQaq9nWqJPgBmvJlYES9W2j9m/ZYdlxHJQhKwbf8a
JCzttwsYXzZXuw8JG5xdd6naRjweBNR90VAKDyRji5KmpNSY8fzRdaLjapfvhx90kV+8ImQ51v3K
dI3yIh6hi413zDeownBWTaynP3k+aLhxIHqYgamMeXazgsNACxvYYfnwW0NM6HEXoRVAdi9M3C0B
1W/r3wDEBsd6BQC0c4j0AFTUg9l5A/djcNZxOd+13AzUqEo4i/Wy2KttSLtpWyZK0prjiJxxfcGQ
uUEzZwbpYg2ck34+c0gP9Wsd1UKixDvR9by0i9ZzhBe0HO/IfhW3YTTu8PLNhN3HEiTsble2esba
U08nLfXL3T9WNque/CQUrb/gRRwqQPZSkt+zYAfjH+5MvNFDWhTD/KoA+8f689O5TllHsh8EKhVg
k5u2MCk6NtZ5+Bzfx/r4dfK1eQMPsMyG58cfMd68Q81qx48PJuGod8B+VBX8Q1FXnJCj+eTtBSLH
uUsKli2jfg/lakl/R/4Dp9XgnfCP9O85bJbjaJ0avvvIW9+QeRFtYv/m6k2mtaLONeOXSuX40N4/
VNvXn00T+L3PbUyOVB6RZIXzT0DlGCxMksH5n3DDPU9XOtigqbvyrEqwGc00F3dWMze1CApUPwmL
l1puivxalrr81ZHv034Qc45KAZlaGztrtKnb/mtYXcdB1rWjEczeBexIJbCoEoxTtl+Tw7+kL5bI
iTtnZqK7cqEiY+TixCAe9kxCvuvrlIuLcxv3pBZy2KkgKevlH6lDkMtVAOxwtb29FjECjJr9Qtyu
9aJo7Kyqn1/JTECYSreEMX67XGtXv8CzMOGkcfJ7KGEvY1FfULrVMFAMrAK88awoojLwxHkb51Lk
o46vPF7pjKxL7asl5omCtovZB/7F4fN91xa6HJbPd5xwYc/YyFMM7CfXDqyJLSH1l4zmHYa69eFF
Y1u01jZKWc/15tqD25h8/icaJSXJIGn6yTLJcz8zvmYXxQfHI7OfBkQSVgCo4U64p6TKdD8PLol4
Ameo+O0GQP33tpkR35S8mIIQIznk7V/odNYmlICyaTr9oRHpqnOTcrnsGb1sYEw+orRWHvQsU/lt
VrOjj3locpmC4CRdNxTFD+tHNBXNVDQm4ntCWpsWeHdtNShb8wxWXi1ZgXHjq+5aMpR22mv729XP
H9lZRB9qi6fc4MngpFTXzQm+0qLJ5HuaI9IA0vFOjXNV7jGQu3NjAmPOd3k6mDJBgyEAXN8yGrAC
LW39YcvUFEB324EWv9+rBk735NAPLYIm9oFBnPQyZejWKJ6IrQ5B5qP0PT5zYvfVQmke8W/RBQik
665hwJJyZBvLCDVrAhSQHSq0trx4+0IdXfZIhyvX94za23EJ0rRCr2URWCrodbMtNXqSimBtKzjd
M/54vYVvejXwtYYNfft2NHxsp9w5A0cb8GxFFabcOtCT1UabGLdZ0Gdo79lBceq3qR2NksNuB0YH
Cw3jbG9oSEV8XLLeuVlzNJMTvT3VY1ZGXad32PKLad3//fNKBjOcCMTiyLcMWTWcSFj6A+B99QZb
k33eAlpKfNJ2eKdIg4IZ7FfEdemF5tuzm7OZr7lLJVKwlp8jI7doS+QrK6p2uscFp9SZi8n8etf7
Em26t5eRH8iHzT6QK8zHhUPq9pRp3WTtNDWPlmZ9syK1Y/ks186A1IXltkUeZhP+2l1qxWUElTk/
rKWYZc7W4SIyX+WrBX7/w4RfPGiWChjez25EEZU4oQTUIT8YZmnEZuCosEmt6w/VBKBmEkO1mj1g
fXvoER/tYc1SM8HV3t5u1BiYRSrZc0h+2QHFeWxQaeosmMqxep9tytI1/nRBz5Ew9i5On/BPop7E
v4eoGcv5zqoO620Dkt8+B725LQk2LaAIMQY3fp4i6pzosQt3bUWrdWCTmfTdOeJ5sSqpwKGDdCdK
OLyNxGnvWXm4xbz4jLgZTidCHsB0lxarIF8+WzjqmGkwMXDHMPVT3vnoS5GA9IQcUxZYQdNF1Jwd
3MEI6xZhT3aKi1G2xOCk25a3S5v5qb8kNWIyXGl5BkXBfETdgRweXaxaqrFCle1VPBbmIKYOrgA/
bHLlJUdpoTWMor+T53H5VAnWMdr2/EzUbwF7hGHPbJVwLdWi3r3/FA3bi/PSg1tVH1BgT3/eB5Ek
ao+lMwBcn9nBZDmETkrgh7y8Ugx7CPIXh6fxStn++7Gsk1+oA4obPVz3V4NJPcalUZBGfgM7MGLr
1SAI3vH7zTAK20RD6I0GhZQFNLy6I/N6GhDK6MMfOO2zv8++WVI1X/j5eEtb5ekz0Ml2s3kW/VR5
RaPoYyygUCfpEijuun0M2xDgVFeATKRuDV7aMzB6F69gKtybPnUJn8ymyQsd8GGAHYiNZmleBop0
K6s3+z6enKSmtUL1CgfTPqI/MvIKooNAn2TC1dp88RcWr1SZaPXOPc5OW1P+S90Af7/0luS/wNtn
SXSwniRk1kNF/JOUIh/pGHP5LnBTNW9wb5VCKHfbA/oh68D6MeLSjJ+AwURULUYIFzYudhbW0BRz
TwvbQS20YwE2ZB0QpIdHnMlyP/hBbh1i81ApO4rPBq6H7by4QdVetBHSCvBCwmhddnGtLb34NcUp
1zOo3gRjNGF1yzyx3a0aCo4ZwRlPzgGur+fOxyo8lHxewf+BhdAKNyFug4tNhMuHD/hY9EVDFd8V
s8v7KYCIlsln7hDt2ZcgSIrvKzikCaWpTlH3TunwNACaZlOGxZcVlYyawOjpXYuIJlJMb+6CXNMt
bHz0BZfhLuLhExHcz126vSb4lvW4vdvP2Yz3JDAR/jB4CDIf3AJl2WgnNZpmI7PKX85RucId//Yd
QCNELX1Ht8a/qToYQT47h0J8kbPeX2KlWVYeBI1kA0uQbSi8aP47THieY9uw/w0afW5layIwo/5P
2Q3PL55ard70Y/ecCvKMnVPuzNvF0LoIbHls/B5kDj+C2O6BHuEmIhlNcbcKnw3LOV8wVMGetQH0
8P+9Gkih10iT+ruYEecxL6zMDY/dETYQXsZEzvrQg86L/93fvxR+QupEUN22TzrfNL5TeCnScvXd
Xfxds2a/HCvvPmvK5tmsnVG8m84HqhrxdXury9uRQfT4NOwf9qY6g5l8mfzKjc6S78qv+iAVzGEU
CI1TITaK1cBxNXHoaMYmi9TNo8+Pvq4t/1OXORlMY1HyO/bU3rJ3bFsVnfi1d48wqlQNrWgGer58
1VeT81HLQn2zZmB41CBBqf9b8TaEVJNaaNGgNo1lQLXLg150K1acgA2whXeLpStH2dnyNhKUVKV2
jeSZSOqiU4Fr3sF5aiDM7iJCJhuFT54l1SUv7i3j0Kd6yS+7ClBLHsEK8FPjOwoXFtSpObNOF7Qn
EaG/1ti5vzLQA7pE7VgPMCGPYYApI8VVU36OTX6PKojPTr2iKSC7utEmowxxdwNyoghYZ9zVNFIU
anUbefARjoIqnGr0xWQbqiG/BO3AgKL78Ky7nnBmhENG7gEO8pTcqoBQUEfGP1VpyAUMyKfMHa5Y
adFNVrLoKx3Yl9dapfAA199KckZYNtzVdYKzCOs51Z/Zw31ZauVc7OhFi9AyFxSP39KOX25sEJTt
mqvGUdlnGgZOQJgWWUaSE8fOwlmCQt/0b88VxUGMGxVPmV2sv7jTshOnqhVFFyN96rtbWeXfWNHO
Ch+dr/PspP8do6/1VSyR6NN/A19u420lSEn9NJZjMzcTip0jn7RY6DOCCRGpPUMq7oW4anHn65V/
EK25yQbq0ootEEi8XEv9sWDEBkDdkjccFcJOLD68VsUgausQS7YPqAomXbbnBfm8Lchmyx/iLCaK
4Sx0Xx0yGU0urBwsszRYlMGE9DwwnIpYxgnO/GVSzgzfaI2yIPQv/+hdIYLxplVvxaxwiGUVBSRz
AOv5LceTSAp32nLbcmi8z87ou16YHObvl9C18UM7WyTx5wQFb5sldwG41v9Bo3Wcj9UggrzatrLd
hYTt8hAOtoo8XHFUoZVaDRHW4YW78f2XrUU5+QB9fz+yzu+7SJtUgKDB37zkdCy/QrWVK1lcLvlX
rl7ii4s/uRlY6qX74oECDKSR4M0TdTf/3tmR1yOzfcbqM1ulhwFYWG5PV0uDqng7Ys7Iha9VT3QV
8zZCKPXaIl+vaZAiQnwp2rHCL5d2fw1qdAyOJCkOnzlMQ7dKP+sPViETli3QnrDn+35JaGTp8wV4
ia0PxcdKV5fLDRcQO83AshDQ2Wo81E4kWnhigcwPCQbmOm5ugiKUq4YMlpxIcMQY06qp2j4ffNtq
+qFm91GcKQOpzhUIaGSr3IR0CYTZ/BybPjehVvEx2vCgNCKdhZFgg9wwAa0bPNjBOnk3NQigC/1t
b+1/hC7Cv0fJTryZzQT1wb89/UxmV2lZDMHcosDIk7LsWXfR1hXwuki7CFkXfWPLbJGzPXL2iEbx
/cxZ1sxZ0+pws5+27/1dF4fMF4uU2tWWebrL42bmb+kLlGX8g6tO8nW+t3K+H+IdsjbNqtScWiSI
Jk/bp4drKTasFOE+tOW11fnsLN7t4mOF9qezd+v8u4rAJtUQ2pmVjhyiSAHE84FfvuBHzeYP1H5K
0+cJ0ATQfKFwomHxhuWTEQ8uSyaEW7we556uVmjkSWh16Q5g94U5WHaZD4pFTdPNhlSefqvTyQGJ
5XQoyGFmfNU0ZP2tPA8FouIBD7cUSbucIEzYzTgQlBInOD6tA8340p184ck8qHFYKSRQ7Gp0XPCg
d9HqoJbBpD2mrH6vuWLtFU299igbdL/Cc9oRBdJCmmP2BV4M6viSmwApxgs/SePAzIDCMcURZVoT
KvHDEnCks+SiB/zTe/JyFf5hk7JaoUkG4/MV2gOfVbvpAE+YAyle3HXVxFMlnD4D9fWUBhzHEfYX
oKG6Z1CtMrX3oI0BLoAfE1npIwX4mhpbA7d3/L+XXZFQgjJHuaonBVpQGkz1Aju0gMswYioJcpMb
1xZW4Ec/4feHbf/uybEhb/Rzk+9wG7CbXftL0/r5+Ljoj6MRRID2fqGRoQZ8nnw50EPexyEUJ4y6
9Bpi4hWksHUSnQ2GtJcYYDSEvCuCeP9RNCZEbtqf8MKsmA2AhipnZs5Vd3CpwwPzxQScpkRhzhsi
Ct9YXfSgf6jbJwVyYPkQlVhgZG1Zl3TFsGV00iouD8fR47qi+oNnstVdGLYno7mAFgQGLbWEL6R7
0GJkXpVqs4PA6rVMP3sw6kCnVHvpNgB5iYkjXNjUt/RwfHY53ntYqGQhvmSBJXaLU1g7FJuf1jAd
HhHgB67rUF4ba0KcUEVAHNjU9DSCmdxDqefga3S4k2HqLxid8w4WN8MJO5+jd6e35E1AmGAbV64v
VHYaYbggzzTRBIk+QL9y1wCtq2GPHZdNFdQjsGE1Uw5Blnv0dNObzZQbyKH4041OdTW0tyxIHumD
ImuKuFYRUVMORG29YUGoerd++uYmmbQGPebwea7BJdYB3eeF47mRY2j4t4eT1+RfRTRy7l8gz7dy
SLaAtmD6+UolbzbcbZNTlZJxHAW1/YQDxws1Jylbd1olgTFrskHTqkBjd0t9WZdPVwKzg3mG6CQj
ucaMahZVIajEXrjL/fhzKI1JCeZtYIvO77I1ooKeyLHFoBK4dTY5n1FbNt65ZH7vJQ0il+0Da7rJ
I9zCF76h6bEBesG018S8+0Gwk7ELwBjKTui7AhrPHWUt+QPoffHWsQYvp3YSOL3FfHn34Ya1ggoj
XIH6pGWTdW8wW0pXmj1vJSMMi9o9MVzYrA+X2CnPSijAq0FzbCruVBjDrtH6hIvK7nXfpmYU0QZR
CVQf/K7v6JocyrzduEeUZ6c/z5iRxATAIyXlRjtRk3PwF+Xndak4d7n5u5Y0ypSLzNHEyRljFfGF
qMbYSOohHvCaZdafAD0YgWa6qZAovEdY76WQq02wJbZdOGVjK0ubfkwIMJaw+VriQYPThj5yHz1t
oYsAY55QqO8ilp1XoZ5fv2EiAbPo6AGVl5BK1Otq3caLbLKgUVlCQniaR3ppeJq2wcGZpge2TMtc
4heRenpKLCPjGUQM2ktYwQV23l3qyG2O9rZack7OH9DuvPaOBprBdOIHgm3B78Snxiwlp8jOftWf
luXJhglezHL3dWQ2ZI8JnofBfkPH58kixhoMBzxW0XElcv899P8R4G2o5I7a/s9APHycPeQo55+C
3Rt72GiXd7Lr+56nBO8sHnIVTbsy3AieFiY+vJdlx5vzJixy9f/BLnJLAYsz47Jbnu8EEYZOmHRV
XEIycjz5gz/qLxm0bb+G1tKPNQI5lYVZ3N2l2nkHYlssMJ4i/gEDqPzUHkAB6/QMDCLdTlSB6ymC
3UujXrKcoKvgrHh0RaRWTEYvjquWJDo/0tHjTLQuOOm1q7ALzLNP+lyz81hp2hPacCI05FEi7JQ0
DHWQ6WBE8DspkF4YoTsQunoYU+IPtUWbTqlD8J1C6uaDejv470qVRKjOYskMM+jkrvnQ6NXfOdgt
PlpS5KEWMCBu5Q4BZCmzIfyRVrT/qgPCnPatJx1p/3lnzdxWpNOp7BUTHFcmxgjy7M6g+fAx0UF7
UAmLUQHzIUbf1VfJCZ9mzbxqHzhyDvQN7Lrs1poEJRA600kI4oXH++mPBi8F9iQng4Kr2Yp3KqUE
yohFnPa4Mmy19YqYlWqtr06zms/9OWQkGJ+d+2NDeQ0vZY8t1RlbHuuCl+mdPI0OmeQSWlx0TxkW
xGinFy+BcvJoviVqdIbtCZx944abLzpI2jyiSZ09+i9mSImuGbA6SB+G/fcAzRV29lHWi9qvvrj4
mCkaYCtxFllYI8INlZacHJlgGAEU+96oiTXY3zn38BXUSMnwDiB1fkDtAsoe6UlodLMEIccmbP9z
dluItyT1bG3jryQVzob8O9p39rS5suuzN10Y13e5VnnIJxg6ZX0vrEbOnqO8X2BC+quLk3Y55tuZ
Oz9eC/rKjn38KYQAbM56jfzYZZ1FH/HJfQf5Bs0/1rgMz1igRk8AcKaeEsvRmXbs0IgA28krxDEU
3C99ycN5/TDfEDmdxIolPWJHiCLdPwd0pwvmOO2qs38NNxikjbAMvR6TW7fCSEl4aMBg8ecOZGKm
59/R/cLBufRcYKJVWPeQYh/CygnrV+oqpLCzuNRqPFwy/vofiswfYJOqO9uJBCnlRLtwxLKsOmPP
Wu2FNz8TaZ9NFGBrPyrgEHYg//env/E+N8iiNC2epe+vAfqVnnP2b9SfyExg7w6ok7c0Q+lZzUId
Oyxhg1jYiaNJHSoWqccbDXs77wfla5kMsl1s03FUErFF2KXqUxu6CuPjLUOUaj4c2OuPesVQbfgH
0t/sMdULVe1VPeR3tc1co6/QJwn6EXauTvOpudwMWqkg9ZcB+ovxRbhVgjde84brrIAiyn8uewV1
hGAoFjxNTFGFHRRdialXOVeJrcZpvyLdTycZ2LIJBgr4iovRV7uz8hnnRAVQhiiqEhV9w30PubQY
v/F8NzcxTgFWsGehqFc4tHhJoEsjVlCtocYCVpLyIokDYZNd0CH/J7mpaPIVpzzAnI/c6WixiLZf
32VMjIR3PzSte1X+/sam2DjjqtDmp0GoT/vUrGe5AxLAhWwW80qEZIhWvaGLlD+7lXc0dK8XIgis
AVKEtKEZiJi1Ab6MrUUq2lc9FqctMPt/iAXj6MJkng/olQObC4g8YviyHB36lxHkybJ7oqW995IQ
hN3QgUNaaGK5l8wrAZu3WGpBrA2DNwBQap/W8HCEfeef2JFUbiN7HtOdUCps81+gMZiQQ8DogR66
SU0vSjSexxDiEwsEgGiuXMIAZyoIb3ee/G7xLffjtIwkyxyR8hx6cnAWmcWYPneNAHtRmEYmuW17
5xb0NjAczFzE25CHl4LWpUqrOdZbTjNPsEkoiiV3W2Z1F/gF3YXF53/hIw4dA1yDgTirMdSEuKRx
/DPXTOMpMvYdyK64QqMJpxYQ+trtWmqhkhEKqH5v5+sFSzlQZiSeyZIzo64WB73DV/SXoCDprRZ0
NT+BVnJkKWPIk69Q2oeFrk/UT5Os8odmPJ5yOxL2FPvRdfjrJDXG7DVU5uAJGTw+DfpDoKBmO07M
9BgyrG+plNs+dvQI94T4+DLi7S1L8NwaCt99i1Jx0CoHRrot1a4NrBZ0LkvlcRurJarkRBidGdfF
mKEIYa5AvgKN1NBogn8x8rzgs1l9IrAvHpRY8hyvMCXTKohKZPpwvQC0eXrqjIkL25vjp6Fvw4KS
savYevFPeGE2b2XLYoxTUsjutnQnj1VaPIA0iZjcZ7jh3ves9a/6sZ+gTEYuFZ+INWzd79mQNaGe
7je2lu8yS3AzKdr0MXobUZwsAJJpamnKybWNRac/fRAPl3WX1pGqSc/BqRZ+PgWd8TumUoj57Nob
KwQNovlCgyf9PJyRkXOReGDlusVGOkHHC52stoqe2Yi92iZ/j7coI4SrSWBChU00YEhu3gRn/vtz
tua+lX94xZI0LLexf7VyQbc04oJYFtxj911STlcaMmgK8Wjhm65MnEPKCR7s7ps1LOBCcMhH9xzz
22jJ8svi72KbOkeclXnKdF9Z+EbG0x0c3XuIApvo6mtBwdu3VkDNYoCppj1iIzUSJv16NlswQNDc
z6Y4gu8LV7qdby3V4Tn68RQvACnevZj88NNdLORm4YxbB1Wkoh+aCj2lMHjTCMzqqqZ2ebEf0GeA
I6JV09G1r2FPaSpj+ws4XCzwPpK3FeujEoySxDVqcKOkzYaCLPMr7i7jUpBwkVmc1bCzzRRwgvJG
s0SkVeFGVNYi23fDWD0kTQgISbKd9YCXgeU10YbGrSk1eWXM/FOtIrTB26MO8uEAo4ftuhuiMkF+
WstNQ4r95yRN2bOWdIp3zpl9rM+HSghU39ewEvJhSTh4/gqREjCtFIoKtivmPIJBgmAccY/1O7XZ
M6F0LS/Hree79RVSjTHke3Hqtvm/7Z4SPBe/Uxthmy41gAwthJMTxvg1Wpm+yw8rWoDwxUfk6xdi
hAOCJ/6jIHdCgGyG8AIi8FB0/YhjjRzpm++iMEDcptQKVoJvmh+pxtDyaDqslaAnV8SjxdgZb6wt
odhkFn7LT/q34hFcpU3jrYv55bZsSfKBh0cR+/Gca7oWUKYam8i6mY2apa6F1Lvnb+qsKX3v/A46
VctwhaCfovRh51dCVzFf0U/xKyJFw+K4yRkz1RaUuf/+DSMgC+D5mvgiYLPlOLjN3uYCfz/pPirO
XAUCVyMIDmb+AuSKvEnImNI1AoYnu+JQq9BneS4onLHzfvCoQMVXiQniyZIvt9gTukv2C4z5NOnd
b8w6Gh0clGACyog+NxGdmyI/75HDSPGuFBPCe85qDXVC3dWT5Fkx8KW+e16F0ADLdKVZICTP1tY4
DKTAwaegFYm5eOSydmGDuwIuUKLQji93Hd3a9QGIOGyYOkqsfUUN0CU1ViKuwYgj09rg98uxJ7+1
WhEqG/YRZ18JUtlAfTENDVnZD4AcusmSCXgARTWuzYxBPzNHv6qSGvYyJ6Bx7AM3YQR/YaBUs/oY
y/RBo1Jb0CD3Ra6v9pfOMZIBU6ZvoNI5tCwuDZcR3MSS+gabq0q2eyelsbp2KlkszAO3T2Y7lpUi
qtC0KzezSMC+tZDuQN4/bXPy4xVIZ5IaMxKnZDbkRN9cZSKHz2vmKJtOlbvH0ISCRzyrI9+BaRxz
2jqE5ywREw2nqmXrB3SXRQ2E4MKf9wOTaCCWKbqf9ZErfw2U5+t0/tePFoZWvJl70z75uqkkIBS1
gkDzLPP2odMuLefcp8i7Cx8TwPDKH/C/gNBJgeQaSoODzbOWHCvvS1xFwF40T/EKUhZ1TOkwWCmu
bZ1ohfKcHcQ9S+ySOI/m6kFh5qs9TE/SIUnAMpLgHTHogOE8G6zLHnU8so44z7eypjZcmBzCQNaB
t/JTwAYIS/P73yQTTpzuUnjbjpB33/Wd+KYDpsSI3X/MPyibKxdwZi1ixYv02dEkyOH1r6j1/cuv
BV8PUMcwQyyiEF9WEXS0HD/uRqfqpKSMMEAFrJ8b7ZVMYnj62vCNcw5L+sF4Si3xwQHnRq/HNkOL
f/NayhSPF8xYVpp0G9jgx/PqikSWTN/kNVl1MriB/+FrusmC3IbwT9zk4biyUic1DTh9Ar4qUirc
0xqC6VgFkAsydtkU3mpV7JgsDPY+gU1gf8Z0EK2V9D6uSp15f8B46Fqydygcm/2T2mwr+Qgpxslc
r5qw2KWP32LkJpq07nUB3wONaRN+k9GVjnt4QVIxLtd2d856I/A3IzRrEUL25Yc/RvoQMCuPFiMZ
rbBDQcq/0yTOHZ6JBOjY0LW1t1c9aSG/LpacuPGC4rNhOSw/0pIyAafKvjQSjWdfY23k3ly31MiX
KDCyKnL8zBj9Tdi3KNXQPlnSLwnGWCfTbJ7bGn3Y1ZAPyrSS1O3FUQk3bEh4zA7ypyLDCM5y+Epf
q1X4qJkgLl1grjld5UYY2nn05kp6bBYayRGRlo/cPxbkNVjak7Hqd6MuMUx6IIXac9JDmElHVrnx
k8169NxdUnt0P6z20/hGo9q8+1ga1t15RZayllaqT+xJBUqJ19aNZ2HstfHUcU2oo7faX/fWMzgj
qboC5ebx/MmPoc+vBQ13IrQZ6jO+l5Ed1D0vl9GdXBLnUw0jmn14aD0fcPO88bBnnCh160e298qD
d9Y5ervEXxa2o4X5yzEtijJOd0jjaFFP+RuxrBa2ugl5mirAGHGB2CM4k4zIxZdu8i9tGK3YZQHj
3LgX23Y2Ut+S9ttWedG/TANSF/9Bd0EeQYCo4dOB5jWaxE21PLHRassoqj4F6VJ7xw7TXe64e+oY
o+uHQ+EN9e2cXWgL9l5HaIfp1f2zb0nLgesFLQyx0cIs8NjUt+Nag2owAJtJy8uHjSO4oQgqOE5S
FTOY8zjuGn13gQR5u7dAj3koa2kj2bQvU9PN74Kh8m6iYjXcrneRvH88O8NWjEp8w7SOHfU+ptN+
YMrNrpCwulxx5nHvHML6skkRQjRxK+3jAo2Xc4SFYFCVPhFgld1orD500CTYLjSkq2f+u3H0MblW
gppwLkX3Imky925wtXxAAFG/ARXmzETr/Gktpzn902gBzM5OfWe+c2tEfzZ4vtZCumsQ4uxe31eZ
WtwMwjlziV7QIGJeEhCPxU6Ua/rjRF5+YywCJrcUwmLxSBfvDqtvy7vB5izuu2Ak5YEBJ7Nb6v6k
qYhcQuwU+ehyqQfq89tqZLmDR6mFCIIEuDJ7ttlmuc0gsX10QGJroG+IEJneXURkapC9FaXPahbW
BEdc9/7/T+BpxdgeK1Fupdt6qpHfp6zzc1FM9oUcxK8pza7UjKx1lCJX/Elv53koE2B69loVZRcL
IaB9+CdtYjtY+36RVGwYUQobWAAKop7iyk0v6oJErEBboMEeFpGq0aAjK5C+6PGu/OlRt2F+Q4xi
aT33f44w8FIWZtmnARF2yJKyHNDIGx/nSPkPL3vKuVY5dlAGKrf9qxYVLlB7ac7uxWfgW9tgmIBC
2tgylZEpV3L1U3Z/LMdhdbz/CLveQCdHB0zV4GMF3Jzc4qP574jeC1q9pxwvavzXlj25hLYBNGD5
wOUsSEQfl46P1TQG7QpqyKJyVCtxI6k4jnlW3NFr00GkcHK0MbSO2MuJuL6+HtdME5n6PaWqpsi5
mrbpRpx+vdJp0+WZdN+kIGD1+GdI/NPhpfo1pDrrPjGEOO1IZ4ZljnLQ+99HIH0Q9qXKposa0ZpU
7U2AEvcPnbAhBQno5qFYeTMwaAO549FI3xr3Zt5DIBSWBA7JaCJpPtcscj9+us8g4i0sLEnoE9uh
fWEtffD3djTrd8IoIaGrszxiWuj42gsOJ+zr7nS/rlqHy8pD9L97zWStwp/RKPFaFILB/a3/I91H
Etf4hzf+wQLR0E5AGAKeCVNKoNsBkURBpGwNpXdd6z/T1hdF1ZwtPi9zeQ7f+EdjPKimABpX+71l
tBLQzQLi1ahoj/ewQrglmzBAj1Rj4gzXuXVxitgUCsFCDF5umaI3APO5ISOAlgbddjxABHyDyT7d
SxujFYgGEXsLjalAKHNoPYGioNNzXDc+wjiV/WNmJY9gE4t6PQNsf9SToa3tFDFnfoHrbYvdTRW5
01uePu2FTuzkHE9EtqdeQVB64l9MoFiEyx7DheiPXR0qfrw3dpQ4jsKpP0Khgf5bkkHk5NyDxdIk
bxRLccMbLRsT4AYllf7B2LdQ+iA//hdHCTLSvTB1OqMIZmMcWuRD8j4VzSkGF9aIgm5c7i3p1VEv
9emCdluHFz3tBw/+rJ3B74qEWG7Ia8od8192uUZVA7ITf+NrdGflU9S6yqBHXJNhQj1dp9alNjnL
ULg/etrPranlT1JqTfE2b9GNWg3Qrgl6VX/rX9xOHnli7XbrCPKHZ1gwp6m/FcSpK7vD8RMpyPFF
2rJXbt44lXBso6GHzxvdJWDSa4JEKRSlKBo/CY8KlfX07nwzw++c19td58q0wZckcSSDpyLTPw3J
fiaI+ysVf7OZV8tDtfR9C0ft0Pb7ZI/qIXlJSfLZnm48vNcN8VK8h9tzWKIvXPxu+tuv7rTq18En
sZE762GUb+bj/yrPx40v0x9wftiHRFdcD9UHh4iuf8L3idqw0B67J8JqhMhshwFx9XHuEWkIJ2Xo
HBwE0n7UaXbQp4/K/O1tepk0l8V6X/AplC0Sh9bTBBV7yEYQ5yAQzjPS7lyFOMOu1J6E7vM5m+tz
Ef04eYctckpyQxYL/EINE2HVfpntBz5nhaRptgLhUrj3SXnaxE1cVGONCDXIul1QKXROTO8Q40S+
ofDu3QgYd1S07sGN0Q/IsimRkot8B+OYeujUGoeWU6utuN4wYsI1cfX9NLZtycPEfqffIc2YoDzn
V/RlwQNyx76coH0GKYZ2h2UyL0WvOaHWZv1JQFloRWau+skR2U6kfhGjk5s79Gmcn9TZSx+CIgC5
WpjbRvbhX15QTNNStmZMPyjLSNq7R8wGoyefZllMDKNVWbHITDODCGkYk5s7BuGhjOIk2gYfWMVC
6k+UyVF+0Dra4KQmDHmF0xHFdu1DwZgmlTpJ9pGQS9aPtxF2j6kx6BdPnXQG5qnakQO3rdFLDK7s
7yjJQ9iPPtLsmpLTXeJdjWCzDPmGa2aWN1zJJU9NT8TuB2H1oj705ZvvJagDZuYlKJ/LsBjNKV1+
CHxQjNNLpJ/6QDWNKkkdhZeTfBowK3YAUU31PON0Y/W2qEMbLwuXtCCh64RI3Cxe79cOH+BWGem+
3zGejZVHbxJ3uQg7EyN2YaGe4LGYEl9CLyG5d6TZHr34tyJvuqbrNpGlEJpMOXlX0oyj81Xqulg1
X+d3k1EvFUjNGNRUPzHPDM9r0Rz7So7c674NiOdjR4St5NlMxUqHDNcjqLtsYlzX5xjOmMLWvCjR
OFGDmbNonWPqcXLgD3SD52woFKp0y3r3qb/AlwFdl97rd5xUkm7mSPEG1fIOHcHUWbXRybhMkkZq
GxVCVV74kXTLhf6MtHR798yomcXB+tAjSSgCY4b+K7L4qnOcmhwR4Fek6UqfSffK3eWUxsvdQb4Q
pESapxh+Aj1GfsKz9BxLJcuPUOcCFvQ/MO5ummnBvYIIrCl+oNH6cM2C6XO6fwB5isVUUkOSNqq8
sqX8TbycAyo4ohJT5cHtHHKBdvdRcRrpb+Bafo0WBSrvBjZsr1EVcWEizhiEZBY8non8PtUCkjoQ
6n0H/k0AGqXkVGX5H/XhmYmEWxDgxKzc03RK8tlui9j63CYyEhQeBGfpSjVQpCqzSqQZnNeL7FyJ
S6x6E6OgPuiGgBaD44JBco2Ml7fIZcUXEuWuKjQuOBmxQe+dyBwJLD+WbfZJmNjqp75J6OiJ3g1V
5ulrhQMjOwwfG9ZL1Z6eEfsNNBOgMBvYGIPuvzxIuDZnTVXiidZy22s8HX+n/Mg3Fn1bVVmaelgS
DSmveg9/OoWR+g9/co3KPSi4URSUNfUR+FtK5xkPte3Oytcv0OhTDF+QUkxQdnJOER5BqLx4TfON
+eHmk86ek/q3kHZXtradmsqzmft4w+F5KBIUpFHHKMd3K/GZv0YDmT7vtF+C0mVlifBQ2dMih5Ov
TpmMJnZ+wVG2HZiBMPSz7Kg+S3lb/nnj3QRawA1Hw+vG+x16iGXQDAq3AByYVmVCrRTDtpEGkzqG
OkI7gf4TGFq92smCbzKKCZS31eQUrOQiE2Rqb/RmSepr29dikWCDOhAWdhd+MFrCD63cFGaXkwAS
MIrX+/FLMel+nPEW8UAiYRAaN4qm+61d62zELzv9jkAEDJwK7lhAUxbeNjquckfycQjHK4mcbqVM
zdvkHxvTWvbW7QCovIfhMGiKjbXF9y+xvBfnTdv89ilcUPc4E0yEqxKH+mrYGVbBXKEXndabAnzR
o6CrkQjQI5gavyD/J5KnBSKnG6E51zQ+mGhwXR8hErYgFQO1k0n2D17Cu7OVRws9YoA1CaQlS16R
Wd/v1wtYRkJEYSUCCqqfWgK19s4E9mhkrjubfRvw6ZVpdONf8YaYeN0pC3HusEK9lU0eUJo4Mf2A
tSbSPc530D3iR9kpWzW1VezntFe7MTQq+alZsf00Ec5WgcVLwiCGi6tsqqdFGmqx0eQxF7zRbL+K
nDJP8Gxx48x37JUutBaYTPTvkRC12AAPvVhH6v9az0HkizvdCPTOuxbR5pfx7HgIQRfGEnl53Qzz
JxjwYGWhfWoFB+C/VhcbtmNsk0g4omNr8NMnLrhuxzyDiqauqnPFyVk0cANSFI6qVrw+DrY6lhjI
q0cDBKw7XJ5byMobYe0iP31vmmeXuMbAZuC5c5/S3CczyVCctC8eOggZ7shwbFKS66tPe9tKk9pv
azTKtnNVRUnds63tXEzke8Vh+l19+EPTrH5/7iA0sJGJALmKNXkgf05KA7KVybJcjATfhUlaGR0Q
nazJyh1PDrZwHIdpii90B8HB5/vdKzeWzms9eZLEv6N5mtcOoE2Wt008ALoZUGqj02jZfqH+Id8X
8t1BLEmaFquZbYOMdWXxc/ktLJ5YkYa8sF5oRyiqpqMZo0M2PH2dSRHVbujWO1ThdzqzB817Dec8
DsQervZW6O8KXGudk5WXo7sXnXYAxdhGO2r+a4OPjfYucL9jXrhr740TDly4yo3aOZ/GzYW/ZyYN
PUPUgv7rr5HAyj+6uvXM1fyzKHGsA972kc4Ph8vp8gGfSTRtGiW/OrO/rV6dZTcNkJMfVvkSoEqh
W4Gp8wrEbEoZEW4+z9A4QIXmZLJQAsEzQBBThAz52P+wlL1RkEMBMbLdPeelNdCqwDA05A4ZfEjW
2Baolbm8lDko0WtMe+XOyVsGzOMppU6a/EP6at8oJKzLZzG7U+vsIqlQjSTkItBPBy6N/QKyYqU5
o06rInb7EWmHGNuOj0ftJYh1Lh0IjQwFQSqCvIlzPs+Y+EET6rr0Nt1l1Ah/tYQnLaoBaMjEAzho
+/8jbHKuMVjKM94FZbcqVsNPx76/E92nWT6Q5iyqeXtLBmAiwPKU2EY/36mrtS3S/NFTN3z9ZmNG
pmFbImhJjpWtvbHIjrlwzuvAfQhatAyYHblRjDe3qfCtK+KSWhLJkJGxu6shQPsdCrMhYDPAcjaV
o2k8xQl5Nb2Rcf6ybWHzyPKXoFRNY1QZ2IfOPFh4X10xwxI27qY3Tsb/bSn2SlEruJVu55j8YYPI
sNaSZMl+A9i+JnCeTrvN/n7/Z2BbSZ4qOPXtbVoSKfdObVPqBWxjEbObvxArWTcXzuzIrBSdDH6E
RMfh7sa1/PcaG+VhapM43j/jGVgpi1nSMaLF1+SA1ILYcfSsbw6lQ97quGxE6Cx+QK2wvnK8I7te
6JjppswsjZzoSZj1b6R8VPWN7qWiKnF2z0IvEWEJNu+GeQ970osRhOoiRS025dBRbN/hqpxaqxIP
MdsG8+E6TfjSYlpfnsa7V/zbV7o5XY7G9szdGGmHGAIwKkVKR7zywUuQvvBXVI+J/QchIVhk61+C
D/HygTtYcLBnWZgXm6F8ofrHUpGY+XtqzvGg39eH0t86/beDdvEcrtBeMWvmauyuKee+9xW/WxyD
OK1P3eZcJ20um6NXK+Dw5gadgoRLIkWHb19Zh31MibFn7S1IIqHrMhOtO4IgzWxKhqEyBsI5LfZh
qTkKQvc3JoD8KQKoc7cu9e+k4eujAVlHlO1dPQUp9P19R1B80ZkFb9AWLPQRH1RuS2N2UCR2J6pM
El1cHpUyXifbZlTrlWxYb7mj/wbT/IYCQuDZtDiozGYTQgDuvqY6pzyEnf323RnWqZQuoKvdIV1J
GoL2PfS2i/86gA1EImvyC0UKfLp8q4On5zaUaO3NjL797hydJ8ketsB92aj7S0u7gDqK8cRwuZLG
Z1UFeorqvfm8/CHNta9vmPt2gNK9sicg0lUKaa2HtDSq3qdqxuJjix896cgptvglK+HuBb+Zf4V8
ykC5nRjvLDoYiU4ZK4mCoEkduge+oX1wAiXl+5nV5zB38rkIcfyo2r7LInJIf7202WjZIh6cZxea
g2rQd9sLznqqLeige539nlxpuTztrxCROABXTIqF40sRFSn3hvXy0MYjJUpxEfxnTccMV76Qpuju
Zjgsh6+zTJofYVXiwhRgkClC+K8ofy6byzov7W94B4fsMyiZ+VJPU+haOq4HIjw7d0xP2lHdfU2W
LHtsXBLfNhI2t2tQoyqPOYFZ5LAK1HP+dRCXOzrOZgsPRzKGPf5LBSTgRKsIl8853fh4HdXwHa+/
fNIoQApwvmLJXZM+w6OJJxNNL5lIaFp3AtMFJXjHmT5OqSAYdbn2VZYmTusXRH32PSIXVRB5P3P4
+5YiCBRF3kfQvc94Ff68ZbK1K4RpRvbm6Y2PpwDy46TJob5E/nqjCIzYZKDAqOlusA1jP8vNophi
cGmQfJX5FtYg1X/4uIZhktLQm+t8IjYigXbswKq8b3GQJDeAqYWYRGKmFFrZVIuiuWNTFw9zaUmq
vlUbFJ7U6NwV27Y5axdjHOEmI4owc22D0Swxe8PwpdgmDOlaNvKKKB2uvrG2/WKeOqSePl6jVm43
6dB18kktNHk/yj1ceg+EOqK42XJbgpPEQsGji6GKTzqnQUz6RO7QahVjISUcKtT+p3bORD+8Y8X3
m3d8M50l0/WVxcmZcM1COQQXzxFqqZBaX0sh6tsl1viAyAcJySet5GqdFGc+a/XH/9EQntbb3ld5
Rl7lWDvkfuT1w5BzcpUh12j8p9PPExY/LSJR4DCEHaNt98M4EzOkMoIcLENSA4KLrignL9F8pbX5
tCD7SSoC6Mk91bKzJha3nD2ZKZdEzMMCGruHbtYrSONdTVL9baijqnmfgQS3kh80PnEUUP7XnzlD
BSd+u3tpvVsr0Dq82gpsUtjGms9QI3eG3xZulrXG7kouEuxLQdxh/8ZQwk8S9BKTqLaGZGQWpCx1
aIj42WSMMXlAJGeJ3O9sQkAEUSWhfiLN0/N0fZES7KFn5+pQUuR+A6tvUx3GlA3hbe316S8cfu6O
9slpwB5YJoFDLq4EtxGs3G3wra+OUXvoJ21gt9v2w6RpVsBYgZ5sGPvsJCuL9nH1YIY4XKHlDqLX
k6v3gMAY6h+hj6SaFxTqBVyEZLh/EK0nZvrWxo83EpNbBLPNddTBggvUvE0DwR6Hy29Z/OfzjHTg
efTStSQQK2511cB9uK7g+u0Cnye+VmRLA5ZJiMfOUhSHCHjsU2slE3Ib7SpL+RiPdzqhKgCTlRM/
XQo/JjUPl1TyT8RV2H7u+E6szoohcBWqJMYB11m9tubRiEC3S73eu1wRSqkhMD/8kqRCq5eAJUpc
I+qp9sv0lzx7O91w3cqUcy5Ctx+m/MqM8/n/6fXwpHXVvyCceRB+wowcdEy40dDRr9GoRN+ImfI0
LoM9Ek/bhswPP6ziLPX9Mzi33xDKxuRwjB7fmw8ZKQvtLFp0GeVsVTfzbImVKm31s95sIKJHjl92
nYGTSPhQ98F1DMPlrVtkfYCjIVNvTOhjwsvAk2BVgcFPks93uaoYuID0EPm6faIv0yRZ/q79SyuD
5Q8RzGnJ8SCPLpIls1pcrv0x9XDZdZk9SAAtPokp2o952DKqXDS1+GLkqFhq/5bFy/OSQaXNxv3j
eaPUlOyVNlzqfPzCiAaRBkkjZqS9lq5/NVQZCbXBEKRUZSZaDTbkfSLxdUNNlGXOji6jy0XT0tDX
J/iFr7xoC5ecbFlmX5d5pZLN12rliw1N2hYr0tSR0Wdkgk8Iq5uIxNBeJH7IuHxHLbtHwKyWEA4s
4+aIDIfycZzBslj0SodNX2cw8oPc3W/iNkUWlslF8LBT00CwgUMz/dwcGKOGuxYVw+BjndbOn+ZH
aPI6Epd5S3Sr1H3EObTBy2WuOxeRRvdI8TAw3IvipRlEnSpjU1RGQB+06lSPjOR4Ctgo1Sh8zWoD
CpJvbVJQFdokOv4h6wOnM5tgf5dL6rVDrLHtUXc9HQcPzmiv0pvvfdO3GvVr4Gr5eNX4xrH6ilq8
Y1OaoydkWKb+2Z4qqizscoLbFwcszw41UCA+QMv2wjrI7wJBZ7Pv16hQPiJLZYycP7QiKPPJjCnI
rUJzsJIGoqPGnuFxEa68yHhv87M5JHNYeCq2RaC9JID6+TLSU++Symmsr4cSf8YYoOa/Qh0jSD9R
kA6W4ieWdJl7QOiz6R55eVGqjcfsIz/hW3l4CzL7+qac+NZl5yD9PZw5pDnBYE4sNJfOhOIV71yZ
0BVFf6XUSHCrWam/ZxNicychkHmKnjTbvSUD3t1+jv636xgUjDprHXqKmGkk/1dcNvKxlZVT5lJE
gSXpzUVtUkG94qX65xbiYO3Z3N30IlUPliG8ZCoaQ4519BDhAUGms9/Yb8VKKSjqdQwp1Wazsy7Q
jAFY1OjpphvDKdROSvGcVx6T2dU4kzltJrFtDt97SG0KUAEckixH7DORE8lStOIUZF+Tz6Fz/POf
DaooiQC7GhpzJWeOCDwbI/vaz+w+9zEQE6fzqpXsufFvST0Vi99aLWJZKKtLLb+S1bSnG5QZhoAg
OYNjeCt0Utmef+wn+rFP/xyozAZq7GXvYHwRZQRZ4Gby96BWlvtHxblGXNOfhj1vfU1Lfm/E4ySo
wlkTbT36k/p7zN58qRc56bm29gxQ2OGTVO5ppZgiiz9IwyIpiNEmUEAxSbeXM7NZ3HhC4SlSiSod
SS8VH+3qov0gKrhHL3J1KEnTO2iFEqUM9mZbEo4JCrPitauor2jDbiRENsFrzNFH/J0KBYKPRGod
9r9684bk1nt8AF/0sliOpj5Ru4AUagiuZXq+yuTa9C0UGwzrcOzjVACkYSfV5yunzVCCOLOI3w8d
TTnG8W3mazdfKPY4uL4c/ko5fdsrmWnIrSqWOuii6P8qzlO9dWEQZg3UCB6d5WW4mGslpZ3A13+b
x4etbE1wwBQ8wLQGEYem50YuwMvAOVGLRkQMIUiKaiaI6eENauQC5oeAeITWa6YK+/OvAZdjXrUe
MYbYPkwyVBrf+97Bb3jzqHa8jxab+6j96XakIJOuYS/59hlmV7fB0S+Y2J0bC4Bu1ifM9O87sZ1y
mzaK9cf954gPEGZnYg0B45BUfSA7E4PykcXmEeFPOJ8n9+mUw4ExDteKZsMjnZ/KohLuhpVJYSFV
6Io5Vhq784ftt5vzPVROkwIac/Htz8iAFzzGskWdr2fEWvSBAc/sOpyge6laiZw/sukZQ4btCKsN
8Qxz1iOKEQA3SpOZDk+ezPu3UH80FGQjo7FGhDB8mgaZh3HWvpfk53qX9eYMIxRCXgwRp2wjvZLM
d45YLpJantuauZBmw2xLsekq3FOLACdW1hAvvaUPG3wehCSaMbUgh1jAP00iJIqzXR10CZfMZFpN
rzqJwX0qrH3n2L3sMlPXXNAkY8se8iq3mBNMTfBjNw3JjlPV/ddWqjZ+DtUVzvnOqOhhOtm+xmvs
qx6pUCphcBh2ZjWcitpL5n+cx48tyweAxTN4fKiW7YKMtWoqf6xD9DuAB3wJ96Kk4hmTg2kJ4d+P
MGdyzUl40yQZ/xu3gCaxMcdSJ1oJDQeyR6VNj7Pjev4VO3KCnYcyTGHOFvtSvgHNZfGApeKKahWj
nwnKqOab9QWztiYxlHQy+2XIuNUl2CAe86hH2gr14Xslyi2MWrRjUUxZVp2qF4kshIiVLTK+95Ok
w9aEKydPNGPKCfy6s9XgacFQuCfTd2cyY3XWt4GSGCvXM3RW4fIfZS8WJl7Coaypg60loFGVOr/d
9ypb4FYKHLEC8uuvLzUdXlsUgSQa5ONcnuDu+F9HZ55tbsQ/mHHK92DzmE5qVl/CnTyviHTsWHH0
84B+Q4tYET484GTbddQPdZV8GPtki8yhKinfVshwOMhISGRTfWGZAW3uiqWHPbloqE/yQUNdDsVI
/nmmxT8kQA1/vIqGSfxDBudaCf39I9mPKbG/Fs7+bsl4trx4MCfqVwpebDTuAvrmPVx7ixVgR4LI
qdg2UGi0o/f/BC+Pm9BxT1HsE4I2QS+Q70lF//MRvxx9RyNox7zBAmVq+10DuGbfz6gP4GXmZ3UP
OEWt7NqTRLoJ8prgcUg0rJ9BlwvjViBQ8X7uzUPw6EJMWCi+6jEHUEbZh9vs+8r3W04DuF0O1H0X
D3E8XbvHSWbsvvDb5QL0l/6xOuv6ALUZuqO5aPLtVk8U2q3joehOUlwH4TNObhCfrKgDX3i1xxDC
BwNblDlM88FtwpybshtjJdxAF6cblZ3x5HbYZKaItvw8InCvSzIrfY8uOZ6idsh2+nV8Jmehtrfj
0WwQZ80+AUAOSeAtHvCy/DDVyzNI3838FnDvod2ybyBWW5OFxDXxx7W+XuRpu6KmwipXNzA2v2qb
dqSbSBeoQRnKh0nA3HjcqYOLkfXHNB6/6ZzPoQetB7LLOrStzB0l6mNu/FN6FI0ks2nT+ZVmqkRS
uQm+/PYlRpsW78IwSpMVQJAtuMmfMYSQkoK2sRxSVbvhyeuEWK1ZdYyC3JYOtYwWtx2roV469i48
Ar1ki0Es2ftt5n3BOJQEM/exgvWILWJlcFbj1ZDSy+LdaV+2SLk2vUGBMvZvj0xTbOjBYdufD+bt
zd0pl0Wr5cHWmmBQVxKR3Guc1lREz4IJfvh9rgzx2pw/7X2MFE8W+OIbRScpDYvNPX7Vvyj8i+Ou
BJOfwE9WLo5eaaUuPgsY1foT0x5jq7RVh5D84UGmOiamb34iV415ec4pdX/NOpUZZ3stgsIVM/XU
8mdnzsTV+HpzG8DMXC01ph3ABd/Q23UyA6oNvN9/6qzWu6y7cwL50Bm/BiXqcCKVLq/jgd5dYT8T
QuDm/AlEyMMPcUbhFv7s8C6R5tbUSMkGXZuHJNsqav1AtIxZk0GIYgSSr1aWRp5mRdZ+vLx7n7gX
WttxVaRFI8dECyzX3goTNBp+bccNxoBBM7T/CVc6Yz2Cpqc9n+JMzYmcbCOgUUBFEbrozcIBFma0
WW0JJwgqWD82/Q4rU4PN6+CdHmbr2KZfXR/5FTL4COsde0+eTKuNj7HXWT+oNG4it569yWYdssWC
cE0z3x9YdoFGdp79sOw29JxdOcExj1eK10r6Lf/VDBM+XqUjjVZf5SMcUdPFvEC26JVY1EDXKBu1
8L6ZzD9c0KXs9Bqc2/Pps9Xoyjtdrdsu1GRNBXXCG+iVtRoWTRiYbfCErHNppc3JkvHBWC2avU+c
BpRoKHbpVRt8B5leyHuXYXEz4aiS681/1RCoO8Mo+qh/0WU+/d3k/O5mmmZrbELogkaKjy/nTQDx
WNMeLgGdyKR/KsOXDqN37hiOEDhCY6dvUjymR/T7hWx6xhZiXl08NC3DukKTrLzDEESGOkCKteRv
7bYC8eVsj0Mbx4pb/nrKr5E6izasqr5e8rf0YbzRvyWUoS67hinAIvUOqTeXluQU/k4o+JD/1iMB
K0Voe8YbEuGmqLSacmD1l4wipjNOETXbvks0BA1ItcKnDbkodYl+nujNMtmlTaDD3MAUkaQ+RaDK
nFjMJ04ycgR1gYHHWcW7NK8dpeVVAPkSXeAJ5+p6TgV+zAIBEtH9ID/3wn5APIXlxMZFasOK/q3A
TL8D+rQEaec0v9j1lb3Gtqv6OXwULxdJR0bbSLb6T0v8qba+SYh8+CyuSC98F6QqN2GN7biE2LmA
Ey0+/oE/oDHbYoYCdoM6IhYzU9Aa1ZF31TdXFX6nc2uU9Phlm67eegLnt61NnC3FAkdRuLnXMlLO
QfEeo10dzWKmBc/kxChQPtnQaIZq07WMaTo/LVss2LyvPyllaKgO8tn/si4/Vclm1JyGMwMsLwMq
R3+D5buGDdho0Tj1aOffq38kpo2XaccZ1mYCmEhpw9uL6spS+tGcODrjT4ZK+yD9auK039IODk/6
eLwOp9o9Mo2J2oXzJHfusaDIMo62WJoYKxtIV27o4ryJDNqy7UKz1eoQmgxChN1z7NwK3l3yBBWt
IWeDZDhog1xTv9XNSaLlDilhMXaisEAFOAa1Qq3Wzr/Rj7HsOfJUQrXq8ckygXW1OR95pz0G8Amp
3do7edKapOf/HznLlbKBNoRKdpRI2db7AuFvKzWCY3KWTMWZppBk09dnjBLspBPcCeI/ELl8QBij
hN0xv0Z898RXEtK+tZQAKnd+M0lVp0tumg+4oVnNr5ewJGYzPkptoi1D1VQ9gfbvtvxqmst3xNRI
xaEu+m119+138BlR+/PM5AKTKNucFeNOQ/QpFE4nsZMkARImbGfFuzoABcDP0j+yO6qgKZzmckbx
Nc6PV5wZ1IjFBosJFDc4rYiemYDuSlzdvOlI+qbQ/V12yrqwOx/CGthcxcHNpT1ysrE9KH6BSilf
nsHCGU7w0r4DhIsszK77XOVig6uOadp3tw5ZnzIuDxDrDz2RzS1R+kjwMpGK622qtHfZU8oTpq6y
NCKLu3msecZwQ19fMjTS7CaZFAcT+YyhsBdenuKEO8xtGIwy9svPEJ2E8AsqGDaUoJ/K64mg1VBl
ZN7+4dcc71wYy1us3xlNRZSzzgGnWrWi6D0cz8Yn55zrtljDHl6dowNqblGnzgtUCFus/S7938vu
QLc+cSVt0rcV6dlhHX7AGPwGYYZ/LDlzrQ/UmDzsdaB3OMd3TwMKdu07SnRKM/yDmQo5rB5wAWV8
mFacZa5iMZQveGTaLRL/5eWqL/JFtBP7LdFUBIgob6YbQn8WRuiPwWmg2+9xzV8IIwdfbJ8nEDYj
+0IafUyYARHllkPkHWdYsFpDRYnvFFE0zaoV8dLQY0dqhH5F5oi0VU65c2jssM3GPuRy0AeKGM21
XDe2w8gWokux0NbfbjKutEkd39N0meyqvdQOim8VI9zigy8Pigszae3Rp3E/f+VW+0v6/71fS9Zy
cflpbvfqox7YysnlNbokQ3lciH+IwZtZZPp8q1fYoIW44uCrgulGToNyPi4jxhXcOIJIgowH9kbU
Dapch04S8LVpWFV1Ly0f/9AWJ9W/X519JMNGba4FwUmJOBcZJ8PWaGxqnxi8p7rqxowYla01kJ1A
1JbOdRpHiv1UAgxl8DEPvJ2e1gni6hJBrG0lOFDWxzP0VGTcVPPzngcY3P01fRhmmUom/J/SUlMT
2JldfjLyIfeYeaMA6pbT0rHQq0HsNXhXivcj3WZpnR8yKt6Cdi3KGsxa0lbsrM4j0pBsyK3KIsgd
YfanY1Bbon1Wv8O200wxhupc1EJGiDnYcxFkfZuraLwhj9gJ16wACItrnwLohfwwLq7kEP27U2zq
IsZmXbQehV/0XWDj23bcVE0sP1+arJFbxBoNJ/dSogbuqrPQatU5Z+oHp/9XPbIJRl78sjXJUQMd
paP+GHNCixzobUNqDgfUJ5hzS+nb9djVxsMBlThtJ0MIZShSEodiiNoD9u6d71EvChe9axxg/GCC
OvVE8OjmfWJnoFJoIqOySPXRDxEf4eCrjQSxXG7ToL9SPw+HIOpC+Nf9tuLJpd09X6+hnNLVv6Pl
XRn28/9kQQq6R2Z0N1htnBV36VK2+9e6qv4gMdIf88OAHAwyTW6VLK8EcvdFcVxrK9bp98TQ9/7Q
eXtplbfrMpQHw6TPdbEoG7xvzCORjDlqPcvnZhZu4I4lAHPS6rwac15npjWO2gjvq6vnLEDj8YVN
Nl0pZ0znD9YKiWFlgf8x7EREGfL81zagVhVB2JWtDqAk7zCG5KdMHcPlszBCK2qEwFJAORvinAN5
bLAVNNqNXNVugzAyo+CpKxpnWbX8eGQRZk0OL08/VlZoCDoBHTAOYHhQX+hdzkWFxwS0q4ipBElg
eoJE3rZXTKTJd3TRja89dwUNSUPjFt02DLNRYyALGbMkDw61b/7BIarVepPBqsrGsqi5L4ATD1nH
d2CO1sCJFxvMHOcHwXyrPNvNGJk3VYXhcDKlskVSm8k0rGSKizR7trr14kbvddS6xH8mHQHat4WY
m8mGhJrTJY+llY9kgvRiatBd5+dan8eXW8HcgbKFjn2kvLQ24YWbUi1mx3/ri/3f0d64vPQwCj9l
EozLilixqQ0N+CJwQxfR7nD+CBiRftiK3eMZbPXZPt4+6qXpx2j4nrxSJr4pt0GJnmcr6K88oy0f
RPQmy1KVuq23gxjCoJhB2z4Yh3eGhyz2txpF5njD8il7Fzt8BchDM53KdzLUOKLk+GRmuAtFdi2z
MK4ZUF6xopaDzvYp+a3BnvZRVL9e0Co9n7ybMfneLpIt7kHmz+DuR4yCCeL5E7l5sJ6zP15toFHn
9ZqSqqqJKH3m+7X6P59qwtIWiF4AEMfvxupXV8ksKRNQ1puj6joRGM2A4lR8IWTLkfunx8h4YcY1
QvnyO1W9kPTYKaRiZAk/yWDLD3dwu8IsyrNEl3iIMkpZk8zNrBoDamJATD7EQL/4RqPULQM/WMx3
3ERVpuYBUW8kdgJbMQGsf33sOGCvK65BPoONq+XkJWFMa8TATbgbGor+69DJlMUYin1U/jVXPEA/
ZCB99lzTVZkZOQBzqyi0T8sMYvtoYezZ31qLO9nfJLEIDRyS4lITkDxpfevKoIK0DV4pLPA6/Khb
wJOBF8wMPLJRi+/5sZ5N4/Dxx4ZjAc3lU3JBMKCXAT5VFPuHsgJVijCtf+eP7Ki73pzx05KP4Ij4
JXup4Hjw674gQed0238/aFqHXVSHPh7QwhE76D3Hp7OwZ2ilQSriBVYv3kY6+mSDtptPD6Jyp9KP
5h31pGDNnTefPPCTwnvg7xAOC/u/Fn5cMfY6q3cZSzvOxrJcF2bW33yXtRkRBN+SdgZYM8iNqZGb
9Rm0F1XVbhIuPTk2rd9+05eEd4LU1S8qAjOAEnXk9jCOx9hRpf1ORJQxH0iLQ+raX7WmVquR7oHG
PftkBjmTFbkAuQDuFB1nrzztTozhUSwCyJh0LvXlGiKoKZuaV7vtFqineMwrDyFwcbvz7jDFIGLK
eNU7htWauImfFq8glgTOOtqAQ0H2HysC3jC5wnhe5FqidcpHJofCL4MfXrwjkFSvQpz+OuVqlv5/
mN+ovAJFxo9CFBrRuK5KolBv5I4Iyx/1GTuEjd+L3elWxc00QFjZokCaFVQaaeNMDQ1vH1HsBcL3
Hn21LZe39gWAAcOHYKZklJqBndpIds476b5G8tOm8iu26OK5Eqm1HlcKnRIdKa+ih3R2EXE5pJ7p
+pWSXATsnYlC/fwgQf+P76sIlW5wsduMdTUdOFNf4EACktYCRCIedNzJ0KOHX4K0M4fpcLHGZVbf
WrIhvTciikGaZYN6+nYgXKLAu1PNN69HtQhcmqXx4+LbSwQbnSZ2dYuT8RndpcTeY1jfUN49+poz
9Y5XnfZ904slsJwgyr1062nSAdHvvdabH0cHLkpzJmY/ZBR8oa31LpjtihbXr98bcF3rJ0jdaM3q
oTaguf790G8hMAZl0TsRCERJyNZhN8uYwI6b6vx4W89l2ztjI6cXPrhkR+S7kX8sNe4mv72TcP+s
RmzkizgkjRLg5HrSXUGpq4YF5kVfay0PlxLNvDQrnLHInl46q+bVok4k0llaRbRcIfeyforogWEC
oi1u5uKm++Xm5jQDl+rujDMpVd8hn+KzASyK198KzVGI5zOhnOlb2GB9PVRVj8GeYEwlYwQGx5a6
1iqhWh0vxIl2IFgBTfLOIH3OiZHnrfWZ3C0hF3VkOT0OT6oURPyeyRthNEXFyP1TBnMmFClK3Evi
QLk3f2uChOZQfY7RtAwW6R+KpbbuQCgnuEbZOAVIFGQtJSGs+ultMXnOF3idL3hLeBqwulbuFkWG
Qj0DnA1ei9E82XBuim/0s2u925WxrWwXB4CXUCw0bG6GlciyzwfARj1NSl5a61tp9e1b1N8dsWlN
ZUuIzzYgcxDckTtBdHb0A1QtjaLXZ2NWfLRTajtjHh9bRnkeL1g9+xTwRIsvdxU5q8QufXadkt+1
Sp1kfOfmRy9ij0iDigNznPl5JfXT0TCOw8oBtb0B09vof06iIoUtrPUwdE2+dYsJF+migGCWIUzL
tisFBphfnZhvzcIt9w9n4AfzdoAqrDARcbWkfODFw86EqGOPqgFqW+sejnqHItds9VQW8HNy09IS
gnuup973ebjR6kvdL2/sdAeM9ROo2eBi75RSbp+AW3+VFUhWbMO7ZuXOyc3L+uzqr3z0H7ijzAyf
OY90uVDGKcKGiRGg0Rm6AUxKzSgncRlfYTPGYUt44k108lzXMWXfOD3izO1n35E+hf/ExwTZBlIL
8eRLgLpdksl8WdeAtnMq4acLzbTCKh2u7WcWvAV3zvgnKcFtykuiTN/YneaI7MpTYXlS1zw7lN3Q
3TQV0DZ1wDP4h/FhQOEHWwTkyTJtsC/V5ByJ4NQ9eTr5lsk/i2M4ll16ggis9JmLcEi3v+2crF7Y
jbRxbiNFmKHkn4KJWKfL5uiLoPlo2ui9MZNVWla2IvE8fyyFiFzlZsg40ZZQoGNhlt1PIOglw1D3
ENOwV0YMJXbRfAVDoPQYzDVShgReWf0MVWChPDmmJo20kfkpd0LhQV97kXAIeA5rpwCzhZS9VpfX
NWLoij2SyFbI230FGN3cu0O5JE+RZQHGZuKKmnJc/55plirUxlJnN3n3t890sXwI89OQ4FgXvllK
hdrlxCW9+6kYz5yuH4SY2rEd+UH/DXodVK1eyQdxSczHtNAjwRntTY8JU921awuSoS77yvy9psH7
Zx+geUmNFOA7D3ww6INBCypfq85l7MqFQgyvoKl12L89Nbn9uw4NaYibaqaVGYTFEjIUSwUKFaCi
AD2dojna7iLxLBHUuXVdZNX517pTFUFTWWWc5Vw1x5/XWigw045aWFyLAA6dMPqh1vQJ4tYSNL+Y
bBk1Lmuwntom1H81MLIx+pYylWw0cJxILVyKFrTZJzXxGqtaluqWGGRCILMsUkOHXmD9F4ZhGUBR
sICNPTKuQOPdGTV5v/hPVs7qSM1JWDnn6fA++/F43XWbFUl9aCSm/+PDUW2kCi4gNyAQ7e8f9Ozz
NJ/YaoxJUNvc+0287tFzOCe6zTHKywYU4LKCj0rJq8RU3I5A1k8qAwADbtDQ3bKGt8ogFPlEjjoq
BULY6SB6t0dmDudcXXKOAqFIGvgl82IMB6v7sO9kI3aDJXnymlvxmxnneFBFh6aCVBVc6/LnQkqd
vORa9S02Ao2mbtCLm/RJ4S4xPf6Rxb4C2u3bUYSEZfA/U05Fg3yNzUbVFAl7aInVuPjWEBf+yqkh
ui7GACFSMyGSr5W4yJcBJqG3Bn2nGkL2zo8DWe/F1bQS2zN5qBu7qrLdDkizATVMPsApd86F3Tfn
Vw/jHBN//pKnnreg/FjyPs3xGEtuuLY5e8QyXpkmvHnZ+KdjWu05W1QXMT7mn7JUv6tTtpYqyj0s
ZNJklWR6kykGlF+uAPJJrUKjITA3hSJpY0b5h0cxt8n+MtlzIHfO4ugiZeKMe77vxXMfLvJt0wGB
KCig8FAzfSFAMDHiGOsbQqGejnk02ZmumHwVe3pM81yb+Xr3+fUxgm25wEp+ZHHdA9TzbQBiyApZ
hws0F9Wi6x7JnD80rPF4d+GNmRgfwtfzzcLKuVlJ2cWSZwCZTHHi0GppFPLUoOQ3JVO2yI22IZxZ
Sq7loLyoeP40dKulLKd0ozPo/aj7QDqdMOSrVT0XmYlbm90F+gTDt+zCz03rnnkbw0mPuYrND4hv
TrUo1W/ogkEPEUpc+KsCzRhzrXHXEUNUvN7n7pGWBgtHskPIu8b6vfJj8MCbW8mEuYzf0jS1nYku
N6FVH0B+ixr8Ot3+xTQK/w4R8r44LjYRgNht1Kjlo3p0xosB/xTAA5XXZdwbNARZMpadv/ZEEqNu
muHUxPO9xefqlcm5A54Z8yPIrBOyQxv5j0Fko5iI9C2typb8amLET+6d/5954VI9fVX4xY+FyAnc
HaPR9FUorcUAHxoTumgMx0bE2scr2Khr+tVZD4eluoQQghFSJa9Pm0NMVEUzBaWfubDiyaLPg+Q8
hktV9VrI/Ob0r2hYr6ZoK0fWvW0sf4B1nPpNjPHE1hJdLdXQ7z+OrUvfFatpqWufKrxCQ/tdmS3Y
Nf3iQgrXKzvHmI67yMVqwQht4d1/5LsgsgjRTGg7/AkYJYyt7o7Gl/IwZPNwYH7L/L9q8IIqyfKF
sG80Y2gBkM+k3Wu+s5u8EHGFHTjtqYX1qHu6ssqWxzYKgt0ifHCDU7WP3kIqCegLf5WPhOhktwIv
H8HZR+D3qOo1DvFPVQdxu9U9oAC2tGmTjBEDoTVlKd/HLHMNbuInqU4Dv0ypR8dPgLkJ1Ne/aFW4
fBpA+6oAau1X7QJ5XTP1JXHFj/kJsu/nN+z1Pk+kIv7B4EWWeVKVaw/ksi4t3iCIMLZsIsZhYDp6
o2vPvoH5Eq8Ye3copFWut88srLqlEwu1UEUBb3MaRXAw/ahrkOpuJxDRqBuAY9xCuy3zi2T0mpXq
fMBK4konJtB/dw9bieK7+LzH3Sp9wxO/thHBnR6GR0m0knGSqDlVwjDaiyYaKdPgeKsdG1sIGG30
3NkCxQOhWRTyVyD+TQOK/8aeF/bObbF8l+MK2ksNfEG3KqOQp4c/xRG0U7torbcppbE75xIA/qNu
6zyj9Zr9vpoHBo8MRK9/ZtMtmz1Qz5xpODyczb42U45ynhbRKRhySLnqIdFXdGYJkfhwhIq1lcnn
SXEEiebknGoJEvDkH2XJHKWoXyt4ZYJSA6+mbLKDefierRBXiErSm9kJ1Fd96TD4JNhrlMuQ3a8i
6jfODtvZsuHjgtjpEfPIZgklbDEQatr1/rjiDrRGr0QDYVGFmH3aaQhVPRGM4Hkrm5Brd8BmQ4yF
24rjHOQh/7DpTbri9BFKHMiPJd0INcGU1PARCj7WtFFAe3PqUEdRUtYk+K9B96IXLSL8qYjV+6MV
ro0jXWXTBkses9s2RyqRZ5++EL30ND93K/kEVuFDTR4wQDAbtCnV5eeM+lNu2ImDBIvllFX6Cw09
7Ka84Ze1oIbVQKwUpx1soJD9DxKQwF2Vk9SklGer1+An64fgNH0cjkz2InP1xv37dBljSvaQu7Kn
vlCZn2hhJuBv1zE6Vwe5IgJ4YhU6ZtHP53rdcYP5s22X30zu1bO16oftDiTDTZqCYMpuH+mWrwyn
FrB1ZI3Pk+Q2EjzJOm058+NPOWHZWaqSvnhxpPZDoWAI5rKLurDGpAzp+PayCCwC9zOnjpwV+DkM
32DuLhdcVVrkAR/mqTJzqqZsORTIjJL5R6XhDUG8MRt+zG53ows/9VZhKz5gegeMF2c0pP1y7Jvg
5Ql54gab7GO/BKNZkjNygaNyamKE29gi7WINbPkMpPSYJ6kHapm4nrYYNhIWrzwdu0txk3JAo3lX
H1RomZAQ1xhlTgtPcPH7xAfHKB5PruToNMGSpnuW1bzl4BZJR0kvRiSu1fVo+FwHmix18Qibmv65
EjiEzjPX9nXTCLOib3GnC1PJOYwe5/jMKkReSnzHWAsHnKtAnfFooXBeWZ7tKdz/z4XcvMHawC7p
ZpFi1C5JT9Wu09af2402Vl61S5NJinGu1iCv7OO6XBEfaW8UYVod9entQ08RT7ZgcFBiaANXp5At
uBHEcLD+Pnne7WyQOhGea3C/DFzWeKQ1uRe+xWxf18mr0rqPi2nCNDEjZpuG7nryyYSS2gS7X1E5
yLNWLz1w8zdU3UelPlG5URuC1Jp6O0JpSxASFwRgmZ39hCKVZ+2LCUk27cgFMisfjLNtrLdQGU4r
2VSEISf8lLWmyf9hg3/2IsHP2pDsFEuSvojGAFBvJQmSD8iJIXU4SobL2tXMAYqlJVQALd9uIG5O
5leiEOCqyL7n1UBJ9TkBsYgQRhtYhI4XCkVNtIorOkQ3uwetjPUUEK0JomGuFMzfbZ/gtABRVJbt
uBpXcIVBRKNw5bVSkxPyIb0ohBNrb0eOBqWOz4NzwQu8nVkc6gIFRH0AdWP42N6f5YWUiMUVWeTq
pBMGghTA1ALEmApE3mFU+sW8jRVKezbybfYNi/kC+dgePaU0ivfdGE9HXO3vZK9AfifJxX+A3otU
kkvw8O7jpStIU1CUgHrMwQ0wReQzaYPGYyQZVWdoN676pd3St8AAnqIR5gdgXiFfrLaE3+lBKuWi
4QpzwViy+4+Cvc9dKPy4qRrrjtfut8LiJViZerwo+Cs+RM8o/LjGHn+l/jSpBENmRFfKflBdtkrG
x/8Jp9r5OEdKVEeBomQ2EvfDvO3YS3QAzXToeq9QLk87YxGhZB781yC0oof+VIHPNtLO3JKFiwC0
iQsQS8TGy8SzCcEFI3TnLZPoRiVT5r2GCEXcRg8GJbjKg+N4iV1/SA4KTayp8R5TRSoK0BDY3oRP
a0QFyFer/5wCyyv52pMrsp//S5NRR96UVKyVeQxWnLv9FIgPUq/EDPiPLwQpcNjbsjWOZIET86BT
UVsDADfmMue9Xek1ieGVliQisT5LQnJQ5EP96VmPfAumNzm8RXscZ5cYVfZ3exo0n9TPpEs1JJB6
OSTkhY6Yx2SYROV4xGXdE1yZnFehQaBQhUVbJ5qyzt6lAm2puRtMsuwHiKGfcwRLsAkZ+Qgcftn4
0D6sH+EI7lM7owbXrhgF1IchImLcRIRg3wyWY+MvDOWI2iiHKsgeKyA7DuwomL6fan0bY94khTbd
1mU+CoVEnwCSImtfI3U4/vmo4g/24TsxDB3zAEscNIX6KyK/av/nTYd/lh/hyaC6B1OpmYnMrMax
bIrbx/x1QBQaeTkKtnxKym7ojg7rNrzRAOo1fwZ0Z/LdKuCR5TR+l2i53LHrCRx04JNPp/H/L00N
J2y7At+eCrK3jXETsX2UP8JCsfeoM8hmMWF2A2hWeeWD+rBOZ3znSycRM7R4NQI/3kAIW90A4QsM
7RM5VxOgF/fVG2bhuKgw3fxMzq2hdpkyzTap/W22GzBk10JIQNwuBCm7Kb/RyjxRWrg07u4Vg7wa
Ds7gJlSiPsmfnfRekFbR7M3JbI+4q5m+oZo1CU45j1ErlX8mkm3O/AQqo0YsA3vnRP1mkJRONCSy
tTIgep262v0kmm99hY6v8DraGY7J5fn5l2yILL7EMDRq6Tb/rwAO1pge1FgtStH31tBqaam+Kagf
B3W+MHnIpJM9FoaZlVj7FgPdEQfb2DxoQGO5M53GLcS6tFSZUayzbrntRKTSMUxlNM8H5pN25rhu
GRpZMc42mkKVpdf9K0UtoCWng065AoE4aXtYBbQ3nKe+QOwO06Y6nhDFZnPtfGBeXLCPw4RXlfGj
Vc6nszYcPKM+PVjbK/q/7IzUlG2OsGs61EJz2UZ2rlYB9JXDMQJgzTM6fAz+7mFefRMizsLxbUkZ
VSWCAONKEGfuMbKRQ1L7hwMyi7XAagmNxLYI0INt+0xXkFVmqrjuP2tkajkb0WtXUbXAKK8IyhJN
XVLMxrwhQxPbiIcHOHCTOR3EV/0THvfHUtv7GcxVQA+RzSz53/KBDk/7V0bcVpVlhUYnSkqv2Qxp
Wt27ppJP9EcyobezBaLspOw+/ylMkFl6mNUlDmyl7lw97EFByLAqVsJIanpgPZ+/XPzGqueBvRXg
7eRMzy1YOqW8IOcAGgechFG9XSH7/eJ4j0HbcQt/hW6JAdSjWLLXqrDeNTsAlYy2J4wU1R0fcdov
Fo0zyU1HJ1uvulAh93AhYxNxuFzsbmFdxM6oJZZj4EAU28Xqvjsy3HBepsCTTMv7JyGcYjjEtoug
4bFgvG1jv8NbomWqgsYdISp5862FF4UP7d9MH+jMQOJZ+Uh+UyB55ZgXpsIKbD3vEbPPJWCJp07M
/wokp2Nz0ArTJJuTVBsltkbdzWyjeq4NewaEo2gerZV9JMlOWsm+81yzmTcSpJ9bfdmW1xCSDKh6
dHzzl+HPDRTDi8HeheLL++zNhzC6dbM2PsB5mzRAwX6g4as4DZRz2uyOCr0dhnb4NJ9/UKSK2JqO
dNR2ewe4vp7do60ML1qQ82kwLFrsaT0kHtusLrdTVYP/QHoCWMhJnvjHdSKjMKMjIdXfsY7hTsZ9
wOcI+svp2bpLp3lvKx6qiPRydDE2RyRwQuBWEg5stv167vOVA20B72/fWOJW8JgCkt8ZSx9gclG6
x6nclNHK23IUqSkQGm870Rc7TjqchUTjzRJ4fAJ9PhA6cOJYYa3XGw4swPTmtVIgcx6ZSa4C8b6V
85Bkej99HPzTUKsxyYiL2Lkg+TZWpFKCunQaFUaa/hRl3qFSAqcGo6RLAOiNAeKGGJNvMGP0QJJZ
PeRAHS/AlcrA00FEEE0+b5x80u9etRRg0AfJKOxPQARuh3wjRIcwiJ8QH6ZdautYOyu/9SCYzGlg
i+hoL3gU93vot+MVvQUKev0UGCC8t/oedI6WW7H2xo91OUancchCU2KVPZV24KJ2lhESwHdCLJUT
RaHb85ALxBEN7l/KSchdnEIW4ebOsdFY88kO0GsaxFNQ6GYure0tX1rRaij9HjeFWMJURKgsCc/P
22ezVykXyQBHJr6AsItfI+ir7UuuqCNy4z+G52HAIk+5QtTjU/iyaxdzXvOaYyIrteHsrEVNB9yQ
XcjvYkZZ2LaL9B0dSRsU3FiKyx7thfb9lK5OfYMuAXPzJAFMhcvHWKmCpWnTziTbtUk6xZ8KSveE
n8DqIDMbv6vo23OdtvIq8m9mxyBviWp1aZXu1tkVAo6gvtsWVFxbZWbD9lmKYUrmFEVgMcO/FyPI
Sin+Bvm1wPjI/gBsa0XqzU5SL7FSPl31xdzleH0p7RMbZxL6g5XYcFSx2cUpinC2UFps8O/DNrp4
A5JJ1S5HNT9wdYtzsi1dCPZYLtIwTG/FfKhBxk+7aUEHYJ2LxBMiI74EvAXjqIX9rBUPe1EL/u/1
W4pST6Mi6nnwLsMF2zAbajtcKZfNAfsLoFxCOI4+p40eR3gZQEvjMxEdDWVAfqfXt1EirC2RPQfI
PziDSIhcRCa2G3zxJazCwzgNwDeJG/MQm/pg9gR5Lz2vkPUM8sOfBJt+NMiyU25ck7EgXMbOjTJv
2opwO33QSISbsczEeZmOMHHZdtSs51nLhh43Ckl8Zh4SBhsU8jPN3dNYGh02fV8Qsuj0FFEc540W
O7I1Cl0KUD5FjHZxeWqCHf6zFQi1/mupI1o0QrsShQ8ydGw4gIKv499ABw+gObkrUp4FfCoF8MKP
LXROrq9FURR27RG3v7Jy7WO5X/QD25NQV6Z7c77mxrZn5KeXRBDgm0Ls1UqdwgksNT9yg/sYxFAO
cGnvXkGblt1KMOwW+281kp9CPPfK6zqn2D6eDjn84pfquucGYwH5ny+X/wyHFGMg2KHVB16i6t9h
zY2/5x1mFNB+99rSd+pEIipo3qRzDkOoUPgXnwxBLfOxYjUuFlIROfzgpbdx+2v7C7ozoYR+VLhk
xQPRUX8/w+smfMmMT5j5XHuOlVb5uiXeAbL+hQCv+l0/kFZ5VHdiJzsM+TKUNlrUjMeDNuGeVeXK
7fO/9v7cDkhkUYuVNxa40/5gTB+gmNqouqEivpxuIsJooTz54IGKumtwOkpk8oXaUvfJv6hA4yMg
CuaxSLtPMU48LjZNPzN9LDcAmqkh+SbyFg2rxb3nSghRLpSeETouV/2fQIzCwAuDfmkv4qziCuiN
rJpG2hnWensHTzIGsYWYEG/Hw0nciwRpmip3hFtDDv0tAY5rw4BlOdwZUxMg8o0VPPQI0kycAPTA
Tmf5IAu7xGsy93akIkDSgCOrBmK88JfujGfJWWFK374NaHcUGmebE+VBzn5JSyfN+EQ7a1Y/bOSc
tUywgMHVi8LhsxtUAgJELZgbjXLw8ZwH1xmg3ru/4CyCu6sKZqtSPvOcYd1lt89ex7oTPpS0ODS2
D7Z1JUJ8vJKsxiy+Y8ugmG843yLx1iF4OwxgEEikiYEBTu/tCNFX3EOb1sC9MuCWf658EAtadjaH
xEUhWc6ahPoOTXcoxLtXNo92y2p+YosnI77GfDjC8QP7ld+Hfpmh+Wb/xEQAFWUNb1l0doa/iIZE
aPfNEJs3TzusM5r/e04hOLCs2gQ4hI8a8VExmh9fJMSV6NRELzo7R6VE9RFV3ouXegbLg40CYPL/
DxTEMp7NCcOTk+KnId91XjmFkY4kP0QzbXhzp7E3bts1iJfOsPLzm803bgmWOd25VPXmrlfRj3xe
qsyTfwnIOAI5fcAehCJKLfAMvUU68nUr/7G60127ivGoHFKOp2GeOPAUGB0YBbeAp9Px+9jEbdwC
p3sOukLgOro76kjlbb34tw3MJY6qIltruKyg4qycPF4zQzue4/Mx2/eVi7szuqhCf4wq+W9GYA8s
RNn3jzxQtJR/B0LHPp7N2UH3tkXNR7+QChMQeK/M0aIdxNlcIIJ8XHeq6NCp2G0iRYY1k8wCMBlk
gHEsZpPIjvBPnKcUfPQ7Ti96FS67io1AsRLbbQKjvJYJh0AdvaZukLP1Cvk/syVoKwlC6RN6hN6W
+8NSmVYbC4GzuKkabQ+zZXJzl6KXHmszYd9WghFxd3mLL3WUqzNHbtO+n7qxo7X2nuovqN/zSq+Z
brZtGnD+un3TwhXfGN61mKKCmNRdWN2Su/xtAj5PlFCbOB/de2UYKXirsiRT6vGKIHXn6yL9TOBY
yRt+wlyMiiuxZrHoPV8Mcjlnc0NvJondGBEHpnMpRG/4eG8GprKGiU98SmbBmkUcpl9zxpGczzIW
Jg84z/TyVgvhWrrtHGRX/RyHWMJK3hRJkRFYY0RXdY1TUpii0QqyNKi9OZlQvFNVQljMS+onJ9NP
5sNupIGG0DPczxSBmXujg/1za9j+/gqSaGgfN/KzCia8DTUYaHMSOuCfaez5ax+W8/Zti34YXPKf
5fhDufiYA5N2jcppNzyXbpZp6w77+Yc7lVWFUt/gOrXqvFEep+yt6y00iQ/dMJ5c849+cqWAK7PR
sr4jOTCb4KVSp1cHI4o3opZwfkz8h2Z7V7dmCVpzEWocawsWrx8R7giA6wqhNeHN1UryozTuGY0G
vzvb/T6+tJj0BxD6zADxna9S7MHcJzlrQQzA7AhZrpcnKRXun6sEa8CePwSbYPONpYgxEDCq1Tjo
nMKGJrCnLQEsXED3m7l+OVmGJkcF4oCIpu6EcAJytFxJO44fC9T6cqXqkSSFCxdGPAJez6S12XQx
wEP1WpDmv4SlMvAv2Bpz+6HmNAqMZWJoq0qsjN0Ilxr2dNA1pki1IYdMki0nFnly6WZKa1Q3Q46S
20ypOVuSJ5PBlM5a4kntIuuBqLvCz4+6KZgNJyxMpJJHlZA2Yc/DIrEWO6d3ksxC8+F6w71u1AGw
gmMPWH+0srU0ERvVsvsMZx1LKoynKheNDb+Q/INgSFVw+TlLtF0Df6303dk/pTHymYT93U8qCkUj
eGK2zSCo1Pgf9EwtjnO4snalE2SElbn8zYCyNBSAInlLbJ334D0kDEcTfalOdttJ2d5wYatMM/6w
A457TZnqHRKONn7UJcG1vXP9V8rED/uV02rvgwpnK1Y2tE0oIazLExV2OMdFi92y70xSsryuYBzi
hCdL/6vOYIvo3ZUzeshH9hLByBs3z9fRb2ZqF2xvOHyj0bxhbb+cEKaMkmc9Y5LHOiBTMhiXvN8V
WGZTDgkg4C1Dv7iSenKN5wLJpD3G1jA/cexhegkZw9ll2g+7ExnsBaHzboz0Z+QbxrxO60ksAsC8
pc3pQThQDosciTEGqkzt92JUq6BgFt5p0xn9SqH95CwsDCFeFAiXtRsnwq6l7EZ+zgMpTTBwGRlE
DFFzPQQ7IkKJIGLiWiMMwnfiygv2JHOngqBIDM3NqrsNl3aV4F8itEnLWxmlK51gMjmW+hgsljQa
wK0YTaBdRj9AfkOQ7gvCC1EKT3+VHzOadPsP9M9xYlXBLMeJXjwbwA0o0iDj+u17Nw9/KpoCVjpx
0DzBjdbE15e8EQtBj+fQ9tUMsVf2pvubBN9VDsyKYenjU7WWaxxT18LpKjFLTMLRaKgsc8BUVDsN
rIrVjOiUrCDP4iFbQVS33+YSdFlI1abpckagQ1ythi/3BqY/s0FX3nIOp/+6EJ4uY7XM6MfwXg/C
vy7t+n1lWO00FPdU9qdpQYy4xIkS4mmJUVRnXHqyrogvKyQhJjTQ5qFgZu/iAe69oSJehUU1DozM
xFR+SPzcbbuWY/BhhM8CdUHZ/zJZHu8Qej8F6K9mtQYfe5pKSI7l4nKMC0tyg6UGknLNHhsrUYoO
sBw/yAm0j2kPF+TaoysVHB+8AK/0lSvfeXsCfkQLHbrTy/3T0wi7ooZnna9P6BmWsVK1lDuWqyoh
EuaCHBfKtL+LnE/KZJdxta8SOuibpCs55fb2MfllrWm8YE70r8fpz5mwz3HMXbeGnC5gRWTd9KFY
JucmXQIzHoAY3tv5b4j427sKeKjzaoyqhUu72cy+MbPcOY/N3FkY4fWdEtZJUYUGFglNNU+41wp4
FsCDgLNTQ52gQIlnyZ7wu4HF/9yBbweMtB9RWVdmwD1omVBZo1+tn/HZZggG2u0AND1MuIXD2qed
A3IVQipz+QcrnH9k96Jd337Tybd5Ird+2SvPiXaqDOb63WIEVlVJ45nya5nNq/oyaIz668+hsZLr
L7EmADGJOom3f9SwpQWrNeVki2fFZbf+aqbVUV7Iy60kFV6ghmyGH8QaJP7yM7CvedAJgEQBOXuM
KOlnEq1p8eK4NnxrF1X2ncjEFmJVKMceVyEUrn/UvaSUa7sMwGtEe77yTWM72WyDozpIJGzu/b6b
IcVAf5kUe4LZ1+ktvKknxGZSU8kbgtZgbbSOGLZwdUYKtwTR2V+k9slsVBv8BRwhUNqVQOU2/No2
0FcvJSPWt9BrsHiKCqhGTHbv5Q+5XehU2W7fli0ZlONu8O5G6cUNKUmKM104K4lNJPx5cxlq3q0G
NW5DmGBIdJsUtd5Vhi6emMHhfJwE1HpbN6g/KQsO2ugt/bn6AwqvRN9Xnrk8rrRSC8AeHGKvfxdx
ShaNX+3fIPxICHS3txoQkOWgJ0WpW8aA2jvPj05n5pGJIjmyirSx5bmiFGEEfBaytm9ad0MABp4r
147BkxC5AwVzRm4z0P1KSeWf1hZy8W1BfhBCft9W7POdhmkww5dJv6HeOI8lUIgAbbymjVZYpD8D
M3GVfIEwOQRSO2x+G5j0EYFIMFT/Cf8sal5lEVtWJXNm/FsWW2UYFJptoE09286ljHN+acl69b4f
1k8uyBJKaprKehhm2SUGLtFjySN2JSkWXKjrDyKhtAI2MAGwqv3Dvtegst8BMTUPWUH4myTz6+Ny
3cXKPzDKgyFyjT1ZDAKHSzCaNem57lZxwejCHZssrX4kK5iscSBZVhm6W7iNY8Dx2b5Uh6SLByHo
EoRhbGMzqX+c0bQLzK9oShWOghanms4Q2QQeeRf67A1/tdguskHnp9i92/cE7RwLIuQmfCiDBGut
wIwEF8jyZEz+rbg++tJhX13wMNZLYWAQmI9/5MlqfWBlzp9oop7xK7g0QwCQXz9mhZmuwfS91FjE
eW6vpujjpBXMd5S3m089kTx3J9H2eEwJj5sRQKSNjFihHbciwhwUtbCuDiFqfpyFG0ZGQwYRJt+Z
x5KF7BOa9HrGWdzHjsRerZZFaV7YX6Uvndtgsx0CPiCiP/W3EZY/iE3RLn6IIIjutGt4EwXyoiLD
p84qPA1ecUWN7K3bR15RotP6wQc8qrzM6Njfr41VEYH2PoJrzeKa36aNgNs59RdzBK89v/vQcrXs
HfzoYW0dchaw4gr31XxQhzRnhIv6AO8CNAF7uyMHuT+LUVM7HCkT19GSQEi0M7xq3wtWD7k7SaG3
6t7d6L9ZwRKgsfROj8BnhAayPvvuN0W/MBfPaYBhyjkGsLtpkhkRQ1LvNNjYJmP+yUP+UhkhZ15S
Q2zmv8P1jTVNEgEM5g3+4gcp4ZAKzpDLipsA3ewgdeAcRMW/XIQT6X6l4w33bWQ8lc+pfXM/kFK4
977f4AHfgOFV93x2UiH+3T5fWRMEcOIXfvH/qjHyNDSomMpQLhnQJB8qg3+8/bzf+304agcbPb4A
cnn/7Y9NxGnGxZib5lzR0ZuUyPuGL6z9hiGQx1KbdERKxuvK3oN+96mrvegtK9U9Ug6w/yESVywn
fNQJwXJs/0GQ1peAyb1BxTuFwKU52WTwgDg0blaf+ePOjvixJmFoF66QTc5HoyDaalxI5kY9zDKx
iK7dnNsY9IGmZnuFXD4V6Hu5G35xXmjhM7PH78DiTO/UgkFtH0wZLLMAWNZ1tCaM1Ag2YPz+PBdg
3JPWEwKpllkVeMSmJxbG5KgbT0P1+cHYrzcGeVWF0U/3XZnZUPVkWt/QeJK7NgGJ6T4l4sbOgoF+
83/9KgqGIg74dEwyKkkbUZ6l4kLYdMKHvn4ym6ACK659fz92wdorv4z52Q3ShiCrAMS4OXW53SAR
Bm8rdjZEXQ1DWkLSgqzsi1RIjnntcs/i8uRLWbn9N+1soqVhUV+jbqBEavZFL15qjroCa8Q36he1
v1ZHwT81NmlJ4b9IGooyhaKSIyjvv+k5WbIQnXe5u1UCyXwiyCLeosgyagdnjxcjiKRMMmyk+J06
qDM/aXyBnyxiDWO9taO+C0t6jNcdnUyS1zwzzKaGHZ/gksZSxWW+DzyV6pUSH3Fb2sTJdmoKhgnh
TY7jaus60Od092IXNpOX8/oubOQ4KCbmlNL7rqlRdxdNKJlOv/d++w5kmV7XIOTTXb5blow4xkbP
sGoraYn2MbTIC0UtH6MVhPO3CaKJEgo4/gH/LdXqXukHApaC8Pdb5G+m6rvhUdVDDWA3M1zTXt+4
P8mQJKqfzc0d81t+4Hkzm2i/w9mNuyj9qsSy1M+/dsYi2GH+jQmGfqJN8PPe1kS0xJeaVNQ1dEUq
AukOQaNqYuyiufqQUJxzJlgkzgwzJ74APW2UQNlbrChclafjuVcfu7IEkcssn5hA20Nr0dhqUK1R
kTshtEMoFmdM77hf9y9hZ0FfXU8ZooVc2Tk3Pobw9gVihuiynCUlxJ5UAFEtIK/whPyyUJVUotHV
kfjENlDjdIB/DO2IUX/S/8ZG0MLGirtpEE3U/v3RntsTcd/bZjzxQkGGMfQX6EeWtmEA50ACnVSR
s73qido78WMZ534ZEppakfNurRYA7iawi5Vvqq2cX5heYOL8HUo8VyXGaZ1ZnS4oLA1WjVc4xI74
ZNUbN/oZL339SJCpvoANhMNEoEQwfYFUzQRJDmjMMOr9Dic1Ajp+HRHnDtNOaopKOaYqt3UZFpnd
k/s7JNaY2rhgiJTG9YaEggJvuqFV3cnrq4Q5BHMGgctqN747OeFy/AQBZwOQc5DxA1QBFZBKxDYa
c3A5lk0+agmCIId8jSb7WJOra4iXZGVAx4MUdK5ZpehuUUgS6ATtOWsBAV1H8LRARNylZVQDcGsO
2jIdWBpObW8HvTSKoWj0B+AeTa88OpznaUeR+IJVpOoxeAJLou8JZ5Q+8Jht7sa4Y6/MlEwaTT9L
quBrE0178LeS8whFA6ld9X5s61mN49q7wYO0GaOn7GVwDffRwszCjk9HohpI4IQ7XrZc83Z9C56P
ZS4RWN8hkH9wSujKKNjgREgApjJ9EL2mAOOQfk5jCze+t0zTHH4RhL/vJrQnjVnxTXdke1TErMPU
Gvw8OavnpFx8fEZ2ct4inA3lvUn7+HH1czTSTZlbvsEtIo6I9Z8k6G+mwAs0NLCo+vByPcFlifSE
bk+/j1G7W1prYvVCuktfn1xPhOVhVGBmwr5EHSf1hQNMv//m13aB2DsWPVGvhEgg8eoP9oujAj8/
G12IFg5UVJ6yrLog/pHAMFRrXeTQ7fP3XsziBEkJkjLUtvi81a6vRmNMWP2RWK8P5jkVvk5kkYGW
Z8qXqtOec43F1/ULXRgMOnu8OuX3SSRlQb7O4bUbXtczPy/DopFgyCNwo8VjMhkKfBVvLvPl3802
+Qs5OtZbGrArOrtk3vSHcKERKqnW1yCUJ5AKNW+XAmi9Wlj5qrYQvT09ECdGqIbROwzyLMZ/Yy8n
tvRHrHHHKNkMYveGtKJGcchQ5nl9zubyxZ8LaVNeE6cBmIckNdQSS8z9QWwRrUFqhwHFwbq9ycdx
Efybd8Jbsv694VOF+HpkR7OJssum9yDrApjPo5qeHpoh4Q70nxVSS73H7PeGs8chRtrk2GXCs7rH
7HPTRViX34KTVs6jGDEx3KfzPKymH+MlHErR4sr9keuNUbSHY+WC/TcgFOHM0aRmQQgRZundvaVm
m+UFGx8V4aBvJ/r+BbxCAhx8ukdUkqrWQYEpTBWmMdpJcjZBi8KZTtoSEOfI7p8cI0qhu6F+jsH6
nE3bUAc7bxRSlu003auPEnXtP09qwLhyadKXCTzW5lWS2kmds4lR+MYKu6cfxucceCNLZHnjjqS0
AsyAqDMirYrvTYYdQYqvzDetRGk0osw/9eKXkFcGfD/pZzyar1Xz7NzpyjvnNVYOxkcw2KKWOMIG
sM/7a0y7OljK8R69bQBqKv7ElDiIQtIrJFk98PpmxfAp+hzmR31Soqyx7PAjfiTMPBWsWIapIs5w
7Gke4rGujadE03VZ2h23EwZPRqZenZdjPHIU3PoJpVb9FtRuQuL5DGop7SRR66plPLQddYsnwmRk
kHfwYgz03QUtIeDzeVKY2dvc7tWjlnIrw7lYoE0uVrotulImvlMoYmxagZ23gZml4W3BZdJMov2d
wn1NYOcbRU8tni7NiL/4CAySZZwaB1mTWEnCBUTCIaWL6g63wOAOOJjYE852/H5PjH3cJkVa5l2c
TYZxYx5Bj5DR52BMkNapAO4daR7F6ojs6tT7eGxBF6WOOzMiMIHJhko/LH4B5qhehWuLIHlfbRPV
ewZhrdH3KjWGFNigfRt4xr5J+97JGsPBSuxingFWy92CJjLPomN8Bc4P+b5QynjvpXhGuPUPXC4n
jtZtue7WkAJJqea8Dw530KK9rNefPX9hPc7LRS11TO4Izfjx0kiHXFf4stDNd9/Dukt/NkIXKp66
TMWPIoS6V7EwXJv+L8URWDu0yoIouaqC07UesrZ/PMgg43ClQobcd7LZF6QaldDuKmmoFC7nloDO
68u8A5zyaDy/RxPv2x7FX4AotxjXfFVtsbEAbLPifxKqzEQp9Eyw0fw1XTZHHT8g7z+uSiuJtn/g
Ftd6qvvGPsJwRNzcf8Z49Jqa3mBz+b6Kms0y8ioqGuy2Zu5r++TzKMrcL8/mAu0YbzkSHBs9oS5i
AZQXTk5G8oBLJctEriKg+2SFsrGRonxgLRpVCwjNWHDAjBkxGTe26R1FmRzmgZ1bX6m5lFm+LGUE
yx4noaRAoJWlklidEB472X54gd/Zl8mAVruRtKxILrCkes/APFvvAyfN9uqHHO7S+TD3Fe/2qFQs
vdZfDTq1tUwIdAMR5eD8Upbi5w/+WaRqJAI8RMhSXZ6FAZlNeX06Cl+ZINoX3z/0ZVEcN35Hdn6z
G1nrt2x1XXeTmh/LraKUWfk+XqJ5N5aHUYX+bpTXBWCiG64U8fnT6kd711UIzrWkNd9QomjcC3p3
k+FqdSn2CbaMb0EUYWlc/xZBLmLI72armbyhV6bsvl7idcrQ1lIsJBfzEJgIxFvjwF2p1DaVUwgB
dHmtLeas84JdFu8to92VzQtgvOiXsK0JU237BtkIlVey7ZM9/dOxcKIntV5lrthziXIgpUDUWmSi
p5v/lulgOW2HriNLiXTb3YbIujWmfaA7+G7ij+9+HkVc8GsOVfDPcIADIqLkiprdWc2r2JwiLMk9
FB1YvQBl8KvxyU2i7v2LIOICQc303JJ4XZAERiv8IyJwNE91q2Pl2kTXu+PBhQ+dez9UOXFbWieY
W9sqk8IFum1ZD1PWgWIUUbO5qXWeT6ru/FwHZZ6m4RZPwta9arswf8C5MrD64e4rlkE+QwL/SFLX
ewKJUYCOlOQuJAw+u7hwwf3VruTZxaBxEcpZ2lFIYvuWas5OcvAjJlmf3EWoWtVYS10o23KWWxDo
HBgXI0Ptg6WwLjxotqIPuwf3zjzvOOnctZhQtHpbPLC10vMMvEhaNNqsEuuuDZrx9GGrRU2Xxdh8
IGgrTWulU8zanVWrEfWApGLOyEy/Ijob3244tt+Gk09JK7Ag9nVZBJkPE5yt5XdHRrRKaD36iY4Y
lphXZrvOLy833OKPnUayDXQvRWOR0SMzbHwonRp1lLbVadrazaesel45XPGQOkwLArW/QiIRPxaP
/ddHFQC+qexObM1JFqmVKBUYhLY9EMmMhq0OUgoverWitW+JZQeBSD4vpW0r9B07LQtZRSqu/y/W
3JQuyXQDJPlh1YEB1rK4IAc2KUTxbLIoAQYLtS3Ekro/QspV744a9Hz7g3xuM7r/RIN5waa8HAjt
tZPd90QsgY8+nGza4RuKBlegt/fJfsNKCdkPcVjXG/fvbdR+XTV9wRkUG8Az0vgi4qDn68LclVKJ
9aUHtW/X6UIio1lZ25NDRgcuF8gUTeX8GOaMXitP3M7Q9/ZUh3ZsdqQJMPHT1b9wvhuXbeywuvSu
wFBbYEIc7C2vcubbDYYQ6V+qwdf+e2+ppJysnML3FEsSqQAmDAFBDHFfWMUID9tV2zLwZlxi0qvd
/+KsMJwZx7SK/I8n1G4n9Xd6SYtU9REdfGBBJhR2cFKRLL4EbhLLd9dDh6TWOf69ZyHgEg3od7DT
U8lVJfQI7/iO7e3o8+xKFARQr8T6QKWN0uXIQFvn9x7xzz8krfZxIRVvNfOMxbWk3n82saiQZIIy
cNWymyYaajNdyC2WN0UstEzyQ1klR8htJ+gSiilm1fJgCC0qEsHdo02wKd54MxeCbE0vJ8UO3sbb
DV0v/t+gWHB5FsS1vjNbn+h820aqzFqc9bhhP8AgJBMaBIt0HcnrU6eq2lt5J4KBh/ox70FC7Vdm
YK2DC4vcMX3iyHF7NegjX33W4psYLJFFEXdDLYqSnukEEEqv55xyugeBjIfbKUk32xnOLbV9Ox7D
tCkNzUYUFLPDrxG4l/yYZzQILWByNdMlYXdP5w3wBzVPcKIwE7Z+h3Aj199ZC8N5rJtyuJJcV1xP
cq9WEQWwX1oUOTayClso2GDwdlBifWA2w96DO209tgzL2j7gVR1cB93MrIjI7tP4ebL/wnVaYQPt
wEieSrQQ/Bzynt3ivXdh8HAI2ZXdZsInkdF1GOjFjDDz9Jb2oylQYU2RdzVrhE6gCIGSOzSMyVHP
T8Q9avY/fatBQP+FoGH8NzYoJFbeCrP++6prSYkik1AU2CfwUA/Gd2v33VfkIJOqA8UmjhJDyL7U
WfNIW3Ls2j1kAiliQDcI9BCtdvnWlnY//dKfJ7OxrZlPFLR1kLz+j4tGYqZJ8o2ZaRIA0eLyHz2M
BhC/fGlyu9wMkdYrn8CGlk4/t0+Gc0tNQrwJBi3GQhP9WdXQKJdiaMQKIaYqkcSmWdE8fEECL5rg
ig0FQKHdqWvLn6JdAZuIORSwDGKKaYrxId7ZUnY6lFQDAM8QZR/FcUJ0fGRltNr19xmRZBrgdIuJ
MJ771hhcNnPtzQdARny6zPd+S4Rf5KQ06hNeAMIY59fiVhOOzkYNwfy0cqIE/ShnwtaGBMxzIvur
UYpFG6zFsLpTfPt2DqA9AJRX7OV0fyOQkVtRmy01q8fYCUae0mHjy2U7dpprRcIt0P1vVRAzZ2sp
lKrT+CBOMPwVrFJ2I0J6SDSBjxRMbZ5tplHUiQXOwsVNzS88Bcg2BWRnHQwxxptLm+X+yoCQN3St
ywrcF5TmoHMHlS6+09hSVLQmBxksR9IZBoTQccCfOnG3vXUS1liAnXQghjaL5iUN5lyqifDTozCv
EiKoW4ERNeRnV0kawfrjV4S1oVGibYh0assnBLXCbYPNnamDxHZAfNcUb5/9PvvZyNH5+i1E6v+s
nA5FR0J2Fg+mvUwe2Zbd8311geWmkBHfwkRqiD2HAWdKuIHV4Z/vtTEK1qlZUY1waUjhye4fvLrK
DueqHUr0YBB8pzy1izjvMu82/NJjDdsuT1t4XoPg6wVdUI99CL+oW7DEVSlWgdv6AFlfm6kkVBXV
kGJM1YNZObcqal6j/oTDX+AlZdzfgB5vs/oG0Qr5jH+MBJEn0Plenk1KjtO5NqBCCT0P8FSVmcEU
wgy5ndVR3K2bj8EdEugpxzNcQtyhu0kM2CZGHGki5tTSR5S1kM3eReKQHD2e7sbmI+44odQHkQaC
UQvafdNYDL8+pmLihY3YMe921pnnPc3RM1GS3eQTfoCcKnKBZxOBASdzTzujqFjmO174PVC70lK1
QWIx5vkA5wgnW2RwvaqgcUk3afmgJNZhOPlLynDqVKLVHRFJB7a3byWmTKXzbkw+BL6YMLHVKG/E
9uEyyghF7VTPYbah81xRBgQ/vCuqQaf5HB3ZEs+HRC4hmzMnHr5zaA4NEOyi5xwhdxoRJMCmIM7E
uJxLeFfpJKV4XGYsdVZ0KTXCeWJPTezJR6DK1wV+rx1QxuwgUMx8Y941sfATr+cE7h32faO95bV2
fiU2e6LB4xc5BBOliMI1ijSz3ctEaOrsVb9VXHtWwHa9/7GtsKy4z18TJWPsDqtNhBsZwm8CdUXV
f3eSGU9nAX2nS4QYwlKIaurOm1GJbSXqVa06hBLooBHeRAb15SkCclTDofu5X+xb/rHEN7ROM5BK
dIYDo+W9+sOz+Pox+ih12da90yfAyvDyo2bKXmkuMf6VRjl8pVp93gs561syp+JCMC8KkuvpUb6z
3V1XBtIl3RzBgSbxar6SHUZ1JolhzFWeDODT+lKS/j1s81Gn7SWyVwpwTFSN+0BDoLw/cdHgrrjF
1ih/gDgj1luvrwFV5agFbzigvYCg/rtYt8A02WHj4wzHR/u5RAck/jXCJWI/aoNKdOwsBpUjnSl4
2i9J3GVzc8sKyVJxW6F/okMZiRUDK/mtJLJwzGUk3Oj9eKf0ZSoyjLb8jtAwvdXb0+wuGYPokTr1
yotU8T96je6vhZcwJCrlCuy8LcXODa6EPR9dtpMa215DW8TrEmIierMkR1JVQqZhT9j7xCGeMPEg
myvG7IojKtqfWHkdGg9cLKX/aec7pwDtKI18tnyY10ACXPIds92s3BLP/3G1szHISUgyBBJtwuVa
NNAqhVvJig/R8uwoWTJUJpQRFZ+hZToIvcNg5UqvUdiySU34DtkeSHfzpzBzBiifJ7b+K3pn+nUw
f8HmGV7PlsaXxcq8i8L5OtnamcE0ScbKMJkO/H5J/XTnuM5dkF2W5gXpkks57ese6/JQBE73wRlv
pk3Hs1mg5a6neXvMLupVYS7koiTcvQFKC94WHUivFhJ8v9lhyvMGQ/VMg9dFoeuNAaue79QxFYD6
vXn6sHT5Lhe8xUvAZPG/2ziI0apn+3BQ4ufV0oKUmNDVx0E7w7qiD4SQLBswsTymlbgqmuL751Fc
3pMBk1Y2IuL09DsxGKg3EJD9hdUH9vdFy73nuuZcV38/Ae2XqPeF0zBluUSGriRgQQPOppuF6mkq
FsEenvZpoiEY8OKbO6EL/saDt/puPQR1rFH6oaPvMVKhtytWK2NRYT5CqP0SozotMewlW9UOd3Nv
Lfh/l3gz32BGm2cwbejQ2zTrJNbLbAbSOfhfNQXf8VEyWhUjLezm7s2RNn+glmnNr+o4wO4Nt2uQ
LcjTBeYEv/L1auCM8bHI85o6U53othFYw3kSn2kt8aUfksGJG4Pv2292RwuncqYQyRVwcUaX3Ko3
NOnafbnYWS4c/IZoLufIjwRcNxih3eyCR2rqpKO900J6wdPBJnlLLsWK+Dny5EyTBmQHsDDXdXYA
nVpSGiCi26kUUAJ2rHTWxPrvaSRyLll443WV+kw6k5TcDylQ8o5SxjyE84IzJlFnSQ4mGS764qUX
TmSo45AMgPFxJr15YlNpYs3XtW/YQUyi/N6V2jAGNf9th6hy9XRjRwH6M4Zp2IaTGMrDYw8Y08Pz
V5zDDIh1q6Q1iutEK6BUaFWVGTYVtF1ueRJKHvLBUag+zeOqNUIWshmeGSo/TGcHxXNP9GeR5vmB
tZ7PusU7fvgtYqgc87f6rH77FJGC8Usv3+OodsS8BfO5/H9woQjERJXbv+J1WPWhbKha6cGtAd0q
x/xxrm0tN/UmQ9xh3pKZkaHG+1PHl9mav8H6GlcsZ8RPVTzekww76DfluzE5A2WDXtNHwlLDV09d
98y3czR9y4++rvv5bq4N1Bf/D3r35Ym+RzgUd8u9qIK+/9Kj0XmkNxfqF7jAL8XnvneZxdQTq+QR
28NOoAed2WXhvxd0zpDcgGqzPmjRuZRlR1ug5pZV43cWTDKLBn0/2lYIOSjF4aZsgKRrLHm9VwJ3
0WJJTX2lIq9mduipl2UEvii5Mx5tEpqMISYiwAVSghmKlaNccsEFKH/UDxz/cKgQMSdxXOfuwHr3
jcsJbfK3gbEwDKrr+mWtbgBGFUtpNYCKi3ndV+ISk076eVt5Uofz6LuMcVrHr4awq+GEjJ67B++a
DsM4RHGe0cKbP54uU1A4XGQTXJMk2Btgp8HYDx0MfQgV7p42Avne8TjiDBFi127ea0Na1/JngTS0
Vf+En721QKBLng+XMy+iQamFl69EmQvNRIAnt+rTzAgUWOpd1u+wbJboJdgzm/r3MXalbrlOMybl
O6NXmqrKZNNhC6lbcUrUvMWYjl7L7j+EQ4YtKfTAkxrakxIvaLAtohZvc2yxwA0B1LwFNP35Y1hh
ywG56Kk9HnK1POAkyipUsFgKpmEF296L3CVGfmSl/A4csTb9I9PHw51JZ/IpA8xAMLHQwrhqppaw
G4CAMypdqu1KXTGvbVx5oNgLiJ+Qw5W/+mlgYxMt7aRyTf+aWdvPtbtw9MfLWQPvqe5JaXrpNA5g
XXvuAov4sC3aedRzWSzhNvFiF01emVZfTlxc6x8TTEsxP2NcScvSXO7spwap9xH3/LdEe/8Efaoy
7gdECzi+d5UWoDqtSRvhMwn0Ig9kiJOk3C+wW74FwYmsdmAyipBpqmXhQz6GCGoLAILkIN4KpLbu
O8AXO7mJd+sXnIkWQVBDfNclX2bGLXD2lX58ketu5w7agKGczGOFyo8c16S2q2RIVMjyZIXLTJeP
Xz+VGzyn1CmRt88veysHeKKlsCLC5ciW+JEztOGXtBS4EbUBlXqi5uJlkw8WsdDveeD3Aid/YXnd
d6jMfFxhpYhTX2F5g6XICJ1TPIE0OvBedwk5wvfQiYcgHpVpAUpIfX0wtos1IJL9bPVRDmnZyPpt
VsfSutTMEf1mNicM3wv8jzs8row8j78FRIOKjJOwIU5P7Tevml4qHBK+U9a5chKL8a0IYDm8hD1T
WE5/wMC4Cyrfm1jIIuinjM3Bjpe4eUSLgxXCCL3GUEnVdyxWaUjXoVUDb22pLHRDcZNXjCp5mIET
HHKdtvSW84LAnaGBLZG0SRhz1Zopc+Wyq+YRSCzXD2MOXH+gLEelsYi3Moc2p+wwTmWrEWzaiJ+2
h5zBfT8w1mEEE2CtLdg/+TOYwK0jOrZ+uY008f451HG9zsy7t5PJJI6EZU7f+prDcLTxoEn6hZW1
UdhYKetlweFR53TlwtZxRq/6dTTT6TKcaRcw3W84NtRwQG/z+WA3fa4hebdcU1Hr3zOvdrFb3wCp
iPRCwIKezqVp8hspb8Ugfo4bo4R+EXzHZOp8WYsIH0G5ZQj01I0eGO66UMzMpm4G4qgsf6XH2GPP
xaYIMjZJWmZmzlLA4XVTFQTBjeYjnwWMG5ptroJwQt5klC0gosW6OnJO8r8o+K29kEUXHLXn4yAm
qbHIwulgntUphuSYQ3sez7SEbG3DUFpXKlhbeVdMxM2C+UaUTDU6arXCywFRlSWZaYH1rWvHr+hF
B1ysOn3JRxtoB9ZkQY2/4xL+FtaETkPUc+yQSVrlF2p9RNFolb2ijHsJDBJLJSUbJ+NDm+UcRw+F
SUUKAKx+CGdQU5F4T9ErvmuedG23sffvyEEj7IglldjECZ2DdmFDVX0kwS9fLQiWkgqUE2OgEbyV
aL7iMW9mz1+KzXdRnc7nkqKrzoPeY5yiQ0IJz5vppHTKZJzdn4KeoHPH28g/NNC6m+xJNPku2Wnn
Eoek51UyXELtGgxP2Nj1VRJAfQHVAaxXaW38XWqM2eZqThj2Q+1YFEKnqoM5iGWLU3KVBvie42DT
3WMgxwW1J7BicsoNe8dKtlAoO1HRZSZdHX4q0mftdjmZgBrUWhG0Taudlt7qg2LHX6HeDIu/ETwA
ETNMmn2F3AJTUklz2gVaM9aaJYIQTl5avQ5oNMa0oifAxVczAGHZyHYaVCaWtHLFlxcQqKgpDo4V
eNN1WnFHA3x5sIzFxuFj3McJCH7jjAm7c6vqeUt9J0+0rBwTqCy6J6GuZKDCcU6qNnkeUSaE2G58
9+wnOo8iXiMpPxZQBQu6ReVLhb7hXw/qwHsXAu68+BytjbB7Q9TsIgWg4w3a6SmnCG8fXFAznGCn
IyHQVXwUlRQhke4qlDry+YEFCvOiS1eVtOSaVTQHLZ+iLDpCDRgBSUpOJN2ClfwEUrclIzMcYKjU
0QX3HUm3EYJjCM9rSR8MitDJNWcMpeo4RlFAjDwLMXHsBcrO/ERxl6sY0lPdrW4CL45muSmSXppH
d5bQvYw76mx7fnkKBHYE9sgVvhmb5YGiTf/LgHY4VvBdlLf0JmqxDRy7HPLaKTAs8oVDZO/3dglT
u3rkFfVcivETaNa7hBGYBEibkDFkgZhf5DqiLzn358tYxjgwk5Ck7AxvfIM/JN7mEezuqeR/n2ix
jJkd+z0cUdnu7YjG803/4Goh1OI8BDkiCCIrC1K58x5PuXhh76rKh6BwZO7PNQ+j48G9dfyKYyqp
HyX9d1VTjl6nNdtC/nvOt8XqiQ+AtcmuJ241BgwpvryZHQm6EIiOZ9cF+VGZ6DFQhnPDDrG0V7vm
RER2BgOPfxX25ZobqXyUsVnfH7HuplTl1bSGNA7lZJ35ZLkgMOynzazlWC2rYv4rOTo6raitEkXj
ANy3EbtzEwMPeoojmBQfpvX4DRqbnHzgkLNytyPr1c2oc5tSZXOAV2E7spd5fOeji6SXeOqYj4vK
HinTtOHH3dCT3xoeSdeCTp3BdSk/sPDj3+6Pt41XmCfufS6C5mE4fLFHDwQMbHY3sJVj0LZ3Kn19
OBzDrT77FxZusTYs4dfXX30882WLRfzF6ngFk+7jCtpbLJTOfqIdtNM1o0yV3x/0HKAPDR9dLw4i
OAGgmgC9haOYGrthlZQogUUpQZjr8ggx+mRCMda+6lN1QqEH7cpmy1bafBPysmR/zk4yCjkGrcqI
1z+dd9AdlxhYgbUED6z9tpoHDdFhJyxLL4iTdw92U5hv5dzNsL4VKP1nxPhYyqY25aeyNxc81e0E
a5kANWwA4/f1LePiivdcWAY2skNpdQwdXqtfr7SSGaVe8Vho3n3E7umFuGfZTdzWiW3ywJFdGAP7
n0PZekef9jLsOnkT+3oGrfS7z8oCKW/IPNCFPhfYYNW2vWyIjntKsSKX5YvOumuGBYI+o6c6JW4+
mnptKVIxCjcF+qpsd2Ds7Nq8pxhKbeM7gzhNJQZ9+rTVUF6x2PnykLI+VJx46P7C60Oxf46Ol9D3
1qLkfvDOLjjpsT8I1KgAfd38Gg66OBCqikV9g2xF1ihpIdvYzpiLy0ZrxAX3eQ53vxVop8SWAuLG
I4h4Jy++7yv/yxllCVzzpRQR+Aso+3bpr+aPUWQVFqVdlUb1XGFTP7uZluypXx7p9ABj/4ZdSQsJ
OSrAMgQn1aMnorbzmnSks1YfxW9jXxKNAPm5yxSG7v39DaLW6kkKB1XrdFEuKIgbJaL0L//NY/O4
51yFbVR9AShni4GMGzt0z2UcyPKcgDFhA87x/bb/YOxAP/xfb3m0Or7Nzbwlg09x/4PyBsXSG3Lh
6zlkPdxfSIvk1Gf4zb8ReElyeqWWIV7/K33z0kUPtN04xcu+v7f4oCPzAMsMiwbzjcS9y+WrIGcK
bwDYwkoZggdfKLLoaSdNkiSrTN7cWOkE/j4U20RBHYEU2XLnE2S12xbJDxv85WOBfdLxg7c7SPKr
mT4VM3WgSy+GUnBIFUYKNH7sW3EhljLKH4OjaqPsguklMuCaQth6P6pO6L72pPQMm6LiMu0zYTYZ
+orNJ+7T0Ka6eh3Hos08nFwoUNL2VB8/X6mxjfAHZTsFLwqpFbQ9Q20BiXk3hvXPtntai8YslUyG
de/nASb6fkjpFCr9lpqOwtqmbBNquASRwS+0pY04v+sshEqO69jZxyDBRUT3PRUab0hJCIMDdFmL
aFNJxRyLZeAAKrTsR16MCMw7PH3ZEZLhrQfVFWtvJ2Idb/p+y0fdZeTz594EHqoI+DIt1j6zBSbx
WTA6JxAmbn4wTzvii1AUKcW9j4iqdnviegQAjuEuVpd9cQyNZaSCUZ8KrgdwwxduuKI6hfnhfXOQ
Q3rKACWqqO5pjIQGUv0ujvG2vt+vOl4hzPmUC2bXTer7W5GDH3ywt1FC3i05KiMhuOn6NAFdwftL
M0OmGsZaHgyKBDg5LkQzBG7q93ziRPQYZ+ivFgL/t+IxdeILWYRRdi/0Y7Gz4k4CDYFYuhTv8pCz
wWOzoCvIpMFfs8mwbXaH9jC32qZ9a9nPzBc/Oe5/JDWlYQ8fDezo6phALzpMGaz60CcCIkA4/UCX
oKSmbyWHUJM8uECKA4ZfH6edWaAaZxAgJSRJ3mCUQEDg+jfyZC5lNaiFtdUQzf5sRoSugCn37S2j
BaspfVelUTPeMZcU0iSYZG/iWtLGBSQmfTSmk6OZHU9M/6HGCKkFGUH+cL86azi4IoE90F8DQ0G4
n/A3dIDDbvuE2TfklsEONDP6vmKrCs0SX0uaonptkMsThPhwoODMnaEJrM9hRLTarSwLjuOLi35a
mj/4a/H27FDF0CWsCgAGCVUhwV+4KbSASLup91B6qzesgy8ehbUguDzwrFt86o+YKTf0uN4WcngB
lCgrEmEHgOlXYeVhylUAJEvvzPRraSfLcNcJd75vcavpol2tCZmRQGdioVDCyJIgVgYb41FElx+g
PjKkZp6MZCIU2TF8NVrOPeUNMMuca0ZM5NxRatrzG3gq2Z4ijsbGDEk+gjM5Me+tom3//WlG3lhe
kvjiPUnoMHSONmp8mOenpS0jS+FstQOl3kWmHx04nDcwhSLr6Umw678uPEHVFk8YEYUVQwH6DUvL
QF2U+ShKpNf6rWrl5/pyKWhsTMZPuFHl9s3h47dwuyT6Y1anmaE5icF/UAW1yjEmv8l1gAWgAl+6
cxUuR7ZhG8OqsJcZn8Qv5/sv7nF3pDAUpD3t+jreG0tBbVx/YxVePA3C3IADGE9YeqQftXkepKDX
3fOifw6cvgnNywULb3EiKHZdveW9gKTL97EWocPuvUQmyTVyqhO+dJwGpfIx24Vn/+0bUU/6cPWx
QTDWADDO4VxwlRZFz2ZJtrJGg3whcV73vJQnohAuQdUxDptEjB0JyJHwNpDHlNlXDgMcJ9xNMeuj
APf2o5HY+o/L2IwBnzroDy9KUk/vZNeEoI0JXwWnJsaeJSAMguKjuq8T73QdGQucpEkbXaFNRI3l
4CVyPa/y6kYeWY66FwligEf0LxoJaiae+yVDuhI4wpnnW3yWGoF4bIj6hOPD7Z3CFBfjXYpnHGYT
pNb+rE5+7tJzcHqTKhLtU9LZ4UFeqhWAe7fNZP9U8MHd0P/6lfcZmKJPQ1IlR++nBP/FMt2FHK22
vZmFNjV1UKWZhOzqA6WX8oDz2OUiA0OgZf3l/KcHEdd35pt+by8+e0VwvjD5JstVmcVhQ2FHvgfD
bizrePqf2ksul/e88/9OIhRygGWqiub/GK7s6uWuRrcZ3fClPZH0yB6OEhMF2ivGYo8W84crLMNR
mn7BE4Jtg1b06b0yrx0EBnPM8aGUE+2AvknsglZPazu0lk94OITlBc4qaCJaMVrs4WhV2FPxSyJf
Sp+MNk/4N2TddoCIV7wUS04cR4ytOw87vm7QGGI+0heWmfAQqj+yA7S4DncKAtHBqrWD/DtSKi8b
8UDtdsdUO41VrhjA6PDUNRRJwIgqddBsQT47qU0vFGSvuop0fMRLj/rdBFxQai8wb8RXgavuA0iS
waZNM/j65LSIe9GUdVNrGdU4BNwKKhJJYfpdgXmBNa3JfBiCcijtcnkMMyJOdqNWji2rnuBb2TtJ
YSDD3M3aGaOhEGI96HG1V/MT/nZPzd2SaBLuAz9E1Xl11PLWMbBGCNLx6I9LBS6dHnSA95YvKA1e
H7522PaiA6gOc13BcrnUdzkH2LikTb7J6uJ78mZOIe7Yfh3mnB2XIZJv57FVJxkOhN9t7BNCdqdr
lEJzCTKWuvOQEdFs2kuks+JVfc8SIkDE+CVvHxA/xbUY0ff8viR17339lxAazcaprga0D4l14tei
/7gQUk040Of/LY8LuPk+ZBDyL63HTAiRI27QCTOVF59I4UFBeSLm2gC5bcCRnaLeiy0LNuFV/CTW
OsabJLSWijww0Cdn0TRussPqXFRWEIWJb2qgo9zVZdMy+JlLS9spKfFSVxJobGkVxJAQmt9ih1pF
V/5knZNi3hK7Gv+wCq/cl+ZP8b3IqA89ZCc7gW7aLWlm/rLUe9m+pGF6zbDpEBf11huDygcdjdht
4GriyIL7Y5B96yyDdGV71g18AHmTE9TInFIi6w1alZV6Ntj6O2kwrUeZxPC/39NruSi5KS8tWXcr
b1aGt+yVU+mX7NXsJP/EUKFRJzD1F5/fih9o2pprAAcXpVR1b9hUTIC3cxlYbJAybwvGqGOLoA02
sBGL0HaaP3UzaK3i4uwgYy77P1c+UtYAYus4znYYCLbqXHJDUH7v8crK+IP3jw7S7yNdDcwwNGce
kdrCMD4WNxiHPBGOVJVkMB75n5SH/CA+M963qK6FHuaKL7WvNf5u7SKVBZXyESEh+aLR/QDjoaK7
OcBeI1A2jQt8tPN5g2VDubRHmH1Ip3OexANYhjZwzaX+OwRjw3rLbVfNs0r6+3ByUgbdO50lBcfU
+SI/5Hs1PJwURIjeBQLdjDN+IMYcIiUyGVKOJ1f49KCgR7WmepGtMIqFGMsVC88fA6aXhqR4JUs/
OaroFtlkDXdERQsEnPpE1X6X05zYXxLlFaftwT4sF6eS5s8uLh/B2e4PAB1TnYWRl9j6O03ngHZn
SpUTQvtD7AurLWq0tj2JmaNzMp5ZPD7oyTVG6j9MM9nU6QckLrybfs5JTjdN41J8VQqIc83pbQzY
TGagV1xlhewjatCWyhCq11/BScrT04Hs6+CgMliuQJu4UBs57RPX20dzNUAEyYZnlWHo4JqfMD+q
ADuKAouFri3IjfHbc/eCL4oRfq8x6Pk9ze4ypPeCc8Yz+nKjvbLGhStFZurmp2Db/pHgQHg715we
NfmSkYBQawJ4RGAheVhTnz9lI6P2Up5rnivo8vthDsWmGH/FEBUW5TiYY12kWAJVerYZFKqzA43Q
tJjKyEMrgVnJCw1u+pGCdV2sUZtr0KLJ4CalptASbGwDzvbM9eAbAD4Ti3ZD4FWA5I8K4CB3rR2C
6GbzSXH5ZgtLggiixqCbXKv5U5ATCNUSer6akhKZwfz5C3kkqy8RXZ8O4C7Ae53bNKEDbVc79saU
iuZu5YdszduPlRRcMigWJ66jyZZf23OwgQjAi+ac+MZ3yQv/8uuweQMlvXpA8F1W2kc9ohEXFWt7
UwuStaHTGwfNQ//GsvZBvMa8KAJXX+k2WXaqXDD4HlCfkRoIY/tlO2TBEJfpI1NAhVp/5pzeYscH
/Yxt+9uY/XLGQLp7ag5tX+K0MnotxRokpmTtMW+v4cVFhhF/JgLTi1+T/zSZMLuZ4nmTDyvZTF9C
JxmrzUs47bHTnpqjevuIOXVwTe9APaZxYXsCjhYgEWImqjZIQsGcjHGu3avaHzNjvO0Odb62kEN1
YrBLdERNh2KRdEtJ3cXDmx6YrXuza2hDzJS2SRync2HtGzKLcrWVePJxftvs2TGK0DMUcafDfGNR
eLqqIkF+D8bE+baGsCCkvDaRiCbVK7+eyjT98Kx6kzOs9QDb8/uqEjKL0j9RvmahuDh9197Oj/0Y
laEdmt50kZ8VWVD/ixh+m5O2RCLyDFceyqFox2tMJJi2a1XwVLzpBJLM93plOyyNU6tS+lSzXvQR
dS5cNZouFLw0W6n7Trk6MvfRPWZ+3uviODhs6EUbxlH8EBRmT7Mfy6v7CFi05scw1qSyZKczqYqh
qDSIEcKVx0unvqHtO+T0DkgucCvW5b9jqOmeno/m1vEDxlgLMSfREZmLLh0eJMm48urkE6nwuaII
Xd4mgXSuGLKfGePESo90Cax7ShCXHlbbFZtJfMvUPvQCQpB0xCo6uPEzWGimuW1FzQ5PnlPusOOM
6A8aR+koFVvv1WMCKpn5C3ce1CBO4ALvYn2J6/eUG+AAEv682L/9d+XrARK9KbRvx1eupUh8pu/r
Z8gALnbw9bZZoXEbKgjEQAENCXj3c+2CV8fpawhtEcoXgIriQX36KNRkMjZ8UA/ZVCk0froxrjPQ
b4+fVYbdRdIGWsPK/lksArIqOXd5rjYrarus66IfyPn6L8HzY3NJPGIVU+hhBAjVqNLVNcj787wY
WosQIVopeIiejFiuJZT3/GO7y1tiY2Z4bji5oKvbx+IqjTwg2Y/zemK1jbyGJQ8GeLG2hkD4JMx6
W6+yAsmxJcJ4W+Im4BuA3RSzg+IEK3U7w2daO6gKj+m5wucavB69FfR4OcxpETltc8RPw7w1BCMP
115Rc5GTiJgfJ+mv7HYbYqe9iKZODL4x8AvcaMV8YSU4Cm/HuudyWuuyWq4K2CpA8dRiA+2W65nY
ieIFzL+GU4Ucyj4bf7V+0QfK2iJx+KFEPm2+31natHnSc+XxsgtHnCyHItYlAW0rZlx1aitVUXmf
8gWSECrMo65q8qPYnJk2C/j6qzQ1bwsBSBOuSOA/5aLGAlCLo4dP3puEhRe7QiAcmOSD2NK/ybtn
k1bgXAzG7o+hTR5Y4lHKUi68DKTMmV4SDdVIjOdaWCe4IA0Fe6vThZEZ9yNjzNXb6/vlWI7fRYGq
yBa/IHQFCY5LfNJfN/CwVSEGQdV2VZfqRCfqHaqYCJWL+46PX4VhxLajRNEunvPbedZzqx4k8NTt
9GVABrkCCy7fvnVuijgVcr4w5EOg/Z22oe4y0ypFzqCYfaCKdsKx0746PmPLOm/sjm7t8CGVuCzA
vgcWsJVhj8l3CUXYQXFSH5PxFxqWRn7PMnjkvj0a1E3SI/3/QHz1mX3lhuwq3BKVTJkXPG9A/0/x
P3E3d7+eVoHzumZeL4cW35XslgRCT53xCIsdCwytCuZrQCoCwxCV8v4w6rg1grjnHY/zn+yrUWkO
TMOQEP3zCE/aXq8HSvrw4ZNfsWX/lHNbS6Ej27/JFXYWHA52n1e8JxkUn31ORwmJ0TfmtkN4KVId
Pv7sFsGYwaBqj7lxT0zb19fHUmGMu4VHTXZgn5qv1cWiLkXQY9uwekqxeWA0KIGloJZLKTMp6k0z
yxZEBktdr67GwKqmQfepuuU1pDIAkHDPI6rBsTOVFJwjKlc6VKmRo57b/ZKOJY6sWwQY3w1PEQBv
27K7e2hIhSjaC3oXunT+3m6VWasoAopOSsTKVhDvjYhBnDOkoU8xHKd44VgdXk5ejO2ek/mpnQ68
C3TGOIB8TVmsuNoBvCZhM8M6XsMjYXZmiJVvrTZgcBpWhI10uMcVgRTfwap3rzgaXLIKoqy75+s3
zn1r3fF6G8ED/t0EGTcvCj3ZFCEi3lVCioZ3DFicMJOapWhGzm2i6zxBOMPJiHgZ6ahgsLokq8R1
C2Vu5Qj0Ex/iyjoD8+msmQK/TRWhr6XCc/yfoh7976hRwvnFNrBzp/acuvabdK5RlR1UcV8BsYZb
9/MRO37Owxry0sh9DM/bmZU2avuRH2TliGTM9j3WDbhoJOM4TH0Zs8605bKTnFm6/AZjtjCnwPWe
HTT+WxdCPTIpCHwnmTQxpii9Qz/Q3Ga/dVuvYyewDoRKmjV63zYLYys2ZwFJPNPsHBEjP8uohEc7
/vAc8ypMq6zVH7SkgMYKkBE5dauICHGmPJUJWDjD9kzLuZpQCITywR2/1dvmhN+nnycYsjRYA3qK
ThlAYPoado7qjgtSsEY241DS2phoH3Do8cAyQRXSn/HytLxES2waBMeuHjrptkWs7Ib2PNnYe6XI
YtOFKCRJ9Fx4j/Xlr2NqtxSr6fSPP7uPJEulmWoHRath8VesxDVEPRn5WSA3w0/zVLycmpNn6h7A
zWH+7+1jBTKcJQNIpN9ZfdM/V7NDt25sMq9p06JhuQqDXOvHWiyFvYhxT6Gb1o0Csqe+DUrR6NIi
Ilqqu0Hbill5aqARQcC9icA6fMFwuOJjZfJuBIKzczRzfcTlCk29SPWLC//Mni+6sou9nFSFRyBz
YeXube8+7Q90X/LFb7zNIfHP54F6bBxjBsgPCt/EjKuHYmcsGi1sR3soaw50yQ8NtuIs0VD2niLI
I6aEhwnERVAlBesuP9z9eeGqqykRpUiEUAXS2Eu9xGGaw22NALFzYCZOBVDTJ65aEVdQ1xyVCnGO
jMuzZZ1/ywRVuFHkKdrME7W+OJAcsFQjVyYt2Ta/8zTQmxhz8+955LjMeud5fw0ibOxRKQZ5f8KZ
HQW00G9vExKohBVuxRAeh4HDF5Ena2ZIVQKgDWbY3luRF/WWCBK5Wr7lbb1pxFNYVAT0O//UqgEl
3/WohpQp/PfrJlYZ/IzK0OoJryhD++9IiNmaa68/6lXt6v/zAVoytjGRCKp34izxh1WxxxX4yFQ2
Bzwm2Kq6mzLsY8nj3HsJTM0welb+j5/hpiZy4BOS6TqAbkfCw8KWH3MYDh6OiegDaYeQLK31XPTM
SvOYVbFCR5/FrS86dZk1K0UbRovzw06c94rRAJOEpAgqIxSB0XECjDDMwpZuDhnL5Bar/wySwtKC
1YY5oD713oM1+32aIs7cqKuvTQx2BCnyh587drgJkRCvve6vayK7u+dfO7JUePXbdAymLTz8SXGj
RjRnA6f7eHWLBiQKtQGhjF1AGMLLnWjCtcjaDZIIm7b3U1B54zTYYwSxEswdZTncuAvzppmRFbJQ
FesWp5Q6sMSDJvUSYhOSnAMoGwxcQCbdJ2/FWBsoGlNhQ2zSmYjzU2M7KMa73qd0rxrCj4TcflOz
77R7Vs8LKh5ng4n49rIgxCypp+rBhmk+vxwi5sqA4JD5it8oFgzNhh5cUgpJ7TBpXY+LGHg05cS9
5/m9vJuCwhHEjxFKBCqMWINZacoiRDzWJOOmFa89PtNZSK7Yi4uj5oNFTXRyl2pfZhXhwzzr7wAm
mqlgH7gYBquu4yrJLq8tqp5rqxRb4LUGyw2LYJQgF0BlaE+SosebxOIr8CbheCteKETEtUv1FWek
/iggTnFmmL0jvsuAa8aj3CcsAEdOK0vduy8VfoTlXsSy0E+vcljkhJr+QlJzm8eZeRZUjzL/tkpF
RIaeuwAQh+lXoPY5lJ8iTthTOpBjtKdW8mEi4laePhS0sDaNlKjd20+YUEoWn6Lcq5bcqYh/Wbzf
YoJc3VbCSlbCKMU7egS1L1v1t0zoQd1SCfoANPO1CbNl+jz4rpaoRP8ecaMpZD0ZJNar9nmfDopM
R1Uv5in/xHHBC8guxeosoSIkP7/yBYAdWR1ix0WXeFhsiAd4qnPQAMtGr06M1X6XCSyY6NMJJNMp
YwbOhPHt8NV8Oe2oT9LUATNf10ZBs4HJzogli5KWnpTxeYzzS2JltKxBKqBFS5HzRJ2yeUz1GjDm
epuRhlc4bEqQhOfAosLgPhO7u5Q2ngFa8z4OmHyEFQgWszgh6QHrF4JDV7UZ3MBpJRcM03twvZ52
QX9Z/+9jEZsShUI6elRR0Rg3lNPSRn0AuvSFRUW+W93heSoiib/MVHhTwhQYBp3LSBT0scotGelO
IXMcZc7qlCdV18TyOywAbN1yUMxSRIfqKpWOeS7UMoEBbZFybTJotOzRqeL+iHweR8UijUldlc+V
4Mnm/8U2eAItQaCmeAes1+cUlX6VhRryfc0XOKBBpg6X8GSyo3eWN8WlIbcGXCRylGb7GUywH5eg
nzKZUrI2c+QWRIQ+3p35IgnVXJW8qTr9OK6wW7MLmCqVGHZwF8/hFlqoctD5yMr26JNFpDTkDiRb
2aZ+/Dc2JklLj2b7gr5takXiH4kM+/9BtzK4ioVm/ac13NpTD4gzWU+Hpfh+MQGLWzh160JuMsRq
jUzaxP4nKqyODVCSC512Enq2JMDTBaZUA+4pQafXbSnTa70v/OBNM9IHlsWBMAYE7nGouK3R8u+k
/PXmqXMTXrUwv9XqDNu/nA1OIj5gSZ6TvhkSVe0lj9RdNkP+y+sUc9BwJsK/Fb3nO7fUF+zM5Il1
505RlDtSRnQltrXxdhmUOXdQkrnuebvGIJ/O5bsMoTqouWI8lrBg6ilcQqf9/ghd40gCCyzKo5yQ
gV/25MsPGxRMXzH2d+HeJ3RVKAWDqR3BSgI4ShSYXBxsX5srehmDgo4bn1xD//d+feebqqT24Mhg
MPsM8bw5REchEQdIC9sRguLMvKzMg02itam7pY1zC1eNtWE9gnM0mEdijP7ElmkTj7m8LPjAErvZ
1mNc5yL12yaGombOdUrenWxtKnqDU3Ldv51ZUd1PgCmbYcI7h0mN91UjJTiXC6AkejNF1bEIMCJZ
MeuCTqJSCvp3qJ0HV9GCO+ARj9YSAK63ojJW+t/Eu4CV/apfelObUJZDxuyK+iueamkJrWQoiCSl
Tc246R9suXO7V+114S8Ngn/5WhbdP/jou8uRyYFDmCUFa5vvGzv6TPnsAn7wuMXhaoZIwsIqTOS1
kHVHTB5mnNl/11nZBIWnWi3YacNKYxiBfp3MTqyn50rL/FvrylcsNnueGYAOJKBfQ4BsoRCbxVsJ
pHu1l/NIzUcHIUhehIV6dwNnHGawNu1fnfDroJ3v+xtIq/+3eVRAc8Yv9B6KOdMZQciUblMl47mc
Eteo81RQ50MOCpt1nBjU6ftghTn9JCd6bB2XqdxrNp4q4AhbKf0WPRSJLC1viByJWhqyy0g/UP1m
I+d2BFJHVQZPDpFcJgNShmtFrS/TA8I4LqEPgTTmeruk0hPR2ap9FyPBG0Xy17Tfq5es2g2/VuUd
D8NRAN24BqGAAh/PZz8vsv/lJwtC85jJiE7Ny1BDHnb15MQB3Qi7OkW1oJbd2gIGyZsq0BCKztAL
XrJcmo8awzdqovBp5AKWsXMM/ZO7Vkyzgb0QMzn1wOPr/EvkaK9pD8SZt2rwDaj+xa7lXeUY8pDN
jE3g2Etck8hT+1oYYETR9wZDHhLVELfG5wVWnCQ9vB+CguNCSHtTbPDb9Bht7pkegM8S5dmwjNWD
Ba0vyJJGHX3CnlsXHzTbzdEllIVtQfZDpKCgOFQT4C4fLnCO8Mxfwn5Fyzn89LeI1QvSgb6HFvd2
uNeIXf3QsG4H3sEhSiKPK1E39S6TgXmzSTGrSa2BQRaXNoaJqg2A84xgmnkKzjEaSWIz9Epwc3e2
BvOKHymvTRLDCFLHjmJeit67MSrFw8xoebYjtoflF345mhK1D21S3V0KDoFGdxuGLH1z+vpQniis
R7FU0G7ECf9HCaoRX8YTwm1uEL8s4ZcQvKX4Wcr6D/AnmYSWFeKmZJ2bT2t/vuvOysLPCTXv7WF8
9pBtLcSpkoOkXDbSGUmJwH0dpIDoAOqN1btASiuh7KnipwlaI/9eBwYNIofl/MpDyzaQnTx7snbF
dRogYr51X0pWL/GIBI7nMaqnDkSMtM7OEZadNFoapuuZxVZQKWOvZ4lJMJJxhJvVsmzpM7jLqIhj
LFEeztnF6j0+tamQ8dmVEvl9Y7Xivu8YOLlNaqqauSds+U1jVY9ObUYmfFU8/kOPpSRzekIheih3
GoWSO3VGl8AjuS5Ftp7emEfb3QPwkhoEnVvdfFxCTYxyTPCZEmts0XWScE51/bCxxxh3umyRxQRN
7mOcbyul/GXbYrnnRxDl2+IUann1vonehSwI8HaJ2uo1k3C4eFr5xOknoAAMQVywXG9cOducsHJI
7tocwRER+URVPyhFfwjTbvHx3zMfVn/LpnEksC+z5jKtoi/7br6qF3OQNE+pzqD0LscK+7eWaTOr
iZKkZdND4DqMxEzlNChNrBhK51J4+UpLRBfO7dN66C1e4fYCqqX/9joWy/6oI9fYnK07xv08C3pV
AJZ1+B9/6/cuFPkyHtaXysuskWSeRkhUignB/ria8YTqwVSroB3Ise3TNcOfgUVKbqZjh42jpUbe
vnxMZf7NgJHdZcVBJztfLEY9ydDSqRtSDAOpxPbu7gNALxwedlWtLY3e+ehK1rqI3BIR1bJJng6c
Kh6qXwNsGBk0Sz16MNiWJRRhOwnR4QEiVsamSnSwbwXmw4qY42TiXfWCKiL9rDhDiycBBK/pOH21
BqJzOFVe9Gvti81mxKXg9D469S1fE1jgdG8rxX0nPOhzoJk39Eprnrcb1uo51vfffj3FTFdJxv7C
YIEPQROwizAqbyJQUowfcd5XdrbDE4YT+w7pU8/Hp2s3CXllo801QYhBAGnNft9dPT8drN8JPfwZ
9PolnTkuiXnnJRKY+vv9pHpQPk8919eI3NNn1F6yc4I2nbmyrdiuYDf8iFIcqcZ5XONKf5ypYOLk
2AyQ3MT8menee32Kd/NI3ebFT4BVp1D6T0kJy+97yJUz83eVOqCNkT1nZt2v0WYzJ9XwnBLhJnNw
MF0Lj0IiMjEs+Y9VY6A4j/LXYZ/YNdQGutK2s0XaeupCMlfssigmtyZQpujVyKs0BlH8BusSXmcH
7xzktve+d0CkazvcYlsY49BLHaCHv6hx9uoEcCmYZiW2VsFEDeQlWhVG57piWQp/R4YobJ0btkEP
rHArZ9DQMwqfynNWVpySeCQ2BXO/NYxUJFLGaJl32RbuEI6JfqCNX/xlbvXDyA0PVsd9cR8aBGxf
utc2MzT3mtRCrqZfX1JW9Rj6T0RcAj+ayp/18FPhbBsg4IVqSVUl/PW0mxLbrAl2IusSBJCaQGIu
qFIZY1oEgRsOR08AFztpoVp853rAVGDL0hrKY2eomJ6HCal0kgDISF4ouGvRVEhfP6mPdllQQbSf
FF1WhItuUSiotdaPI2/62OqaVEkSe9jqYMTD1EsgUgvqVBbFZEsZPFWCYHZmlEi47LVkNyoYTAtm
mAwb+LsAgwojBRPLpiejD7pwpVU9I/xgh2zRLixbIdLuRb7TrtHAyxp18bhsolmcqpcR8Pg6z+yn
ZOC0pzso3PGfiIimFrQp1THLonpWPVCyef4nHmy+bhturASPw0mp1DK1eSHnArdYK1rtYx6ZvFUN
eLZxf/2LVXVAkvl5TOV3J55x3VzePRpS7ZNFF+XP56TECdQAg6JjvZrxlIde+huoePehkMuYjEeh
+xYvjlXtSceZcxfZcN3rMeoMUsjyFIERO+VwI0H77KqgX0zYfa8nMwG4tntzaIX2R3P9NuxAPTI5
fL8pcrRhLqUt9p1J43FUddED6N8LuqaxgOTRNTuqm6DP01K5W3DwedSQBg3fcOIqbMWKV5hSBs+F
r4zqOwJKz1wZelCHLnd4i840mtv7xdR6t1YXnxMfRaW7jO27WDscAXNgO+TTnyI0GkT6HtbZUTfK
b554Z/CxLHy+YU+wYvAUb3bd7XMJCFyBGhAlBlj7+UbKeEo2zb63AJWBqOzZ2ixcqJC6c+OjTszl
RrQrXS05UEqX5KBXJQc7qjY/i2IUAScj1qi/hN/GtxfMOHG5B0+9GBGXQmCcza+lSInRGns0hhqo
L64yIwcAYoi+voSqUMrBPiQp0eUpR9sgxaLKWyEo9DC7TkthKyEDNUZSWy3OqWRCAaiborJ1Hzus
slworj/+jY8kmDwxT9rsXM16nt2aoHoqprOa303j8/qwp7UcByLWYhJuH2PkPL1dR71SA8jN8JSw
Pw9oNs31G0d/IC4t5A2jzDZvSj5oShots5KhEHfn3BQT0457NjWF5lufR2FKtih+AjCrMw91zcAH
FTg6I++/3lD2op3+7CUId07GRJ2pHil8gv41w13kwMKmmRgEC7fsRknoJkopniIdJEeEOnJ2lbkU
on1XkJecVo/vkdSPOGMmfCX8s19O3XVtF6kNbgOS/b7xUAUGVv/dGpooyc9GQqFj2PK27xh4IyrN
5wk9JpwmNX3Pmd4HEhc97ovfC4Cn6cJGJafWOSLNDV+3NDqBP+ATOqW2rbLA1ASrT8cMuniXkE8u
GPIrtMmlCALrmSKImavcvmBYH4AC3cmRSU24p3fNUrWJG+L6YiMWZtWfMbby9c9keZq75JgzE98x
jgFi05IdnlmrOZUJV0YHhy5g2rqKgJBtoApecAXC9DVliJKFo4Au3uKLKH7qsHNQiuhekD5Slbyv
wJa2FGAxoN2oin2NsRddCM6B+9MZyoAubIqXQKAk3XtTrmyLNZ5xpLoz5QqBKeUd8YrkWcL4jcmi
VV6fBwrJ63UH1fziJLPeLrn6b2hqGkmBVxzVWU3AYcHCnbBFd36JBeYe+1lrF8YsFyAI+tzqgqEP
kQ5pJ1hNNJDG8c1kTTFPHGxRt+vdcffVD+h9YmN65HFe1TBj0GKYYXmXpI6Nxbk4Isl9/WWeBsNp
991eWGwt50jBg+PRyJGc52n9GYs1SNwp829M/heC5KgNzkEL9PFbIeZbXBnoccUrucCul52viY+k
t/utd3UOAXFS5pur/+2ekz9tukNOFLjzy5xa7J7SJDFXqVWltEIKO5SPtGgBtmRU8SWHlCG9Ji5j
zyOngnJGrfAMCMYMDgHcXSV/DQofKt/fUPbIyQAhasgDtSuLZIlQGmxjg+/24YLvo/fGpmI9XGZ7
WifxtbdovBZ/abHe9o8hIpdfiZ51Lw38kUblyrm6DQ1G18rUSCOesidSF4GW0JdcBYst0Nk1NkKb
O4ArEe16BlsB1v/OVHDJLhWNm3bOcSnVlKvAdKtV1FOdUVjuPg7jNyPHkeT3AajpXklbRQ075V7M
UvuiHbUVVKFDUoFfD16Q4w7msjiPtsYQ9kFN575Pkxpfp5vFbjci8LkJ64SkMUNF4LQUE7PsTY5K
vAdDOEU8Rw/ylt3VnMyUsqv2tzP2+abCyPAMyrIcG8XS8ZLFmC1FS3TWbMok6jKvSfiqk8kq9bTL
aV6rwqALGC3btcE5qHH5dscjzSx89ILSMii7rgFCeAJAL6iMaA1XeV3rrhMDP6GOpQy/hi+636ht
YrhwQStcBmyo8NqSLVIFjcMFTGr5fqAkMXfqQi532wp7pedQIL+KTVVH/btDo1apJoqMTSvK9dga
KmG66dFO9u7AWCKS8qbDv/YAn/Y5CcuYA/19U2LnwoOXq7INlw207LkzMTX9cxjAqf+gwWv3JvPV
0Ps+DtRf+h8JoywLns2YuQnpW6x9+zd8P4mquxR+B0iN4oRResuDiep3sHDtn6fWvQv+Jxf9W7O1
XF8ftJQXrOwuuUKoeK7I/4wc4qYU5+rCnXO5UZVFjHYN4Gdx9vzxosYLHFI3QwVTAZWkzVlvbzSk
0/vSqw9Z4Ei0yD6g7q1rgiNRXjH703El888xrjEd1i7mo6LapdSLtxrfvxtzPrJOrjPL5yUeDVRw
NjCE6vc81nMqUKOq4iyxVjyCcz/PMPOVg65+CQf8zD4HFhbSRIPc1Bnl6saNtejgucdSvjNZHZGq
UIJrQl1Iv+8V1uQ2y4SU6V+cE/1a1I2Kg2X1rEHUN4g6iSRLh7lt3fdZkP0bdQF3mQ+HOtWFRh55
aG8qxXf3jqOii9VwTHGmysnGkYzuA58Yq24s7ueLvEefqHxDV7/3NnFsBfFjpLQgrQXRPo0NFDUC
arz+0lufv9GrzRUHQc/7HOHJMv327pgdm8mkiCw9eAumvl4hR6HD1GAHoE+M8HYiI/XyWI76BLHP
WeGIGAQ3sEX52AlDQ9YORr67abjyXhOHDp/M+20FrQiQ8+lrGV9BnVoo6vbRg+dIaTq/eoOR3lUn
EGJfHKA0vqMn6KOsKBxoYQMlYovMHqzG2z5L30Pi8WXQDySmghvuY62Y4EaTIeYqfU//YOdR/Akp
Sll0JwRjBH5s3osKeIU8g4s7et0VTt4PVNkO1myLobfb1WQzJAGk3BOfkrWnK68H6JDYcTJpgS8X
tONALVFNztOYQwea1wN7XzaTEfUge+GQfA+ufPBaoSLLznISKx6gxCr/dn0ipTHavMW4KuVHW5t2
zeL+4N9WdhY5bXXhYMaKHIxBpqZcWRrzOz3Gk3Hx8/jfiNIcJA3gjvCiJQdiqn3fZinSommJF6QO
7iA2nySn731OhP3y7j2mwBXPrh8W+NF+XPMGjztnUmCLFFKRte2IW0ufKGj9/QU/ysdeDp6qlKiK
fbIk5SVOhe048jiRfoZItB1iBreoZvKFMqc5uSqSExFkdmlysJMCk3Dd5qf4iJsnOhPvpw9s8k7a
FMCjxBKgGKMUZR4yLbNjRxudT4Kgbmm974TH+Q3G/GQbCMqR8LWFLtAUNSQnSh1+EgBReysjGLP7
QKeuXDogWxPNtW2/0kqWapXlEiasrlUgjK0Kb6qUs0wg3f459Co90CJjFmsRGN4gg9q4W73IP2Ut
h5pNdSlywRvHEt9t95Jte1KvuYYejJbGQbjiTBTtsfc7zdr6E4Bx2Zbtf3vK1s0Cs1MMzkt5ZFKr
7En0I9086jzZ/h2gVjxxv/43jyPKB8oblRaejl3ic3WJBc9L8+e1QnESC1t9fm/esLPH+binGc5W
3mm9k1TrdeqW/+C/5+xyPOLluzTUeXGRzVJnVemvSUBEbHKiNH078YKC3FKA4xrr1VNC8motVkyY
XmFaRl+P9hM2HzUwzdyqCj8ye54ZomyPzuffJ0s8UmUxsXP9goBG1dn0yrqLL+ZML8DqFIfmodIH
Cxv6s+x9/37sVe1a/IBc10PKrC81G0zzCS4JWsrhUp/mTrQdPpbCtdONqjH61NJ1H8thspyDR/3+
QwDx2y3Z9ECfyis2Gee9oeensbBfBRKzbsb+fIn6N3ohtuP4AksawGZeazORcuNOOMbd8BhRjggp
1jKGV8q51Or78YAJc/gjYWloIpP8sAVY/xvB+6t4Slof3XFHsSLWCSn8j1ptNWdYOKZ6QA2uGTRe
PfA7/Ua95Fw/OAdx9e2iIjt/5fsyQjc0dyv7HWAMXSX8jQ4LwHmtjSlXybzumjhTXCCnJBEHbiWS
woErrrhsAq/NXWc0OJpqc92FCdl3ZGCM5Bdui5HgZiAYeN/5I6HH5dI5sjf1zMxjYa5ztCL1KAFy
WhQ9u4UV8k3wcuuTWXU0i0z+7RngsZIGGnGRKSWVJB3C/9nqNqieT7Rk9DxYVaeO+QBiXn0y0FcY
FG+eniFO8Td3tJW+QOjJQO8fLSUk/mgNu4jyL24qcVk3feRJudCRtX4y9qQHetzPl3ec9krhcN/f
eakVaiFHpPwJuIrqHq4r10d3XqviBVMmnkuJ3ySZxx10/m8tXRf0CmIF+U/M7K6Nb73+dMDzPiqI
d8ios+KUOIxCKoe6idDDswhyTu4RKDFQFpj0HTSsniVOCi969zgugp/V6p9ViJqjnq9u/HL9VH6o
V8PNhdVaZqVl+xbh4a8KjogfEpT+FyzcMDR+6rB/bk60H9ySF7gQnX6slWPq3Df/6OZXtDeD+Ef2
kvHPse4/suNZR6FrJ4z2TCOeT3cHKp5UDwdCsht4zoEY+i/v9lr934aJCw6OAwrtM3UgEk0g9lcD
cWFyE2wj9YADwPVXr3V0x0rQR1oi8Dk3ygwpSLpkAFUlYXeZYuYrkrNcrMfuPUK1XGzY+UEInlkT
T4SB6KaYUOU37zdB0LWRnsdE+m/8yajZlyHbogsN1D1j7eTxj+gG2OubocqpcnQZlRgBAMIfdBYs
wggffFbd0JXbSFxWA0xItMhXfJ2VhvN760vnUvwhSxk9wT4Qxcf5QE7hCMQXuKcQsj/qZI81adbc
kfRpuXxawQe4kcp/2le/wfoYy+rYKE4xvygmpE1StZN4lMWbQcCelicNS1EjyXQSY9BizmSfNeOJ
Z3gKMZLym0Ve/Ae6A+J0ymcE5dtrhMlvPEGcPj1bMu76TcBw3Xm/wFL49RwYZTZ3FPhowWjS4RA3
NAwkbOzEGLKI+2KFYagYO+o+uRQKM+onrq89hzRl8UQ8pWtswJrBit3UOhLls/8XmApamkqktT0l
JrrI3FWXEmendjes4K5oQZLYPBDxrQ+b7l1tEgjy7PclBTN+c2B7NsSpog+sEOpRBDY0mxl5Zrb9
utWG6DsCV7igJdCBe5F2v6czUGV2xmg0rr89zjchdNURp5EUF8sc+wyXh/OrRNXpKscRlHA2QvBk
oHuHFATQTaF/sOPuiniYr9dnAemOLbuSauiIvbsn0xymOltvBtTRuMtBCpcctRmf+2m9knHYYzBI
4rblKcuQGIUb/A2YBQDItFwCID2z6mX0Yb7cbrJRR+572jMaaMdDngLzhl5ApKjAZZ7WE+xBAlWT
ogHqSWYZmrKXodCEYH/UTPtVcDLvZAt1nx+YpVjlpsP+DMTnkzgnpNGcUQ21IzxwhkAqsIYP6ASJ
9zYJ2cb1DwAI3qlkxZW6SeHMaEyay+cqfkaRs3m38WzJzo+l1/d6V566AlR55s/G3YPYntPkcsOk
xWSsme/WmObv6lMnz0xYvrrWwNhFKYZ5E5laUzQmQ1wwPLIV68ocB32qqBA8Ec+CwPYJYL0z3em9
BGlg5j+cUFlVDH+kQ/PEqa2AVqDoRl9fbx+9Io2mb7JrAVrBHbs5yDxa6wMdciebLFm1ph7Nz3XY
LQHtZAaYtnh/KyG7dDUbKKJKdkcpFl+5zILXU6eaZGzHAbywHPLP7rQEGBRJP3TsUpKj0z/9zXjA
gZGTbgTbdzB+ZzPaLgSKS20+pd2kybcXlZYgY8lu+ZlboFfjBRKsQRRtFeVWfcLOdCoMUa0x2i6G
HLIEENN3YbxdDp0mRYgxBIKUy8lEaLZKOtB/Fg35snkGt9YnHyfQ1EwscaRIufEyhlb/4y+TL78x
OUyZlnhsPISRxrreO+x2yqr2i1vcZPuZduZyGK5vPOpuKtFzvLRqcCvtKZHbVP5abk4bFua6LYfr
Yk6rU3q0AV6VEuFT4KsaRah1GZIEekkjsDzcFW4UoIaV8mefgRaqI/WH5DCrDijWPCpZ4fz78RLE
B1htFI5CuXw9vysZbWp0TMkmgDF1RStTQd2bP4ZbVEXdue/kB7b07z1YhwtFxRlx3TZ01DEGOB9K
cbfXE0cx8kklyNixhYXIAWYtoVG5PnigViiUaVD9V+9Qzop5pu4/nOqCWjuioyh99Izh1RKeAlj8
0QyoJBL9D4Ym8KFtP6N/pblVzcpC47RGvMqyOoFjUFNTQZv7IRDBmtDsUGaQ3pR7AEGtJPUwpKPw
eoBAaGf/U2MEOqPwRnMjZiCE9emLhggqR93Sv/Y15U1s9wa1ajQKtqyWbHbjO0UZNh1AGo2v4i4i
IWXS6U+jHUuZjqfPvwmoF3mJQENHrC8PlEX0i/VzTUKtELyHeMB8O6GxAYJrAbQM33yoHX/EadH5
KeLNB2pkCnSawGVf7G8jjH/4stIj68axlBXUowwMWtRdtNEZIXDwpd5mk6hHDW7jCzBOi6Kvl36B
1XOim6CEaBFZ/z4HRoIn1iio2uQEhO/jSejmiFckChRAC1gWe3Z7vXTEhI+Hi99L9Fm0UTUA8XsC
Edn80DJV+ENGo7CtUiIOxZmK8MYF5cYBh9+B8suRq4TZdxqedbFqCqmU71VenYRk5sSp+bmjr0Iw
g3PGPaoSv/gOf0hGvUHVn7ZA7rFgHLpxttgs3yxZ/aVfy3Hlk6Laixp58sib7ZKvRvsXRK4E9o5o
8UX5OtAPsWb+GHZsTTTAwZ+SshgZNrEP3zs9cID9obDI8i5lWetPSNEVmAw/UZUyUheeYVsBsvXv
X5b+iDCNcpayctAqXGldiSNx51NFzd5Qujsb8eOfhzWgyEpeyk/tptmGAwNbHPLvkosbqbA/FFA5
EwqjNsyeahJnMLGc0meglHGs9EcjNg4oBI3mwrdMuqyGvwByRqyG+PmJEggXEaTTchpKMl3nRLJA
Cbu6l2VbYc5LqjFJyHwVD7wlkfEbALIlwPrff/Kuyp0M92mk24U6COS22vTTiXmTCvVmAwxuSppK
tV5S1Up3E8C48qqBvGv76IuDNDBa3Q2jLnNnbq8h144O7a7T5EglifmDIdYb4YHWkJcdHH7+rspB
CAlTrFot1V/vaTGx+uOZ6PD3OW8hyHr4pRr6MOVt4e0Cu3EtwAGGMkiInXxUXVJ0q9jk1ToqR6dV
Giw+ZIEUOr2ADAYJf+l1WPnjYgxgySjsCL1Bd6BrexNz4nnB4w1slEw+TBzZpz+4G7QB5ZGGoaHr
I6sM/5S0E6Re7vje5027pp0miC8nh87o14+VpLDqYjGpaetM+dHRwkWmqtZl3WurcSgCv6UuISdp
Qd9RvlVwP5npsl5OSO2EWha/kH2EHPyD613Bad/q6YrRFgK1p9BxI2wKQxbubP63khX3Ccokvhkx
4SflIpZqT5ASbwjHImuMEwy98E+jafGyRlibtskXzec6HNe8OonBaRFromdPf0SqUKywrUzIzmZq
g1KbnOV2U+4sv7ULIys8GeW+jtQumRunnN84b6w+SOBsmqiTp4kaCtKbQ3xyUUVEfOWmJIMU1N7P
B5DJY2u+ZhqSxqgSvZVSLZOVoQIEHZQOi3ayUCWl/5jQxg7BgR5Kgg/lfoPqne111Jtb9EtssRya
Q43Xn/ylnIn1G8b6WxStWRV8TTojIQvDsjRrbxoijWVIRQIVzZQeolCmSckqXoMRSBea+oeYhPdx
i8ygyZ/16ILGYpWa40SdqCFtl5OPOFBnfZRKkc/ICZE1kV/B7aBrxubFUiC0tI48ECoVUOuNfRmN
FIx71H/iA92lYnvhl9n+bKWW+gunoB9HXs30IqcFJ5Y6zSL5UFvWbCeDNXUA7dVYEkexuTmQC6vL
4JfvWJRZ34hTFWijPK1j/R3LDnYZrlOWyWtR5B3Wozr0njEhMjA7slWyA76QiA5rK/TlIZmNTlrM
ru+cyOMG9H1WWVnxupG+lrHPfPOnBr+Cnm12vDUUm4Lhh5jrcNEPg9thjt2jPeEyST+LaGg4JjI/
kWXLOLyqPRiDi5ZMW8RDe5qt9zHvTklkdk9UalmdWmXJDJOmP30Pg/OsSKofnUzqc8uTwlH3ilvM
FjgAVFZSznL6VJAQomV0SxK+TZg/EZhN6wLuVsqCUNsz4sgifMXxnRdWbOVu0k+GumiJ7tBBUPLt
2yROWfQ7w8nxOgPtvBXh57pMMEFuZ5IgtSBDyzJYlBpQ72NnayV/D+iZjNsjYy8QlrKwM3vWBl3v
SNzwIWkjC04PPGu49lcL/6i7dvkFPaNDWCbjUU+OghY7QTT0kugKd2slqkEfLMcfCB93BOTYQ/E7
ERRFqnZkUI3NEKtqsyAVaJAFhz5HoeyLTcpn8zYaBr5y1EJJaovmkS/TH2i3mWx5BY2GlN1NVw2Z
9TKABY3scDypDclU+7qrZ/sYMNtlFhZxYknrWctIVFvy2hsWOvmkMHunHaatXtQVvP7NdEWCdKej
23sczQLHZEHY3GgwFXFEjiVynAmtq78u60DVEmOehaBKcoFDMNF3oDjx5GFpH9/X/5jb1b4Cfclw
S1CKWW8TNAbrak/H+9Ojjl09nLczHD44HgJNBxR8w0BP50IGOD5bBa3iKLgXksgcg9sAyTAhJB4L
kVa87EHjuELzAUaj76L/nvmUt2vcJbr0GKnH1v8C6qcEhZxtFStvJkyKGcbiNqwzY9epx8PqXkSZ
vPZZZWBEQ25oHVC0pHJSlgXooiGIZ2zYsx/hyspaCGAuTQYSiZeO9k2T6WjaRuqyuhcgF5g2rwVR
ZeK9i1ysAjysKIaA1f74iJ5i4kIWyhyKQCiWco8LpT1zBUq8oYmx8Zt0kcaNfQxCddBnrsvxnIpd
hwBRb8KIkckasRUSpbrZfn+v9vxGh5VNK1kDF5kCz0ezB2dJFMyuI+xNpfrLElOGQu7i2RT0kofM
Dg2mIeREp8Oe3xXCirD2FMEIF0UpB7Uu1HK91Q34zOUFD8aUjJf2mCKya3XlN0tjAlGUii65xQBK
Euz+1E4xAF5jtuxwlzSX7qgjHWNTbpmQqhojEANgT8RuYnbwjkjqFdn4k4T4N+Am9ma3BMKIbogr
etwsG1N9xhkOKH4/ZjyoYSzKmCWMJ99Q684pCPrLn0Yn8zJhcaIdWk+f0IjxXQir+c9YTz3QaFuH
T3BgP8ByHUs6NIYwJkJ92UoNH1gtuNjuQ4BdyAVZw9BEQvavyLm0R+PYMM6BI+C9/eMbVK+QwKF4
3lvKb02JhWzsV4lzO02KoRB0FZqgr/4Q/0VWG9c7UnflPmAM/70Qb/bZyOH9fidFcRwxxjwPIr7E
rIpd50lPdNKd+MqpZ++EHN3LEvL/qDeNQ04crIXbQzue7YWZ0DAkMRoXvKTIW92nw18xOtODtBjK
27LWVrOf9SgBwAWU/m9YGLww4TLJ1W6o6s7XeiMvCrCE5RFbA9liUVcv5QjCBUHkTSCgJBOKqQss
VWs=
`pragma protect end_protected
