
module niosvprocessor (
	clk_clk);	

	input		clk_clk;
endmodule
