`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H3t1c41yF9tn673d+21aDVNQF5dKHtqSVCkQrRl0oK1C48Tl6sKwBqdEXpLomqgh
/2Qxi+ZIsmXfDG6nbAJrFh3WQdOm/E8r3OojN5t4DElGM4PF4S/65j9+N4f6nIaS
oUfgYGCnUdk/0AgOQ2fsyyqtDMXR99lD812o4qEROjw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
mvX6OU9QcKjT2UbA9k2uI+X73O1kI0MJXTT+Sm/DJNGkKgJx18gVkqnOwL/GcGa2
w5SRcQxMLM68teAZzNzhLN/ZNklhDtU24DPOLJU8DybPlHWJBVmQfQQ8g8xDcuOC
q5WN9IsNjOQNsJbRrKMTLWddH/Gb8aPKdjR7wu6Boft+jBu27hd9Qn6Of/vdO1Y0
1xozJtqGaDLSEwLY1WKHacHWhWzrhTu8k3yjhk90+BgEbAeQ4RHvsxs512EutmQy
mcpi5kjVlauGgEYkHRc3LNHeZOSiYJ53/iC93FRjz7pt1qb5S0/aAUdSdbrEhARf
52y74dhEEtsZuoMWfcpXzg05kZa0u/8wfUotc0DupLcR8N6Dy2NWQbZmqwmCrj+G
2vcD/a2cD8S6RiHjh6zlD2TiVzicPwnYgBlIl/W0RQO7W+FPxHpPXiF8HVAb9nAM
ea1gAfOA228S/hl9r8PGiscdpGiC1bLqP4iQ9bW9b4qNbwePZiASKkUpinoAwNEU
ps2b78HDZqJQYFYSJ0r5BtLQQmaYgTHXGJbi2uELBvn8FbOTENhdbeQHUBsepien
S/U9D9rEI9zU6ZikBSJif3fZOS07DGeqVT6/6cl071/tZRBQAOPeqt/Wb/96Se/r
5gEZvmKFYgp54i76RhIXGko0p/h5Mv83u/m9OYr5cR4V6KwXELSBmjqt7ozV/7jS
1Mq5yZvQiGxY2FfM81wcqX8HdIrKrG6ygigpMtv30kz6qnpBUKr3IwVvbp6N9RCW
juXnrjTI5VlU7jWwApMwSkJl6mgi/liu+oYa7HhC4/RneHb6rO6mtNDjgSTauLL0
sxYT26k22iGqM9MhGO338/hFQOKAy0DIwRyfWP7m5NH7hcECrGL5ObNzjPcu6opv
ajGI+aDIRqz2dDw69sKMJ2mc5CEEoxtD4BjAZZilhZxQc75bPo2mmn3VZRz+qync
sFubsj4KQE/joo8GUh3nNbTb4FpJtwOUK8lryZPP6VXi8Xm6CqqWOAuGEoP+7TZJ
y+94z9fT+k+QUpSFtPQYqMT3FBAXng93S0MUpYScmFwvKvVTMnP1mfH1ue67rBQW
SZyuSa3J+MXK5A0v4wy0rMfPgLwIwRPJy1IOtffNj1mDDTFS/9WWEqTRo4Y6WnYO
FMxZMj0RcSHkMLH9vOFuewt5t5JIL4t2q5I38tqejJrTtg4A+3i5e6OMtHBKd3yE
KE3aoZdnXQKrQhOwvFL03g+tt4KBUkJ1Gn/ScN+PI6QHUBXU6UdcqzsBqZlLnDLn
msftfEtNeOiV5NzqwHHe3JQLVGZbQIwsBmM7TsO4EYFXHFxzmiGlE4VXaO1Ni+sE
e/O6TRpxNfUSWOKSx+/nZl7Snwac2eqsCXAsiNyoNsCmWxU538gM0mK9YtO8EPex
fPIKEqjzZKwFW1VThQFi3YA9RxQKWGwRfxBg3HZ3nEXALiPiTXvDquej/z6OYTX6
BDetcBX5AFvMC2h0tNbrtRWrbhhU198pCBd0FDuT5pxbGgZubGkupooJha2/MNvC
4BYwsXwQUBquevhZdJL58ugyvvOZaX+4TwRDFRBXd4O1SH7QebUqOQ+0VvuT2MfD
+UNYrgmxCVf74Z4rUT5Ca3rUv0yLkd75RK3VnPnYWOvlBPBs8ZIS7dH40QzmAdXp
28VCOwvmLzwQklyl4VmRxbUOaVDXMvKgOQ2BtGaCZEmubQD9d9fZ9PIxfRmUftA7
x2mPqt8JyAYpr5taHYOrIkQyfB9KztWYcnxVCQp3C/iEIsklMa9fbcVpOBQvcOwv
eIlAAPjuUobnxbV/hMm0UY1R/fhdrvAIBHqpLg/k1GUqgbUZq4H2Ivp461BNwyhW
5CDavtv6uQeEwK7Xvz4oou3aybLYNMmk0jlpkxgSL9CGFVXEAeaTg3FKgd3uVvbi
yP8IoPVYG72ZymR8xjxlLZ+ZDh/QjJmxAtVm0xd1gEyZDO1goyE5ycqHaItSCXMA
KruH9oF7rfMcLh+zMZGdubRE59PCO81JO6+rr7ce6SZ4FBrquJ6NtGIAn4PwhCzP
GO/nzx3oU77FCn3NW45hFn7nq/jIXJgfM4ALFwr2OVOB3mgP5JVo0opRoXUZudii
KVvWAd+ML8q6zYgWxyza50GOLz54jb1v2R4ck6YmEqmNUsJvcDam32b6IXaJHIhO
POa+RYLqtSQ/MkTmcugkCgTV2JCEDTXYYcBtDOmiQA5DbGO1Qa4GZLMfgeYr5ua/
U4v7HrVBGN4NU5PgSE7XUfef3SpGSZc6Skt5nnW7qrZtzq9v5tu8AdyaU3sKqgX1
tlp27azw6ivs9bubPaitz6vszZCuYHxR9ItpVvIRUUeXa+Ejv5gYRZBQfuj0Or0X
SN+r1eMfF5QmR/EcD7Hdy+MMNWtibcJxIWsjr6jQC/SdhK+o+Gl6AKeIp6b8Wj6D
Xn+0fghTCMx8sALAsBKmzuqCX7InCRGTdwQ/fbi35FzHo9+EoY+AID7hEe5iaPVD
RjChc3VoBW2KE4Txh5IgY17Cm8/PeFQ9SzVWvkkVTNBT11jG1cUOW6giFpI7TS/q
BpuT5aw7Tk1z3R5//50vcjjeC0L7BhgTkDRa3ocWdYW7HmSl1Mxqzhii/3syABEV
2EMPJILySXjl58yPna9ZeLXjWQ+Y8mXQXygmKDbyT45Bo+a3s2ni0fB0RjqusSxA
iiZw6OIPyB9sga0Nshs3CZ4OHcaqrwkAZfVVWTz8H4/nLLSq5GmBkMHQf0vtFsQF
kncs2cqfWNCb1fAHOXskqzjZaAvdtV1TfFmTV3+L9wBGD8W6PKLEFtuDbffNhWj4
IlEtaYvkwEdhkj6iLbOCvxq2vs2rBgOEPz4tRI5yy0Vb77ibXH4GH7PuCOwk8uJ+
t9fKbau5rktbZEI8A0+ZlAwS+gl31KOcC7gABUiBxltPbYP5VqMhlA/JaypQz1nL
AyhsDGFIgB8wABu6/zCoDXGXJ5O0lvbki0digrDP9u0=
`pragma protect end_protected
