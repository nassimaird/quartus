`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ciz/pKamwFFbyhYcJdWEPBw+FVPgNigxTOMJikFDKbv6ArLXiaI9EloQ6iiuGPaS
nXfGF0CFcbFG3kEovEEwqvpqa6rSkHO7jK8kWk2untHIccHi6mN5m7TqHioM4tRA
GERfM7zYL8vxxqb3I30noqHuNyr3qIBIM+++Zr6yJwQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10224)
o1aqzAwKIG/almgCFre1xgkFJZqYADXkvbmAME4OWEbt3geZUYg0LiBCEP8NRjP2
xgAme1Q3kjPnVmfmrSRqdMy+A9i4pOH03nzNBmA9RZQd3UHi1NAtoGcvH9X3HUWM
fXe07Zb0AOAdAngPAxwYvr/iciXQYdzXsI5a6cfsOJv3S4QwMKrqGFhbH4Wq6MFe
BO03MPZZEC3CaciA5/8JAStEbltBsTq++qdb8K3pvtxpW9L8fKSNdD+ERUWBv3Kj
s2NkC0TZShFzRENiau8X0vvpyoLpCr0I6CHgDv321oVbNNQKvSdOdBiJT1lTqyvX
Hv2EyesYKt9UJo+b+EnXv13FdRPEb1ViHGwX/NgXFye3DvpD7nTZRG8too4DisZk
MfytjLWD8hJYq3H9hkJQG5n8/7JQnLjC9kM5Ti4igEP5b38P+3Hh7BkAzsKPJfCE
4M5pH89Q7Ip/LhZ62kwHQUsHWDZk6NgSYIjzbAvvUS06t2zOptkxVbS2sxJMrjCk
Weeog8x6zk2Ol3WfAVVT+uXWX2Ndjwfb+f6Azj1wC6ZPNJTrndxvHf7382d/IHN2
s9H6bfAvFWb6tEYpmAj8dA4a11MRoDgHUd3d5rzIxFvyk1jXstCVZOinbe2HY1zq
Or7BNlEy/GUvJCSE3pkZT7Np7LErrszNUnQIcmsdA5K0amxXeDaDwAt7tPW0q9Ap
qqRUXAXRss88G7J6yEbEY20zkenKiaW2KP3vmOe7lswXk7nNd1JxkAXIIjnRD1Qd
3uSXMrosGlAgaCDVZI3umRzKJMQfHDo0yVJTohl3wLa+Es0XCYiSgckj6ScM5yG7
8fB3zPj+F4UkBWY3MN8jnfyslDIDooiCHUIlsufwNcaTOawzOIfZB7aTDaXX+Ql4
Hhxgs6lyOKrteAXIgJuyp8yY8tZTO/RLFIoruNuKe//ocTrr3ufvLj8fsTOQ9vcj
cX0Eyqem0tO0NKJrgEvayLAc6RlnpOMk1Pau5LI/hrzsV0UeJsB4nwkxz7Au6XJz
Y2ENB+1fyAfxA4BLQDtE4llFflT7GvW1yXjQRPSztsxXihFI4SrciJCAhpvdbo2D
fvg1MYMxSfjsKsDdkkigx2k38ar0kDck2M3PX+1x5JoKueGzFgxpVqyPdfuKCvBO
rGRB1aHtRv3xHBXavH4HKrY0dEel/1kyPHILzhiUlC+4FVJM3QmrVJ+VH50ClJ9z
VSxOcxltAAaISruO8ElBYQnPbXXMiAqSUBVWAMK+7qRKPsdIgUEYBjFer/JzRjZU
jryMqDGEXYAr8ULRq4U2KEFhL1ODRGpY7OwwCZVd0i2nbK7GSbfSh36nPC+xqJ3/
gAF/WHKx9oh/45i81onavgfakQIiU77y3VTbq1yXvzXX+W1FZwagLP5QkgIfPAaO
ghWEY5QH+TkI6WKM3Ae0Y42n09y6aIbSTfC2G1xYmDKXo8G8o/wWfnmEok96Soc1
ab6yl+PUaxJIKfbiYycgqMYWU36Yq2slz/r/reaIgUwqucNbup5vIOn4ASh/XR4g
BW7xGYthxQQBOUPxKHkDEWoELs4dBaRdxfpsU3m0fe/RXRMsvyonLxhRSwIcsjWO
mHtdwesLT3eO/RbhDUfNf3uBFImgGpy1TicwuOBwCBSIKVXeoz1NcaqISvIptSQx
Ou3wR/tMx2hghKdwUIndUYiRmgmI8pZyDe5N3c/7L1Db/c72L8iz1SkCAimMxtAd
ZvQfqaIlHgx3JTYdezU8HAo8MWXhSyUjcpO4JfL3U1m0QRUALGRGG3/cKRDPHxSl
M75rZUVeNT8BZ2d9x0CB4aV4CSY8Nl8tHKFKam6AYP73i8wtb1ISo5ruPW1nKE7j
IcjbcXz20aLOQ4cU5uwESXrG4RPbcZol5TO5R0NhL5A4SbNDibUYcxDdFTa8PDDA
I8mW6pqLm89SVYimfrsYeTNVkAvA/6xxCvHco+onSMfRExxNOf4iKc2ym8XW4Bpd
2TVJE7GSaaSIJmPbSjBCV9xRBfpTjxIL9jxHUUs6iT+vduirT0Dch5vnLyQuvkRs
HJLZ2dCM0JQnUpKvei0WTPU3fJH2nv/Zm3CYHZUwQxdRhxFQnlGe6ARWwVQcZwHo
NZZJ4jG2RNNRdfYb7cLx0KOV/nfz6l+5cC/HJJo+1E+Nk9yKjF0QnZuiZKut09ZC
b8Rh/NXVd9y9c10AYWas6pR8D3Q9BNfPCBpiBYU+qcB+uIyG8lzZte20NTrn5SNP
+9wFhq1LZnObNglX86HaLamxwyzY9RgE4GELcnGufc3HGhrW2/l4yNakN41+wCFL
SJsQrp7nbjKKJkrMst5QcISd2J11AYXZn3rwoYWqipuMvrKx4xD7DxJI8ZXEXn41
o2MjYMyzvsdNAP7i/aV8KLnzx7gof3MH62fZ0G8MG57FDXQfmazZDOyRcYsnxGHI
bfKt11tIe3UDjulkpqDq7NK+01NJb+Uvmy7llOJbDybT9gbmcrdn971+N304qBEF
uxnRTB4k0SwRndTHZzUQiARE5fmmluvC3jCRJcJT8ZcfN6y9TX6uS8rq3AwP22RG
qndotbR+e+Q65UR945nYy/4kjR0mjUIj4dCjMT/S9kXqtHWZaA+hg91EMfIxi5wD
W0CMclPs7HPiyCD7adIHlCsv9yHdnRfahzc16YI7WNbhJCyPigF5ReKpEe+pFXfg
zmuAgeg96HxoF3mTs/EjhgkwF2bjHZvV58ApBokkWKpB0hyM8fO1bcfNUjrNor7D
e/7NvU9akliRHTTkiAfcidwgL/b5EKx++CcUNqLccqRTb4XBGytvitt3M0Taf4gG
a0TV5YFvq3EQoxTfD7Ksy/xEcLEwioNX7AzsQH6Dy4l5nhtgjclh2Xh7BAeUydHL
sfN67CU4Hp4f/sp6DXDtiOJwCxqRJM/on4Gxa+vqlfXWnHqrZ/NJZZKjkwySeUXZ
Ad896n+S0HHjus5gpl+Aq4unvEpqB/NKa3bRh8KhCXOUuhKzUBgiGuk2qcZciBFU
KfBuS6LxZ86Et3j21+IYZDWzznS3NMWCjmES58a9+k6crL4tLmQdSrzw8fiG262E
vDQBhEKcsGlo3Wk/QmHIAijpb5JWHIgwkTfzPeS5GO2Y0zpBbLzxmLxhykKYYckB
87zYEIWoL6EcIIAnmTKOZkeLDYxJ/Hv+NHkg/tGphuxQz92RYCKc1DRppFcnDOMB
31dUQmmdbk3JrDiiN61/TURsxsOY0QjN9Y9REWQjXVfIfmx3Bqcxt0xV6KN5hgmD
zn0EuI8SxObxef7YNKziJ2hSruB84k9JysejUiHFpcXWtLYQ1lvp8AyzKfF9Bfsq
i3b/clQkcmPPlsM4IxucOvlIIJgb7vwBckPleEWrNHPOKZh1aVnSxiiwpWwFSpxY
xWLW5l0l+SFbBK67gHR2T737BqPcKglXWETzl6PG2bz3Hk110thPDOSaihI5LvNn
J8rWiBAUZ2AqU4cEKZtvt0VMj4Jbo21SyvFUNsZpu1HJp66B/5RQqL91zPX32h6U
N5KOrvjHQXwaEK8V5Binbv0B9eMpyeuvA2VD2b6t2RsA1Hnglq5yFsNzjYEbwk+d
49YjlegI5HhKYR1ad1DhmLHLWLVJLhBOuuLrDLNBXI6ymcL9IXipmsXtoRGWt7aP
jbKjsX1n1hCHGywhKEDgifXJ72ZvNe5qh/q8IlOvZu7G7zXAl93LpUMNE3cdawHq
6fIrmyl+VX7WbeznHzW0ve1KFZj4JWRC82/99AONIEXvc3EUaJMizbl0SvpgGKSl
VaMEseDisG6Ad0PJZFjj90P/AC32lZCp8skj49YvGnN208GJDInk4lM3uFVGMndn
aTz18Letkjyj+5iaNGbi1o4+eORYbON0APD/dvidW56BLqs+zQ17karJ5T8rTRhF
ff2sGg5SlIkTjHVeGNwI6xvT7ztXXGYA8w+B60n5nZSTPglWo0Al1rop07+seFOk
UGZTaVHiVestVSovbAEzB3S4ss+zcGbc8lynVEaC0x/oQEEShQO1WE4NbY1BfysT
hM6OohdpqOSBA5UmRlSXXarVxcNITupjTHQiszHh96+lOQaU9TbxWPkp/qxsWvsx
w+7dGznEnaD6z5NKT7mdj+YC6X6HsM5aoTwTx5bXxLZl8lZvgl4Tv+SmHPlJr72X
gtVh+338buA+o6RwRBKyHg6lv3zoyG1W4nwAjztL/nHGig+nJfo97E3NAYUJ6GJM
LtsqTJzYYYDPKWA3EivpVaMBTntUTWBWyQvnD/AUZfJ4kNUoFsm59kd0CdPbceSy
s3CPIeJAfG6fMq+2uo7MhYdstwoRUE0jvyiKOtfEOF08bkZ72De06LrCv465HRdv
zWbqw9U1DM8ZoQ1r6sPlT3YX7pJdsMdVeEYbZi/W0dtAM7OjWDPxNpWyPRvUP3YS
yogz5JIPBw5B+o1GCXp/AG46WFZxeG5BnnHcl1iM+UQzVdcExWhEX8SYZoqAU1Bg
hRfidimv/Pp5+Cfm/EQxYgQDEYY5o0E8UyjQgfUcnv2fRnR5uHhyHF3JbiyDbRop
eP71nkHAMgiPYuwjuPnfQQFJYc3W5GQbSq3wWvAYjzcK8WZgKcB97tby63xc0r9V
EbiVOnGAhxC1FBCQEBuRBE8iyr2ufl8mK0n2Q5x6Z6M1peNahaVi895S4nBwF0a5
4sHMEG3X1K/XKtHzNm6iGg+8f3RUzAkNPQGrZ3Lc4jlBSM+KfRzVSMWL4f6DdXyZ
fH0bPIPqf5sRGpFaBhRbXxgWrfqHN/UJU+wShLBtvgJZUQCHMy04eC5Jcv8c1HvT
ndLNsoOwc3T6z+08oFh1Al62/7im3ip1aWy8yGoYmD6qelJVQfNkzx+excblneOc
YojiJqIj+42M8cH7JCOtLmgQZHyDdJtOtmuQIgOFoH8bNIFuROYUpB9H/ZG1LkRO
bhwbGMzsjsA9e7aakCWocuI0+D+jT2f34nd4Z2q/Cr1QYQgJmHXJulXXBYJmM+pG
3/v2KjFo4ng+SoJyncHGaCFikmiyVQtyNfwpSH0IZJqxKaJsxa6r5tYiQRsvQAiC
vsxUrLnx/VbJ+zqkQqlaiNpnlvLUUpvAR+ppHSFQ7sXE/qoxUV1uSz2gTfW9+6le
jugjLotGUBiXvHU3A2sjSTnvNZMJHZZLL+11iFKOYcN1yLzxIfWtaYRgsU6ykTvo
+PivaC+wvKvrz7LAGmnfIcGRWQ50vHsM5JaPM/y9cqlJtiEg7j5z4IyNstGZeq36
cK/L1z9NyZ2P2Tp6qcKK62a+J1WGq6K2WGPMMaVPLQaYzkSHI+lV0xHFkBcIzXx6
q1Pd3Itg+/+Lt1B6EzrNtX4pp7ojgCqtFmyROa49a7GV9FBnd1+1jLWWHUEsVWHe
9lLE8OEqeovBwXfEWkc/rWLMtHGyUVC5Oo88AQq47eNIHV93GbUOsb064fDxcL5G
SuHE4b5xUaABRxSEZlwopskq62lTRxoiM1sV5DGsRYpUSuvcxiWr0AcE8hfEo4iw
MfWSKXwz7t3Oe6rbR4DqUVbZKMyZTV48L1zr7eGrMovevay7h+ydQTaepgNByNWX
MM6qH/5ZrJC3dL4IQrXhnMYADlpNKGVC5uGesq84sXPiKCmrNQ0RrVVe+8Ac0yDB
G72JIWOsakRbyLeV/EDUYR2U9Ee+5DAv7u2x3hxajTnI/HjewpWPcFBmyftCuxx0
O2MplQmjl/WfIYV4xbZ94GTJf2Lk8yUJxrhtkpVNUx8NNXhb0LT0XaZnM160nMbV
z+Hkq136S7f0kMVwK1LMOdJiP3MQ4gv05Z7LL++gsxxEj9U/Cx65AxU5cBt6FrEr
EVq5Zo/RvTwpjgi7UeQKM5Z4MUQ5V+F7iThEGnYXbkTSt+/Hw5ro5SeU75HpTgV4
4ONwty1uN81t0MQgSxwXEI8zbYd9mNwO6dePKE7+bp+xgrsDrFtpeuWAMne9F538
rM9h8cfrD1Ne/7ccXNxuoWVilUbOCOJQBHd011dGwhrncy2LRL5dzl1gMD1SfzeD
PMX+Nd4g8X8n3up2RvM00e01VSlrIpiaUepd7bdiRb/apBvGs/mZYXkko/sZIuOi
Sg9WWPeczIDCXJ2NDnWYCZsBt9eBL7mJ/HJw8cGH1FV2XQOj44v1aic7upHG2COy
Fd15rFa/sJbDoH7d9OLNJuWLOIKvimJ5SpJMt21caKWSVfWxgjvWaHEeY9o5EcLT
sOluMgT/5bl9m60ZMuqSFXSLE4paeyt1CRdtlvzUttl13RiBMUl7PmZopxTLofq3
YlsIEVnlXW1Pgu6inqFjbIbWG7Tx+D5V6Leco/TUHqJVJWVMQTi4816Uzgo2W3lP
/nN8eaZk0WLMImBAyB3EhX7MQ6T21QJDNVyDTHZ23/ofY5Q+AGuripDICVWCNbRC
8U6Tpn5QyhsznpXNF8PJWh/7h5lCQMXmFk9kfFzzU9nMH7iC9n45oL7IoyRWn8Gm
VimDQ9yaTVs/UMb/XhdpFray3K110s0Ffwzr/1JWi9A6H5FF3/V0BpQIUFVeYAHS
K7ngVphK6UCVGY8LgDeiH9i3T1D8X8Ms3rLgFUrbbBO4+Nmf2oClA66yGfT7G1n5
2Q0qDmKAf+569T+oZYLCo78cSwEqInCtJbfvN9nmHpCiSUKyeU1EAjY/CZpErGL/
FMJiTMsMVtjb2IkocDNu+mZgWcTDQdpHvlmHGvOc7tAo1vv2jDwtLcOhKmQqnAw4
mUL0FWISHwlNbJZ93ZG0yU86Dj6qoEZzgfUdpq2LSBj/DTPC6zECEcYMn2dA7paQ
1AE0jtRSYY964C6jnEmccPYnHG98/BxAWnlllaNTuRekQKh5XIOlv4k6hzzrb6fe
fhY5RXzdANJMsCh6gWstC6UqFCIjcGfUxw/SCHkWvtVPhkLTv3DOZ8NRNH1dC9gw
otm8ynJu192ujm6IdxMb+mTkiOLB8An1xorJtTVRKxwFbRq1VwSjtvAMIxPPIAJK
a71VUMxajopJ9ZVMrs05uKH9b8Ye0G/oHatYB4Z8s8fATa3mKXqq0Nx2mmNazxm+
lQ+5Q6m50GjBlbeK8neyGSugEjBPOjYGjK2fgQYK+z8u62eL5eDewkw26VULLF5c
kBnG/VpzjYD6/PSl/3cnJ5tfHQ4SK2g28HUoXV0R5PRIRlRVAYckgKPY/gG+1JPK
BqQr6d/qO2bvKXfeYwYbU9kIB1mSehjaWgP4arLmYLiabhHwlM4bTp9CqICU3y5r
2LuxvDuqoncQLrY6l3fsdvSMo0Vyy8VVTYZdTr8bjlv7lmKO1PZmxl+6fFVEycS1
Rxx/sP4tp+txtvPO+PMU/6m+JyO4q0Lhm2yX7xoLKWZFA0Z1QaoourvmUTm1Zidj
qZ8IlNfy+xQL1Ep5yzNUE8JVvJ6fFbTSBip7QaFapQ5tmQPDmdC/DUGaqJQdi5K+
C6Snc/1HB+mMnwK6g3K/HWtMbpFExoTK8MTlT9PHuQFTqeu8y8rv1Git11q+PGau
4Kj/ECNoixFqruSawxCmu+HWwcggKI0GG1uroDCBE21EBSnlNhzzndjW7utvKCc2
VHNppDB2jgv5qfwfQM4Doh4q0ACTxqEcM59tz1v1IT1OsnHzEg/DaJIfOhFpruTA
vgFoawJf65272bFWfN4APMw2INpYTLnf1C1RUGFW97Lex6RkYB1Ka9T9E+t4jplv
n0vf0ZRe52ml0RrcWorXUzDG/tO8WCEFUdd017T/EMR8OZqWoN0CQPhgnzhRSpJZ
wC782tDjw4rFdfNHL0vFESWjrwy0zuGYA+uqHydB1NZBXF1YzM2Rr1dzBTAz9Kce
luYmw7lL0Tpm6ytT1XzMgrSBUUk4U6vC4wjBk1VWYhXOomfrAyZNJFzFfyAYKm4H
PJDPnCcPabY9Ga0YMAu89MBo3frEqiHaSCPQYUGJHXaimTj+Yi0V/cvIHnQa4yFD
pzSqSJjmM9o0j67Z5sTzeJKuSptcHHt+dMujaU29T7OJpbYrRO2mpcvOfA+HahPF
15/dgIaV1/oHOMj5fqP6WGeCyj7Gc77p5AkR7Ztn2TvDCWxaGnQ1EoKZty/4Y00R
ObtGQnjtNpvRyTViixsZJEl76RDTwt6sa3buWk8z1e7h8eFYhB5w8Jn9Vr8A7EbN
IJXG1njdTJ6L6/oUPNVP8fZZOWcvqlvf5nQoc9+ne8ktUReAPdoPUr3YyqWeTOnb
fe39fOH93+TlafskZ3VvdwnfpGrCycA3oprZcKI4CZMoLzPBYV/pRqBWBks1ZicR
I+ynj+gnroSzpkAPgHI3UHG2P6OapwIbNGMlbTb2t93LoHrLmLEIEXYtg9Gw+SD6
AfBCi/+JLuDy8H2mtG4SlnItJYb43QMwijVYbST1KZ4ZPNe4sn6MrD+TCcb/950Q
BPmBcAy+1v32/YMho2IiFtIV/0YsG5TOP4NvVBhZlJzbyEdCcoUTyUJwtepYJ0vK
RRT9EG/6kc3BhlTp0pRsedFZqg8FaJcIkqTv14r6eEkOS81Y+frJKweF/XA7pwzU
DQAv8n9jjkIHuUMwge5xTp+7V/8yhQUGhYszPGWgXKuAQyaLy34hqvzT3jviRizM
01VLwVdKrvSpt6N9FI6eFa9fh435LRRALzOUxEEQXq9ILDNOXsgZxpHhTdtKrbQY
RbE+tKC2xlVqC7UJoQCQ1DuK6CdElvMSvH29Ug63xofZh5FrzzJG1kMNpSrqN0S8
1RtvWrHZ/6TZDszeOqY3ngTm1G3VdPFCP8NTJS4TR+4E2X4mAnS1YujiDbZNUHsY
arc2xp3svflz0V5iFw8nLsLHCgNMl1Gm4jEINr4cAZ2w7YlM3CyToyMNF2XQ9+Ld
sLy2BR/Igr0lMVNLm/9wQ8wr3d84MKSOzugn15Jx6MGqECYEmwUJ+Xa8VG/XoFqv
XBD/aV8wpdwHc5zKbClRO7PYbj8fod3YJn3TyW5WzQGqeUfrWdVWCagixf1pWCxV
XPdqS6ukGfslgO/Sa+quVsxl5JGNBrutlwKO7fOXcxPpgBKvVOXlsUH0DgBh7jIH
5HIW/bNd0ZoTUd17TnTB0bPbSnHGeNgpUg7t5jaW+SntREo95K3Zbdr0I4ArQVu0
pyFiy4Z1a2/wzM+T/4lgVbyYaAxaxG/DS5PyNSINkZkMendyZvwIcf9IdEqX1dAc
/qSH2+sNI/Xs4746avcr1Z2PYvUO92PXhh9l70xP8RKACluhM/If1dwD10qpHXRG
gcJPciMtK/j0tm/y1ICxLImU8nQLp0FKWU5/dx2xboMS6XE3KeedZqIwFbkW16qd
flkbhEibTfNCegJsQk0KJqNJMRLer4uL9SRabEL+ghojN8Vy6w3tZDj1VJQVrZGF
oj9i4fokzVLhU2zsqa//V7dQsJaBkDBvUOKV2y8KWuqTf9FotGqEEr5XY8gbpFHf
itg/a4eDYtbg/EFT10cI5gy4PB34jNuNfmTHcONueopfNgZCpg2BpoVwHiqWdb5e
KOujYG0aN/U9CvI4Nqb02lU3E2zCs4SR41sq86o2gxcq2o0oy/9I5mT67NnvaE+M
ajbAfkOHyry5mr/54vKkatigg/WuXwUPGvKf09Ks3YoCMf2AcX7nqEWthdtxChyP
+I/IkW/eUlI3dLmBuPTRZalKAcmLaWyNpmcHZFptf0ibSL/Hj2hH6M7wJ7NO6cQh
eGBt6TtAt8D6v13y8KiDAK6OWYycH8FDct7Uu0aMf7ODtf01Dj02lNl9wqv61wp0
xybpGqHi+dgrjhK6myOqWcIlmnVPzQ+XiUqkzZeVZo+tr9qkCrA8KDtd7f3wPvKW
w/bUwJEFiXdREoFVrD2amEt5EJyz5HOWOkrZuOkAmojVzn+sOs+BFmO4j0kqAocp
2X76OT7451XjknQlv32CXdgkZdFkXE0rpXBKMwBvi1xwUErQWpsd7n4VmpzaSGP6
4h14S0F16JX5q9Xa0Uhjn59RXp5jN1bLBS6flB65pp9v/YXYMlzU+DDKn4I7hWR1
Ub3mTdW4UoHpdgw39iCcNzPzQ6b3WtOLLFvmirruoagOX98baIDKvTk/hOhVSzRj
mwJvGAWEDZwynRkFC96spkPOXKQxS3sRzmd8qcNNr0jkXpqh6BJ+LleGAsAzdMrJ
A050MqZfHqZt6zA8kq6H92qClCLsC8rPL0JUgeFsojEIqCrZCMPC5WEPFUbQ0MpB
9ZDczZcSZpUM0WTRiFjfQfTb2uZodLDXGyapNrNXjSATw5oo/J2DtveTGohczj65
1AWU84mDhgS8Mc4ii8wraS1JVBhP5RwfgAnVQ4z+1eUW9Px4oUTAu9LDk8h4snFL
usEdWBleNc2/TVWXrEQXpjLY+nJgo0LuPcprCG/+BPU/GNQ6ffFtFEmfaIzetoE5
Av/NFG23h1l0P0elIAFb3iwLl6GpEF0s7dP2my8AilyxVNBgh71ICNYTD4hsqMfm
K5RUqkcwl0FT8+XVizOqVSUn/joqr5tHNd16eyfLs5gar/2LD+HAV5oZLI1kuTwe
EiO69aGeFKDERjtA4/xpfJti6wVp6hNH/FUR9Bi8xRcFj7FYqhfaYYCk7S35lXaU
Zi9ejKfahcKXUETcl6m+8mS9ZQgY/wj9jp1VCkMyqryTNM/alncvpIL96qMdxPo7
ChxeuTQWMmQHDiSQOAwGTc6WifuSzvW3tt7yDrVauJ6Ym2xmC7QR83mPggGvabFI
fnLmJH12So4u67g0cBmh/c9VfO5WJhu152S//KIXVBgcLYnd0rLmuPZy4AJecgi2
IjDGyNhaGCU3Amf60SoqDB3A8L4DFNcU0fpIwv7+RvEP/8Ur7yn7VKzcotTOte33
A9mU6YceMrHdlWtMaMbSJWEWOEz9cpw8gK8cCcERIOIQKBIjaXertZUN+6X9UDvj
99qtMEcsUS92un8Oag7CVcNnj3M6b0r1hiU0I1H8me/BsQtyA9jri3r1IVxZB1Jx
1dy8uJefW0w0GI4+rMEovrgRhSCCRziSPZIBQwSNhyhDdfcOG1x1eWS7bHMkuKlj
xnSl22X2ZPjAFKJIFTNAqGNop3NylgiYqna1N4EtGxeeHRza5my9d8lj0YsLv7Z2
ZB9T5u2RFlhqcoheNPl/i1FVPGS4hpsh79ZeqOhQZk1H+6q/JIx4Nk2q6KNqjdac
W9ZVWjMyS2/D0vxbWcnFWRSKdzbAkQPIndZCqKQdIA/nsxfw8bJjADjgPjAr4dX8
iGAmH6pfO+e3d2ghpC6SRleINYmqfC3mFpQqrZPIajIKdKwKQRGB+mKeuSvU7CN3
KSn0HEK1lVz0HGa9XjgYYHHig/tpDH0+7acHfizjkdAwqJYaopZnYbVocvOPDvP0
WpSC/hcye2jri1JNKTxRmtayDLIT2haJ9jvFDfNwZIDnz2n7he7n4g/aZcHi9YJT
wq/MYE+1zUzsgKVYlqpP0aZ1k+FAklYKMPbblcnG6TpSTcLhmENAyguVazDaw03M
vbmvQjeo9/cDvMn1IFiqRr3g14sLD8h1BfmNuOb7/tLRQyHo1zd7zqeBug8bygSf
f2+dPQR4kxUcgxtXaiX1dzQrUoIFgA9xRJ6nPInT7GG6zKWN+oGsxnYFsDdmfzU9
RYMUVDR4WXPiC+6aa2sj4hHh+j5n92hIhvFLyVjWXmB90507q1zgao9lHTMAljKc
rmdvCQIPJbbC+rIhMWF2ULp1I/Jjcp8uJMe4dtP024zAmNNbaRp/u1JBloqSOAen
1M7R86EAXiaCDSjxy9qXl3a+VMnssLAg8s1OwmyqN0ueIs3Ab3E36Wx/N7fqW4up
amuaQrjnFPP9UTfZxNuXL9AFxAtuj5azRsF/Qxa8rCkExUbU2ldgrzboN4Gj9/W4
0uL49lWSO4qv+dYrLJbzn/nfgfaL52IeovO3xSwFMoizD5dpWI/hDMfdV4BPHtLx
Yy7Eu7k3RJXH7RI5JYG1CcfS9sfN4U7Tvj545tXPEDVX2DI7MPDu4Udybjaf2NOz
ghphBL2uG8JTwTnIj2O681W0prbHjnbNqtv8oq4ydMX+S/S75OOA1ydfgOTC1k5D
cb7TCTEmeJsI2M/42cVneoWSDOmBCiOl/tCfrckBZJzI9nACViNT8z55TCtJ1F5g
t3JlEaO8fasC3d3COAJrLYMDeMN4TgNMjDOUQkAlEr8RVBiUo6flPFDfMF1rXs21
vZm2YB37XZcWkSaIEM5FmmXiLcjQUwjrEdLfRou5E9uC23ltjTq9T8e7zaQbsz+m
1iK+lj+QR5vBCHLis1tNfh+tE4rX5q/kpSPb3xWi6tXVSrPR/qvBC4ajBLSVOQA0
3yv1twaKTvZ2Ldg2W4yjxmFZNLV87HnktUslzrPG9Mla+qtDX0ppPEdPndKRjuTg
cBr7Pu2PjGg7K4oXhRxm7eV/bfKio7HuBp3vq6SPbLGWxvbUOGGXVEcRFZPFJV6o
rrR9eQa2uEUobfsLon2AYybwv+hbQOI8nJpnjfvNKDpBEvuYFtaDcd2agkzJ80KL
Zq6+3JnfLeu/SJWi6xsrp6XIe9j57+ltazl5HuCqIXLOCrs0cCINXmy4+WLY9Bhl
MNTp+RQekEfmk35yIqIZhenhQa+bBcUNfRpdbKR7AS2KU5L63V9JKWah1Onjg/9Q
7+m7atT5OU+aNL+VjlS+FJ3hWmVl1Axwsz20g/BzY+z4FA4fLtb9k5QtiXZ6uOc5
so+glMlHlomflKUFJ7BRDuDIt54oMHKBc69nKxrVS8PGhcy8WPRvpA69DWH3NmmP
sOwseCj/UGU6bnYJ2HPHI99ZFIhD8GE17R2KB2OU6GiZyOwBuTzYqs9YIqdXRFBM
Z4lIE/11D8hbpVzSV31WS4wBAqSqt5xAb3BTNH6MowWkEqnULxCIsIvjYVP8BtjQ
BeSUR8UeVpMGN+g9Op4FqvGykgQ1RJfzvDzX51O1JFowoswxFf4r7vNC3CWyuQYg
OY7dKByIXVytgyBhDO8tcsf+DQ066cRGfI7mpnGjCDJrQ+eN8O+FZUNZa4xwXunj
Ga+CP6/13nKfYR54eHL6fD8FOXykaj9pW0MtZ1ISapgyMlBnNF8oocbtWaor7Szh
9o3SencDgcsMdT3BtU1oVL5HQGX7RQY5beu/3DN2RrilVYZAJjAx9WFAfwCo261J
KL36TO45z7jOTeoQazLVH6fE9kG0kwfO0NDCDsLhbdHX+ZilHF0FLijd4mvvtmj4
l8YOYrdwoSGyfiDjPcTG6xGs3Imz88544TwagE4eGD3PiWkaVEc0FCZ2TJnP0s/X
y6y+eh/c4x7Qpwb4zP9aVGCd2hXLuqgOJ4+6SavFU1DmGSoOU4WpWvopKUuBBAQ9
D9+XdS/GTiE64jocgCmgyobnoOa6WuhT99qdKf6PUCyNRYv2ShhHssMWjb241biD
jeTI6cHNYOk//Z08WC4uC+luOxXds/AGEc+4kb5B2iIl8mqGl61H9BMa7KYPDUIJ
Knouc33luXHaJw2kqz9MMM/hTNd8RT9LuqCUhun2EY9y0tDIxJpiAf1+m1O0yPiF
ae8Jdh7CGzQ3bjHKRMjBjt1HsSqZF7PxPNbrCpu2dyIHvvfZQ34H06AWYcsYgmUS
Hl9nUYJRH4aGjSqJudK9uW7WUSK0H5rrEcQ1sEAefuJ0UHsrP3rkqwkjSgFuSviv
`pragma protect end_protected
