��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�/��|��ס���⾟B�9��S���r��"�]J�(albo�YG)�a�H���j�����1X����XDװ)	򒇍��_)���dK����~g����)���O�</�#>��r�}��n>��W,cM4q9^P�f��2��Y۟�aI?��+V�*#�uD��(����(�ϕ�Z����b��	5�%0���ð��[��k�<#ӓw�� x��4��,,��L�lb5��z�/̡�P8᳇Lٱ�ն�8J�:�8�iK���r5�*�y�YP�v�t�~�����V��QHG�W����lͰF�\g�z�7�Y�a�w'B�Lكm����c�&����Q�
�kZ#����n�jp��_�w���w��jT	�&� �$&��I-ԡ^�sY��Tn u;�<n�c�m�)��A �Rz	W]�Q<���)��hZߘ���C\�-�=o��Jᔵ� �/����ā�2�2#���Ȋ��a�~3�Ż�$�j;�}*1�/XH�w���؜tK�r)%�Y���Fj-��t��L��-���!���,��K5��yt����e!�M�a�$�Rw:�bG�� �t��}�����F ��XU�'��Yz˸��j�{��9�����S
���\���h�{�j�;�ӌS��wɲ^�~^M5>�zyΣ�g��8p�FA&D��}�4��d�O�Ci�
��
�ʺ�F??�2ů�s�aT��7XM�{
\d�3Djft��ׁO��I�rf��Q\�oa�([t�/dꙈ¢���g�����G��N$*TƭRM2y�q׎�pӆd�مнo:���`�cɯtٿ3a��yS����u����fN+���#��������B�\e�u�m(v���]凚S���at�#�ZZ��NAoiښ�#��5��eӘ��dH+���x��#�.~j��|�x"�י[]�gRU0Ĵ|㕱d:6�����Q���p�5�� 5C �[�@�\�	;�У����6��Anu�PyR��Je�ulTJ-���qm����ָB���[�I5��ߥ&�g5�}J#�v��4�b���k�e���
�.���y epä*R�z��������p�� |��o_�ĺ����U��@���tV��Ҳ��;���4Q��lc,E,p��D+�	n=����]��>���:�\�[u2ad��v����f���N�"a��`":-��^�)�|H�*e�������r}mS<1���hOm<\��6�v=�)q�BF�M�u}T�n�B�8�ݧ�.>!��uaC%��	�0(��D�i���-"��ħ|�`$usW�쿕�bF�B�֣Џ��� v9FB;W,��C�l�$�/�÷W	�U�T��#"�e�R�M�5��f�oN�7���VXlm
@0'�f+�_��ߵ���:�T�fFҔ��M�.$IQg7����M�)����m�8a�@G�D>��]��HF�'ohb��b����'y�(M�&��4>w�ەcP&L_�1�1i��M�;e� F޷�*n̛vL�5��~n��_�hz|K����
�WQ�p��2f�2�^TK���>Xc>U�Vi�t�:j��$0+N(�l����d �Y���6Gr�p��v;}*��rT�4��!ùb�a���T�:1�
m�����2� iE�S���l�4n�_�C�q��hk9�n��3�d%��`J�y�v���.s��~se^+�">��(��#�3��31�M�H?�b|w���R�-X	i?�^�Wo���)�W�]��m��'o.#��ng�-G]B�}?�h0� b~���e n�U�0p��Z�1����"Z�ҕ?���N7{E���ow�Ay�Ȋ�K�13�8�x+^���QrZ�������~ppLmz��j��y>��Xk�P��D��jI:V����L ���-��e�r$X��7~������'p9g�<k˴���-�� ���)P�r�"D�>T[/!���j������0'{>r5֟fâ}G���B���mz��D��M����)��(�	>�8't�Qc���ȝޑ|@ ,4��J�w��Y�s�2�����<��G�p!�c��O��⠼qݯ���e�Y���+4�m�o�t2�9��>�lp���a�����*�aV���27���{/���ߨ��i�@0,?�tzB�����8��p-ᯏ���.�� ���8����S(#"����\��++r7"E'�M�N=Ԇ�S YNnI�J�h����S'����1Z��.����&���1aX���"�p6L�%X���??�2Lӳ�3��8DC�bO�}�u��[��ٽ�a�/����'�� <q*54w[ve�O�� u�/�O?X���V�]�#U���R=zy��m62��=�!���T: ���L�(���U�m���ڙ�J��s��HTy�&p��*%�'�I�#��9� ��QN+��w�� )��B���2��a��_~�̢������!�7�"��
<��*`����(OO��*�_�~ -5k��?K!����W�FJM��,T�^2{��m�8��e��'i��ݕ[k}�C��A
��~�~u�~�_��j�����h�,1B.�yfl�!��J��h�Q@���]����22G���K�p�ن�����e\�p2��)�"�$et�z��������-�֫Za�
-$�dcŦ)fn��	%�s���zI��rur,��FXƻ�2)�}H!''	+f�=�aq#��������X���̯���"�	1��?n;Fݟ�R�an(wh����"��ϛ&	N���0��,�"l,�Y�aV���Уz��ۂ��cX��+���V�̰2`�x�J\�3� �-�� �wW���i��a�<�3Z�b���������{��~�l��j��mƣ�%��-`�FutU�����P���hPX��,�@F��3�|#`?��ٓ$	�(�*�"�g�{ R?�Z2�m1�و+�+�Hp^�2�+��|���"��G
k��K�n�q��<���pY���#��ٺ�q��LC]B�N���ćo�t��V�a�P4�?��􃂈۵�\�״l�.JM��h:�PX\�⥛�⍟B���"�W���ήmZ]CaqV�U��O����e�*�Y���8��=K���C�ް�.ƴ�����7�=Z��A��ãֶ��΄'R���E���U���.s�-6D�rI9LCp͏�T�h\�i6�Qh!�z��r踥�Y��8O�9���ڍ�]s���X:�!�
�޳�U���X^��� �%�*�#�-�,�5�U&���� v�{-*�Г�>LY]F�Q���A)�Sdmg} ����B�[�h� 	MB��XE����a~�<&����^�X��2�d�`���4l�l���T����s���^�̜����
zN�����O(ΑCw�KH
e��l�%�؂3�5<�Y�˒�:�Z$lJ��$>������]*��}'6\wA�@�8�H���gA�.�v�w�V����ӿή�*���4�Rt�ئ'�z��v���y=ܱ��{��FR�5r�^�� ��F�� �6�:� �c��=�P�[�����]�U��/���>���
�A�Ѵu���@:c�Q����6��'�&N����a��;���K����ʃ�qt�P�;G���eK�2����VI2�F&Yj���rȐe�|kG����u(����˦�~�\�)$�1:L9��1%@$.����j�v�u���@��_jG�C�g�;�o�k���E�˽KAI"����8��N���S'�B`�Mv��Vҭ>�͊U���vb��Era���o?V7��(�D�q���c�|����u9D���0V���9�����g�hj��kR4_(Is�֕�2�����/Q����~8�¶��O����}l%*5^�TA���{��V�qQ_�g�Э�
��x(�1���a�H���,�;�3�0\3�Xni�g1]Ԗg�~ ��˃`��-��H�)��|��䚨Jޙ�>O�+#���V�@�z�Bܳp�}(I�#���Lɤn������V��1�Xw�V���q:��ڈl�d�#+�*�NCe�e�o��T'���B�_c�F|�T ����*�@?Au@��턅�0V�ZR���ק@T��%J2��"(�,���j�d�AXXoae1�e]-&�'m������e�g-C#�H����JkB$�+�5e�����5O�(T�F	�� �t7�*d�G��)��8���W��ESA�F�g��g!�6�:��KݴR�5���?����+��2D�9�^�b���M�
QPlB���"��c�����2Oe���2>?���7/'a��7�����_Z2K�!g���'���<]X~���l�e�wQIT�F�8�M*G�uhn��o�Ǿ��E�]�C��I�\��;�YO�W|�����K�7V�r,����j�W�h[�*"�N��4���	>j9��]� �\�[�c ��g��R�����7��Ce�k���{���1��8"�2�۶1��Q�Rr���~v<kp��H0z3 'w� &�8sEle�n�א@���Af���
72ĵ]�G�A�>����,��c�������#��fax�	*�B�͂U�;�F��My��E�h*.��d;�l��Cx�/�:���6�����������j����Zi^ ~�f�m1N��D�똆�;���ā���FI�y^!J0�����鬻��Ȥ�Iж�6��tL��O2�V���V�f�F��_��%��!��6]����N�e���ݮ���5�n��W�R껏�����,v�>$��{�!V�>��m���뒫�7��.�/8�	`*�:��b�;�������#+7��|�~9-W�_��`ĔB �/,Ǻ@hx�H��g�ݯ^>�5զHX��PT4�<P�a(��@{�'���,k(��!ʕ���4�4Zu$0�F��(q�V���h�x�aH���`�e ��'����D�ڴ�Z=Ѓ�@�Y8kK|c0��p��
̆NB�G5;�QdV�`�D�%v7͗�s2˘���W��<�rT�h�L��N���I��$�.�rV���~�"/�Kz��`������-��D�0Z&g.������GR��-�41��<�a!��e�8"�?�.�m�.�����ڞ1�l�9=Z9�:�%�x�/S8&1!uN�I�l�Xx��*�J9i��PR��ނQ���Pi$��G����.Hd��������t�[���������M��*�g��,Ej�ג�&��Ī�##S�d~F�c�o=�V?*4�=�P{̍*������� ��w�1a����n�-�bY��yi�mIùƦ�ܶE#�b����'��" W���U:[�܂����<Ԯ?|O�iC&�����D�t������~��b	;�ۈ��[Ku~�
��5��
��?��2�e�,����P���f7�i��_��'�Z�?�wL����
��Y2�*sp������ �hLJ�V��nY?�YP�� � �\~��5m	���j��~D�e��Nce�Y��ˡ�����m��.!O�AޛNHg�QwL`�1��&D��N�N���,��Y����&�?҇�P$�e��P���׽L,��r8�B4e�a�W����5
kb�-�W���g�Rw܆BI��^�eJp�l�Ӄ ��vLD�7S83�������]�a�%�<Q:� ��U5�E8��$�5ƞ�Brn��O��sD�?�'�W c�xD�����'5�+9��,���\v�Lނc���f�B���d#r�����؟Ը8@C��FJ}����j�<R3�n�'@1��݂����8��E;�j�B�H7�MS�B�!nf��z.gB����PH� E^)?k{���%�A4 �������	e1z��p�N��Z&�)���d���_i1���Q�cF�-��GHR]/�i�Bע���f��v'�UP���д_�����|�Kp�ҍ�������<V,.�2
�gA�xN����-僨��� �8���VY�!�(�Ƀ�0K�'��{����|ٍ�9���-@y߁�9$_�]�Kx9���T�U��jG�
7U�{� frᨵ ���H@���N��yS"�^�!���ٿ��	2�QOe2|�_X�DDx��gnO�LU��t'L�����k��y�^��m�^c��!��-!Q�RMN�CM	�/�vcs!G������خ���nZ��S%wL׼����d��L���C��{3p��cM��͓�Q�*�	TBQG$�X@	EF��-�Y��{!!�7�|�U���?�|jg0S)[K13&c��IIї�N��ź�Y/���B�_��*S3mX+\�b(��3�Z���Ng��CAl=�F��	؀P�w�����˄1���IJ|�D`mh�u�7X@`���}�t�`Zg3��E�ϕ��ݩ�8�X«|�]��m4�n6ڥ�^�FC�1��R7̍F�O�^�{������=Iy$2Qlu��F��k�g�l��\FHӉ�:):�PƁ�[mr��q�Ӽp���W'e��o����W�Q�DRp�q*p�Q;��䴭�K�������b���Z��^�(��bx5�,1�d����FM3�3*�o��t�����nnj{ى	�r�M�	���r��4�������T_E�O�mș��<`���	��M��e� �L�ث�:R��ZT,�\�(`���4}��e�JU������DR�{"3[�8c���wz��^�G�qz}eɂH�������|2@ZӃjڍ���1�]�����9��gd�O��)�J��?� � |"����]�*n�CT�&���3ǨxN���u$���xp�ni����<�7���1�K%��Xכ2�~Zlb�ɰQ}"��f'S4���wJ+̀߫��g��)Ɗ^�+}*�
�B_��xBʽ?Z�Foj��>�F�<�ؗj=����^�9�V�Ңw�/�C���1�xK~�L��vy�#oE[��8�*�eɩd\�wl�A�����`
GUB�OLkަ��{0V�$��֔��(xԇ	�U�A<�as_���U�,�����	�Z�!^������Ũ�O���n3vҗ�e�Mڼ-���9�TPD���zTy���}!�&Ϲ�"�*;��~7Eｔ�N��WBZ� A��_D��ު���TQ�R�g*��A�ڭ
��5�@�K����P�ej��k��C�Q��bA�,=��QL�kP	�������' �y�=��&ǣqJ1#m^O�\0�4�\��s�)ͨ�G]���g+����f'X�I,ً,Gk,��~��b�JphIf�%�H 
����Қ���#U����1�P�mbQ�G����/��Z'�i	�2�g����f7�Ω�sb�Hd�Q.,��;��$�����,��k�<�kίr-/+;�,ҝP�Tb����sY[M�y�sYܤE	����"��>7���9ހ����e���3�}���n�$��Aj��DcJ_煻��W�C_A�Ž�a�ҸP�N���H~@&��j�<�;]#����Vr�D���v�6&��K��4�?OF�&��F��xL놲&��M�l@DjY�)�EH;ؙ�n�cνp�T��}��\tN�O�p���[����8�M��EI�U6xrʸ4L9��ʐ?��c��i�'���	��#�Vy�Å�w���}Ao/�O��ԯ�Z�6a革�3� ;@�)�em���+w�������t�G6x4ẏ����X�af�$x'�p<puu��T�4t2�GWF�~��[��A��< V5���L�j��k4O�'�F���d�bMB'�֋�0Q���&;�D4&Xz��H���BXVLb�xl��M艺r��������C��4�``� ��K�!�p�|�J��G�c�G��z�����uG�!�n�eH-��Ym-zf���e�[���u����B�:�g��*9�<��������s�x��4h�yy�Rm����n��]!D��5�y(��W��в��`�.Ls�,cT���6�\������1"�B��
�݄03R��Qw8��d�/�e��#%(-��Zh���Y�]��Dnj��iU��7&��1���XFi�~����K���/�/�}x��PH)cY?��żF�*qu���^�M&�)z����VZ��v���_�;Y�¶N��pp��u�9��ԶIЇ*|��K�hS�M����`���{�6��	%� �!�]��	d���Һ�h��8#�3�������Q�g����ܟ���;�c�dܙ�&�5H�L �fp�` ��9ժ�/�f���̌�.�aY����ZƜ�d]P;j����<<��y+s#z��i��Jr_Z��R�ɵ�Ŏ���0����`�q�,���lٰ*�����9˰��K'���a��p%�?6}��v~꼴Rw�������_��V�P�/�C\���Xj�Zj�UP��#.*�>��"�#����E�~ib��L5��yʗ�y=	�J�ymȇ
A�����T��H
P���;�q�ѡ�h����$�hY�]�)��+�"����e䕻joPSu�+��;WsyQxg�*i�<�kS6|��8~e%�]ԀA�����aa,<�2� ��oV0�Ð\�j	A��ġ_��L�H��\R0��$� C3/���b<T�����C�S{��>s]�1��ї�\�H���٪���xS ��i���~דs���9qBí�ƕs_ˊ#D�;����`TЏ���rM��h�m)��$�(n9�_�ª��bB��J7p� ^G�ٺW�>ntf���2���Z�) ��y�Y����G[¼�r��Z("���Pw�Q���i���0r"%pi��e�e��yk�BTF��F�����8Ue���Z��˖� �11�R�����. �V�$"aZ;45/j�҆���>U���.�"1?U��!�1�
d�)B2&��f��J�`��:��={G����	������$\���1f�K�����O��r�q����A�� �=|WX���H,?K`�&��0ۉ�]�YxRL]y+�BeM&KM/o@�#��z�BK:������gAz�n_�՞�L��}\>�y�y����l��HIx�M8�$f�T�1=bZg���H����;���ǲ1�g�|�v�:N�;F���T8c�����7��sm��:�tpb@�^(��t��+!x^��-�G��4�/��\�>�[D��l[1��%O^�t���H���g"��xo�e�q����Ľ�h��/*�jTjS�"�'PEd	����uON���7��=����+V]l(j�!��f��S�Ǩ����Nͽ[ע��"�~�w�O��.��r���P��D+������H20[+MR9҅A�D�a�����p�kM@�_� Z_3�R�E|�Dd���`!�.��^���C�]��#8R�s&pX|� �D���7��9_n�QX�M�_���3fy��֗_���ׄA7�-"�ĵ�������XP���I�O�qг��.��XC�	���;�4�`�1�X�Dp3�x�"6]����3⵸�$�15�'�? ����s��ڞm�Q[�r�D��4 ���,[ň?��<���O�m���.��
�� Ec���=s���3͑QW�p��_8�Z{�Q�nf��cq���ӒCj �2��ƚ"���9J5k$�l�P�ߌg����l��D�M�Hl��"��wGL�JM�*�P͋�"��+��=h�F�:	{���m�'�g�\�y֪�T����q?��b�9���"�>l���#UbKY�`FS~��v�f�8_ŋy1!R��#$��,�L�h1λ�����o>��	=��q34�'+����`��צԂu��EKJ��La�@1�����3�~F#�3�_*�a��{#Ю)��7�m�Zp����B������<�UۿTUN�c��kn���-"�oj�EC�[^�;��D���p`��3�^�gr�_ւR����'���"FN4��H�$[��R/��J�L">���,��|����B@��F�3+ ���*~����W	�.��+}=v���	w#���!])��i0]��Q]�Q&��O�ϡ�Kc5�5{�p
c�a���kd�l�a0�FW�����q����55�UB��h�	&`�io����M��,׉𲌥��P��̞��6��j20��� |_��O���Pa9��+/�).`�&7��_9ƚsb�d�L$�x�%�3Y�f���l��nU�T˯l���xJ�[�J�>�R�x�G5.�J��$�A@+�.���p�S@~���w����F+.n��B>�l��
A�}��(;��/�zە l#���������uy,E�+�^�h����j���1��NƢNϡ%��U�r��</��I+P�_�����������*�`��gk9�:䖜��su���������H��y��&.v�GM�U�i��<P�jR�]>I�թ闐ę�ɒ����0�u6�!� �cj*j1A��������s�C�0�+)�4�5e`6U{ГA�BS2+���cyf���3�ui�_q<5�"�-���P��k\#c�s�J�	�h� �O�/��pzabf���!$���57�y^����s�=��%��}y![�� j�f�jp���gYo,�Yt ���Xd���-��+��c���`�}f�Hb�����{���7��O��Nǋk�#�JQ�ύ�&E#��{.ha˰5Y��ŌW��qy�ub4y���'1�r�.ҧ3qT_�碄XBMh�M(�#iϘ q�6i	�x�m�zyn� C�l,���(\B��,�t�����,%yZd� lg��0�d_|�t����*�;�1.�x�o|���B79����"��	�WRd�t��j���c��t6hQ��e��6�?+Y���U" +����R��c/=�n?���MT�ʲ2�D�e�Ux["�>5}n�� �1Z�`���+	�5#���N.Ds᥶STީu���L������ZK1�����0*�\eݭ./=8 p8Ɂ9��,�_Wm܃�Kb�_�Q���?W^B�[ԱB����$2kay�e��1���'���#�r�JV`�"�-��-9f���IZ���c6�⠸�R!�[tw)5\U�>�L[��2�q"%�qhgD���c'#,0����.f���SliWn�)�>��	-ap�Ŵ�Fm�X�,,B�x�MH&��p�y�V	���%�[�`�t\��S����k�xD���L�`{p�*k�k�5��8U�q��zU���?�Xs�?jY��C�-���c�*��kˀ�, �������r���Ao��\T��������}���������n�K����aI���FFFm|o��,��ˊ��ݳAK�����P�1��+�~�P03�ZrD��4�R��ΞBk�`/k�����y�-X�i�t%�b�����LO�=��:�A�<�b?�.]1�kN/y����a�2�ءuC��2&��'Ju�#1A�$jmx�|��L��q\^"\ER����o�}� 5���yp�1zn4�.2�I�(;�fm�G�ԃԺ�0�Ӟ3tn�����s�ѭS��]���Uk(9r��� �J��驘�E�R�2���6�e�o^����{v�^�	��^��8�g5xV����]��9B���)8@ 8�K�S)PdWQ��r굵��) �.�_"?X��ܢ�.5�JY-��4��+F�*�%UH+�3��Ć�[�"hQ����+�Q���%��q�\mr��:��S��޸��ș �F��v W�'����O,Ĝ�E�3\z�����aq_�S;w�Qg�Rd*V椥���f,�Ѻ���v��[b�pFn����B�T@�>0~G�&,TL�n�%@C�D�I���y��\�.�'7į��5�����H����s�-^[�Φ��d�u �'e� ��(I��[ޥCCk���%�'j�0��m;��N�ܿQ`�ι�%��O�B���1�vl��C�on���35��<�b:�P�ů��lJ��~9HB>t�E��t�C�=�E��cBJ��Oaq�m���7mҫ�!@��c�8�Xق4ằ���t���L��`��dYN��%�l�ͮ���a_��n�h�������c&Y��轤�ɇ>���M�ؾ���n�J�����V�GK6u��)C%}ܔZx�P�f�����aXz�����+ w�b�))�NSS�3�̐��'�	�K��1.0����yY�g!�
��͟�`z�����-^��u]+�"���D6c͝K��Z6�v�;���8�y� �_Xq�r�@�1U��1R���|	5�K*&�!�&�?���(�v�a=�L���� m���ؿ�u~Wej۵��1���q� !=�^8�h��/>yNH�]C�1��T4�c��7ꋵ�{��r�<��� ��e��s��I�4s�h�Ǖ~�_م������B�tH��4eq����͖f�Ol,��ͷT������8墠�	H8�mg��W�"%�G�55HT7�dԓ�QP�7�͆�C�l��v����^E�nP���"�}�����<}�_z7�YP�M}�����8ݸ��ߖ4U_h|y���n�]C�R5d��OY�����X6��+�.�@�usU~S���q|�}}:QY�n#�:AWtqၻ��땀t�n�Z��ȉ��;��W\��l����W@�,F�n#���J����m`Ř���y�z����Q~�xD^�K;x�\�7L�[Z<�!�k�	��D�xEw$'1l@��X�����n%cd�����&�igc�\�jzY�4�U����˓?K�3�� o��x���=�JCZe��VnDf�l|*��گ�3�2��~�a��9��r��<x�jg,3�f��0`P�m��M��k�Ih���n�fN�2�F���N���yf+��`hL�����pZjc�#�0���T�>Q�,U�~�&o�LU�\�9gX�
4dF���D_���a .�vF	�kx���	��m9m�ߺm�-3	C�� ^�����q&��:�rl�Bk�G�yB�p��y��Ye���p�yg��#ߪk�5]�El���߈���a̳ڡ>�L�`Wo�Š�h&�N�}�z`����Tn�<)�(zU�����R�Z�??J����黑���2�H��!�晴pL7O��7+�)����R������v"�_�܉�g�j�1u+y 1u�x��,����v!�6���9:���'�4ss���Ͳm����{U�c3Ɣ���Z~
�����ue�"�
�h7�Ո�ƺh)|H��%�����5R��'s���1M;y7��T7x֧��&��	�>zTQ2g�g��5��e�#�hl��Y��B�\^���.^^��LO˞C��������z��+��]�h=��r�����0"�CNۀ����,���.[�>��mX2�v���C��F��ꯏ�	�,s�e���f���t�7NI8;)d3OY]�<��ܝ��wך,���y�춶v1Fj掷/@�Ę���.�$F���z����N�\|�Q�����U�+���#H���RRn�+��⁵v%��k��Js�R?Ӓ'I�Ӌ�.��B�g��-�V�&��g�&�?��p�p�k�4�X\�(GT��9k}�{���l>↶��2���Xˍ"�����:�&$	�#�]`��<,c�}��)o����e������L�Z֘����Xc�Z_�9Ì����.���K�%Vzp.@;<s�a��>yl�~!;QCk9�}�E��d���t�
\F������]��#����Vz�A�pB��-Y6 ��+�J�Y��Dw����r���0��z~^�JȂ�͈U���㴩�8���ybe�q���m��<":��h�,_P%�"C���������θ�v��������u>��di>aKц�R�bMZ9��e�)�HZS���=�f�� <�q�G��$�S���j6dcX]��&����pr2��`�?/c�����������G���Z9x�4�pп!
Htl�@Q�g���+��cx�<�P��_���i>�!�ł?٫^&���'�G.+��