// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
S4j5VwdY+eEB5J873MFSRGACMGPEFTXecWz/4MR4o1i6tRoklNZVk4Cq7MQFNI5+SL70Q2sNbAgx
SrIhVCatlPvcUp5/kpYRvfgswiGrd8KjAl4IALkLX3UWTZ+eqG9ddmZbfrW3iSwrHseTfauD9yUu
HWGulV0sv+zLv8Ky09rNZPMy7icOzwWXwMsrc2w/HOLajH6/xlnbujh94/m0EWMbXMpB6tm3kP7J
ZjtNB2c5BQi3aXO8kVxE4NPbWpF2Dt6o66H4hoqjo5AJ/dOZPrkP7/h6K8h/kL9+wrCZTAm9BZTL
5KBEgGGfdlTCK+k8/jFKmYojVYsocC/zPnZGmA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9856)
y8FFCblif9mIyZzGg9sRmHheSgLJjIwP16oxHt2Zo1NroB/Q4j0x/9WiMh+uN7WvwLu541XyNmAK
G/GKvnwDb29AzcuIehRfozG61Ghh1O15V8OO1QDICLCYPLXPcuMvkTUrR+l3k0XF+sTANQ/r4GXh
GBZc+hdYwBYptX4dF4QWrjiwkP0mGLhDp/bOt8Cs06hwkUFIobfDr/aiMG9N8zrxhqHdE/UJFZH/
ymx3chps10SHIeZ+inrbefpbnQUCVHNB7/SVieh+wAvRKvzioUN5qHWSd04Vxi9Asx1WDBZxBGSB
Q35LfM9kFGrUzs6D+dujMJP5MAQehFfQR6Xz1zgGgOroxocZGrC88cI+gf812RqKJRojgujrWaym
EobTOLpyce3mezSMDArY8v8sMedONSxHEB1B9zx075rBychJrzOAnkiQwsWPsjwIN0CAilAcqOVB
GLv9tDGTfXxyKd1X5zHP4sWPGFp+xOkv8zU4fklRGWKOwtcWcSY+17kE0d5b8gpJy+9FXma0UZuZ
WAC3p3WORQYNfXX5ry228QalC3JDxulGeqej6i2lgeIuUgHyKTgr18V+xrjEY/HvdogN5PXMDWd9
QfqustL9MXEtJsNwmqW85ho1V0pWTXVlBGYPMpLducZnFXVnSR/IjycvBzHULitMEvKHYEKt3ccz
iWA+M1bVJEOFGWCdOb8LN92vr1VjC4qWFLBqu81qL1KoBXibRoHSenbWlnzH8VMWkPwRaWLspzlW
POPQE1P4hVUR5jqZWWI6EKa7MxzN1BaijI5M9vw2sUz8VVu65xA3BNyJPp4SZ5MYMOJ2fos7dwPf
1RWwKLnGFATQWLOY5CrcS1jXv/m5B3T2IGvb5TZORWx+pP27dXY9+GwPebLkXaPNQqIEXQEnmfRM
vVTA702w9W544DMpOgt+St243sVuYYZ/vGmGQoYuGCMjrvj5g1LMyPmJHYnTD9eHlT1pMKNrHoyI
lwJpBVnW/SMU5hIPC3/VSn8yh1ATOrdEWr4jEv1bjBJ+P57vDrhwDcWTXcIcMceRtCSUbub5QuJd
hR7d43VNDyzUZcQSUOH1FBOCT1I+nvXQ1Ua2s//KMQ++UvWtN/YJMMIgcj+H08LuN6yHvcBMXOeI
GK0hxBeGRcVAKERdRSX9+zPvp/JB9egw0kQJ8K2kdUMf93n7MYAuMVf9l5IA7+QkH4cXwk/IUITD
gjF9g/Ae6LFjxLmBlJex0Mg/RgvfQFkhwcyfmz7eEfZMnACtrmQjm2R0OJcLizf97m/O+EhL0hzi
R31QSCOK5Q87ux9UnUUD/wPSEvgbBpDp8b9P7ev6mRnC+7SUZ5mKEReVeK/5xgUyb1bHISOGIhVn
Xgi0jNKDPqXBmhuTWJw/Fdt0faF1nqTVw34l77Pq91v7YkcoxFLDihez9Lp7A3cHlj3HP4u+FmN1
Rs/1VVPON0OdlQwP03wJl4MccWOdBaFLdd1haLGjzfiqJTfTuDKIpU9CsA3Q+4Ib/aO9mjBvLLQA
6Q3lQkCmM8krJJjkVkpnclw756dYXNoaFBpfsX6AOzpxSu0aaQ9PKnboS0sXd9bsD3SJdFBRvtvU
FzQhSK3ApYltj06hpJwrpz9nXYveFWUext0rudoaS5fOZghe09+onLTrszX3CY4GssiHR9JgSx/b
tklGLiLdq4wCQF4lIIuNYAmQY7AxbsbujVmeb/ICtkV3mMuITMX6xRGpm9UcQ37XJTZjh6C6xTCz
XaKVGwfhOFV5o7EkoeF9VgF1vFRoYITo12fNb8Q8j9+FV92Sc/P8C5oRXyL0E8cdZKTe2xxVZqva
qL9DyegjhAnFKZQCjFd6skYj0x+vBmScU+MdPLQxRmbkNphIB7IyHS38k+pdKcNRUVk/okNuilE2
EKoRgkaGKmh6knLjRRM78rSyDBkFHyMm5Tpt1t9SmAsAQ/Zhdrf9cJW7FtcmAKUG5Tb64cNHQb6Z
QdrHwAsD67nbw8Yie0pGlfnmDnHAGAN0oZn9JsaTsz7TXS3LB7B442mOeuJbvVi57dBI6iXN57KM
xtIVGuBQI4sERLATEofIURIACiq4BwnJLpwIHPfupCrjvORcsOW5FOo7KT7rjiicHlOXcxv2JHrN
ugGT/p26L9h3vnpsymDUBtmzOzdrJnei/8GZ2hprNwRBiI2E1j3njVB11yNpLrgA6HW++PehBq1C
3JFYBwMQwbihawPhIqXME9zGDXLfOwnBFEeFGBaeKpAMtCWX9PeJ+EA2814by5srYtQWOXu6KCNx
/v+Y5uZdimGX9DInft0FSgt0wh0x/kQWfuDClPS3RHy9WTvDcF5r587Eqz5+Ti2lt+moEhiEW4mJ
0p8MUZZiRUkeIRwAFL0rJnPv57tVChnkJtjjeElu9h8hg42jEf7kOIhfDSTSgupMKRbKmZpPK0Bg
AiorwTv9nlL2AzkbSEIx4i0h9qC7sQA46Cin8xR0EZaXzd6BkNryEgZ34GVTF1hEwEglk4Aw04WR
BJZBnAvv5+iWHSyq0pUsTCzioqYKNjLJ/c8OrAwVsdjDySHoxjBh45OnocCESvI/y3bOLtwOr+rs
B9WF5Hm1qpF0kkAEPJ8g/b+tpoyk9hxG4ke6hFOHLYkC+YTPrv4wA6hpe3ieNEGuJetLaZotCDJq
TwKiYSBrswM6n2RYpDegu7eXl7ZfVVoeHNm48YiBKnAVxBO1IwzWrUt/Q8h16hTxFDzsqgzDn/b4
Z3QnZrjGtE9u+6WfdAIq/Raz9UW/QNRzR9re0VEHzd70zACCADqQE3z20VgWetlup0KwGMShytt3
DXe/3aNAa1sDFPg29V5CFPaS9L6y/uD0k6VbOhTbFkE3PWa8w8NIg9PMrupASf97F4pwYb+HCZ0S
6vg+XPzET562NS39IMLVJxk3T9dHdwDAknimw6J61j5bvdbwYG+Gd3By6iGCqBnhwoEKTNCD2l6r
AWcMpm2pWzwAFhA12gcAk55B7SbyuTrnNropZXbo6XZmxCT2GpO8LlURoHTdx0rsJqjzObwJrtvT
+FF/RueR/3YNU/DYdbafw7kxa26SK8mq9hOZv+VIboawGYbqtUY40rJrJ4fHDE6PLE4ADy50zwOJ
D4Jk8dqAkyPtiV0wQ0/2qU5qA96BxvnI59MCxYN24essqCL+IcpRoP0hRhMlvZy4qIZhRL/IWKzo
AHZNVXxV+F25A8cvT1gU0rJqGTs4DYNDCzyRSqW9YX6KXSbTfMnGCszS9Alf1//dbG37fGaGkiN8
7G5KYwr+RTrWViFC2uUOI/2NOnBtxugnWWWsqLQ5WOQTpiwrFgf3/yzGqi5D7ZiWpnj26I8b1DRb
N/P3Ocym1puUNRDHn0Zr/d/y+FEHmS62WDvpuGeVmXnHbUfp9ppF/gXIO15EnADPGmh/K04yXR06
JGzhJghHnUqR/BiQ1ZHh4KwmIx/oBRa8luqlLU6jCzfAf51NJ5z/xw1AuL53QxAwfUOZaMI8gP1c
fIpT7lza0No2o1VphJyUBSSoO2iv/4RpnUu5dLg4oB1W12gXN6zwbOLiXTvCu9d7q3RlvKhKXs0V
RSO7xIZu+kDnu4Yk6w3S1I/CbcxMrwg0e757BtC3zZmnjW3A+hIjUkhNMs5JaXJ08U+9hdXWs5xP
UGNOBY4Rcz2HIz0VD+Hy8HVluTz6lCt8vlFygs9pN6eK3aP/js9lmbt9XmmoxcXZZNsdU3Yrfi3N
JBjyt4dt6ioOjXWWO0DEk48TEEcJomyDLf92Be0mAz/I/pti8KjEHfrB8HFQU8/tLvHC832zUqNG
yMrQpH/rzQRRLZzRWxpPX1iXlK7AKL1Z12PeN8RtP+Zc5lFamMKR3rLGQMhTr9vocCqkqePwvNJI
HF6xLUxaQTvQFmWkyNhEdqtssx4XD7z0g/uaB4RX/bIj4zFQsK8NUlEvts0zB4Bha4IQX/5U+7iK
6BLRwcydHPBORwfQv+hxnpqZSUEaemEgfPxAI2v1GpHbVbm9gIPro1ls+L5RQV+0EbUEJcKcW/aQ
kRsAgtlK/uwPvbVTTGAShz9epYhBI+CQerpXtn/PixDKNF7Z9+EU7Q3IpPyHBe/P/+DchurVOTXb
J43Vnox2P6/RuuLa6SLArIPESt2Fq7ARJ7oper2K/91T6mEeckNpma8C8wPel6vRY4SjLMUtzYGI
DbwkJPtiBxCApG4vnw7A/WkI0Kb6fQslzFbyvjJe2NHiZ6gECNGQXfhbPIMtqtzkiPU3WggeYlNI
S6G/IuEokN3TIbUvSTjcSCXplWOgIAHHS7SUDspDlLdcUN/tm/Gj8lOjYbK9A6V1GJrnFBltY63E
dE9kvInjZi4m0G8zFlP+6qtDZ2fihoe9ilA693EVMPdq0rE4fZ9pFlrI1VbmX8H6o+B8yPA+gFj0
eYXE5qbL9FdMF3cNOe3kHwfdBJ9DBA+62auWGtP0kcZIvR1PyuB6u3tm8hjGBiiGG8vYgsBGfB+H
QFf6npv+FdH/ZaKakiVFvzwiBHzwSs6r4feq5pswRnL/bc2tBZ3fEIJDC7+k2GGPWpuqVlD1/A/i
DjMnIZDJwenn/n8iLdJ5RiV022q/ufFRA59C1tYf0Y5IigLZsN+vrQwm/OGE0RtHV/AWqHh5h88I
vzahHJVtmupttLSCaoWPBbJEjVxt1WqUBMn+j0pOhUM2yO97ROv5o5xW1oWLeIr2BfKx+1mVPEWO
1VDWlanCByGPVBcGuKS3ubPrQFyhO6bJrqVclL4OyMiUEdDPkShnZFOhtNWduW/S/tl81hAqpI+x
/gyE8/JCKi0OTDVS156ZJBf2SYYkiWTUgdNKYHRjuxJn8DMtZKMfyFfHsH1EZf6oFbVG8+L5KCWY
NlUc6rDEIbskfiOkfKuE0XwJ+yX1QgVWC8qltGj+TPT292r5ijXec3qK2188Kr73K/Tsnf5zYyDJ
zm04eSojsUzcqTcsbjrHWSVyCJ1uYP1VLpfHKDj0C7DDs9zZ7/Jj6YpX4WNJpKo18D4Os3MT4EJS
jy1JUTmGm+wHgBL09ca+h7im63VJOU/xoS9IqXq5UcL4QvyK8D3MwoOJXTHgivygbvhmNzXqxMp3
SLRdsKuZMb8XVHGfpJ308SKZYNnnCCB4y6S3dQurt49xOxZwfBkvhpVkmHjnHcXYPfWNpxXQSYku
c+uRb3ne8Xg8qMxXLuyUWXTSZCI9Ovgppd/KfobnUPHf52pgI4yAtwnJ0QtuElrY28i9UXBXVqKG
CJorhakSyhgW1hW5k/NYVDZkXaNVYWf4IOsUd/cySPmC/NufvfkKj1PV2nxvMAG9iIQU9YnGZ19s
mLeH5eTP0rbikr+XbAH18q3t66z/yQp87r/dFj/HsaKPfTSnpWSanYmlKtcnOXEXCtiVKrO7fFQT
Vbgrayd+t4ZS3RZp6yTWtkW99TJs36CdxeiNWX+qOTSbmtWIotpgjKxpAMnKutrzvDHBOKdg5ng9
RkOY2e7cCU8Y8osfzKSqk5LnqVNVkHiJxvoo0wX0wTeWVv9bBWu+H/IjFzZQpOBSSYrwRvJDfM6B
eLSMGVVwcLq/9QY4m0nn/dU1fdaQTrOPuI1l1oKShpHqphDEGYIA9ACzQlMR/U6WiXgzmuRfu/ER
FJjQFZsoRzYpf8zjod+h9Ny8yatZ7XgvfcLb1ZeZ+Kez44m/lNvxaxcZpGE7Zwxq93V22/CIuEKj
CzpCIl2y/55F6IMhmz4MV9YnMWmmS03Y1LmJryGdV1GUDaB2Bwq8mL8BxPKXg1SQSyECZdyLCPyI
ZF1sGsFygzMpIt/kaSZSc9cCXC9VamMLxVdFgR8nScdvo8EGxNWoUrtmcP4xILISrMWV2Empj94T
3OH/OlCi6cAlUzZjDmAGF/tJWpqVLEmUybsAAlKvL6ac4ZagLYcaFXnW78movH7PkJ9Am7dcFF3K
wH6JXHljFPduMAJ1UQJJok1JLgh8EyHTkQQIja5p2Omp080c/JKIyPokQ3uR7okQ2scgNXOxy3FX
Is3n7OFpxbASRjc6M17Tw/xxt4AVjyW7ibQXE4iZSO7N02PDsvbKReOVmh5uZuAnjwv2Auv+qvH7
912wTSrsncmD6XFfrLofqffW2S0nL0IyTsMQ5kX8N8bKwhiLGEDfEij98cMfeQEykftxhtZF9LlM
6QZVYIwr2jDgBHMnJxr43DnnpD/QKb78uUxwl6ps8M4HN+psKdxkQk9tFDa28ihyua6nqPbsCiw7
HCLPox21HgJxfJJho6FZ1qtsiZqQ7hA/DakCysPlkAG+05cenhD1m1YvDHbYtA9JGecfi9wODNLn
BZoW1Bv9mY0LuElBcMIz3wqtrTBgMnCqOePV7AO4OeURb9/F34++c5KvdLPt1024ev7Lb6YQ3Hw0
sUAzYzvEnX/+BH+Lz6npmYOOxIFDklM86oZfzon3v9Rn+jNmI1hJUgyMG0jtKuxXSXOptITfLlMJ
4pw+mUDEOpCkvqz6Hst8TZU5sRxg15zJWEKojX9uKBYdZZ2S/pzoO3FRuCP7EgontwkWH8RNjRAA
M2od86wv7dcCi0uPPa2A/KI+QikTFlcdRaOpBTPk1svY4UfORyU8fPx9PqNdiGrPVqPDsb+1wovb
kXlx2vvoOoChoc3AR7c8AMnwxfsKm/RuuIHghKMAUV0omGheHBIOXY+YqIAjApPk4drKqB5eC14T
oiQWkggs4Xh8chX/WqMTqhYHAXqbnpYygA4Z3uAnQnEHxn/vAAHZNBcJI+Ohgp47JHu91XIfD1cj
2hTkHrbh1tcC5bCGPyi+qTiQh9iCSlzCnlRsUIkYd7QgLU0ZpH1/UblHEmyDK21UikFJTpi4GWLq
uaKY8D3eyun0+6C3+yR9m7+jbKOjuDHVxDO/yNRMRdyyo0d83Ytx+DfS36j4JfTgpi80drfyhzNh
dKgSLftVKO2N/UDYfTaihZWCWqMhPMApxxgtLIG4P4B3HVW/PdeQq3HrUOcpLOEonkNbD+ZwAJDe
JD1kj5GT55pTIKxdNLMcNtoDyLkvN9e3Rj1Zc7oo9o4M9XS1gzAU9bEh2v7e9zJ6D0sDesXcbrK9
BTbMgo0FEVhtsPx85b7Zl/xIiHM+nFnieR6/MCh4f9xSRFoctJ5nwyRFBnTv7+JCiTJ7IC2Vc/fz
fH0gF2BgSKHo6J6S4Z9awYMrvqTaYPixHQPymYyKSpWtpya68+oTs2gXVGcvgKZx700zRSoNxoR5
PFF+bdXercsYavpZWm4Qno0AS2nOaNDxSb2areSRCIep4vxPKKk74Z0b2sqpjT9Cox54q0upanFG
nlL3mW/u1C7D7gC4DLDnWKeMQIzRDOUxjOLIeo3/A9NFPgGyjnlFGvK0pFKCJVcyFDLPuP5Piqu1
UdiOapa0g7TCQNAr5IIRnYI7IcwBDOubskpNGx86QFh9A5Paka2po+J/IS3pC3xDSurTeD9rUmwa
yzGHYZFIbQLzwMR6O4+4OrzDdifCl9Ck1MZEUeRCZqRfr1TV7GBltPMZmRioKscTIgzHaFJcBE1M
aoh7NblKoPKMeN5OVuscJWJw1rcx9ncqQmW5Vk9ZrQLs4bRx6Be05DBmXG0as79eKhawTmxTvBpA
ZOAXq2m7LiXirzujAJ2tKZUzQSl6dn3UWfwR/LgbT7UC1uRCncvNul2qmYW1I9ZEUU+/uM+/BxhJ
jXZ05w3miCcUu6OzbmOcSD77fiYzL/8nywcl7ALAwxaIiHL8w39/t5/f/oXOQPHMbH1K3VBoCzWU
5oaovVN2zfJpi5vJ5DEDoV8B/HCfgYvPdnBZ4La0M0KKddXge1BN6M3HLLStXuvPI2KDwuHyBM37
bZqcWzPxvbppMRMFABk9DQRB8NO6OrPt8Y2dTQpOsruP0zjwh0GETT9QvX7pa3AH5Lp5GypfXiB5
zcRWz/TbhShZfT5JwuPA0RncJKdGttBK1XBGiRCwUae4GWHOE5q54H6Wyy7NeKijtcG9WFOn+s30
ID7HRJteNGabjbwSfXuj1/5Jl6+9gwyBVs51DprePHHgbZ3KNQgtrX/RZRMAp7bDAQHg54HMiKAQ
Qol0ZP4g0GjW8eWQvheMsA2rlvFsxX6DesdWHeKfe1UwjqbWXNLdM8e3Fm1H0zxSspJH/ptTVodX
7a+m8uSzdS3SGE8c4vnl1kqs8fgOLWE9SUAf3r6iH02yGvceUVs6AWzhnTs8Vm+L/TtWKni+gSWD
fx8VXtNfqJlwgvtZqoZB2PzTqiwmL41oU6eTQCfc+fB5tlOqTmVBTzpmlq3WSZC5/SEDNqMIKziM
VOGIXb5s0A1lspksHc3xvooXffrh7uDSIxAH4XeqR7jr4asH7AIxDAjisB32cQCaE80u1nQ4JwJX
m3Xuj2m9wFZNODsIf1V/SUr3S/zyvVrKgm/36lQIKnuHQ5LHLF26UWvcSGRgoMJR1Ky50mgyIhW4
VoRYCUeYt+G92+tawZv4CY0GYg4UDXIl2GUR2uLoanLikEEvqV0PC9t2HO2NXBlYUw490Jl/7g28
rjJdQNifP/eX2NVgAUB/i1VbkrVXvgwRPzolPF+drcGOmngToPWnrvrIm5VGRMD671CbJjteimRf
M8NAlAxu4XoIDH6kjNDzuKxZpg8ePY3KqZNHGH1N2mVB9pr/9qtLqEHl7b+5OsD9KGPlHT5wfi6w
0fDn33i85YIehalE0U82i9WYq5tmG3hyc9F8bD4lhxt58LZGcCZDVMJNBJ6Pa7dzGI/x8EKCsVo9
TPxazj3uC0E1zAovGWoi3JuXGvBmazDpiliqO1+w/d4nNwmy07ELl5+bFGe9LllIvXqYIhDM7SBh
khEx1ls7mh4lXicSEe4LahTZZrlvg6jpjJFJYl2/izjgGShUNJerUhkfl11PpbiyMFoA/j+uBPGX
JslU3nYazFGurEJVbZ/U2vUndUUtWj5XoW7k2QfDswZ9kOk8EY8gVupnGBAVjKGTJ34VyQRB81x6
14DZEn0+d6QIvLSEtuXOlKZ9YEJVH7rZLIA76kpck4iDnd/u1vXT8CLW/g81YlKFKmM6f+8wH0rD
tAi4ZI/C0lYXLT1htFkgU/8RvKMW2Ga40pVJA5jc1JXORLlFR/sUq4kawpflQ5ozl1vhsHVuQCb4
EWN2tlf+rrjLe65++ZcLfluFa6A9uiebce1gE+xKBh/+FFpRHQGsTM7v/OoinV9iFswEUGEfLduY
HyE1E5LU6OwZqKMw4cphgps1T9b14dDM9CQe6E5fr2zH3SgPaSmO80RtaXOYTQR+xpjdjVJUkPM+
BRtPa38EWL37GUelMxkRBg9yB6JOiA6OrWCXTqO58h4p4T+/aiEtbRNJZLX8BSl/4Ud07RX9NJD6
EFli3Ih+lo7UGvq3GniqZ6PhPYz1vY5TDJ8IKPYdy05VHuMoNDDcKKE5cN3FBxJqjkaH3FnuCMrI
3jegmv9OfRzcN4tKt8b5B1KRihmYUVrHzjHaDGRDixVrDAAN/LqcdTs8+9Vod1nhNh9MKOHpE6lc
FL1cPvFKyS/oBjj/cvvSACjYHpKpl+ZfNygHt7/0VqitYpE53az4cp+JJIoXh6c/kEaJHZkYyel2
ZU64bhjJwYKVo46RzaDg8+WqLLlYikGWudVBFp6FqVRnMnwYsBXGtZTs2sVfs+96xUv3jgbHkyfb
hyaqet7N/IWnn0fgA3L9HV1z9tmuLyMr2CtJKzkFJfkUlyC5nfK9CHEzja5UUrfjLsec0KEOHpbm
/L1ExtJJNJ9Y45DU6ZSBXUiSpmNix6L30pi5nI+1j2x4vADD7F2AJSG7d1DA/4tsP23wwpRTx+6K
kAHaEEK+ibIDG7X1BykM2V4jXmwOWjF5djbyFVkdZb6Ve/e7zp8j104BXXflDslKosRTyPSSZjIb
M1/YveF/e5MUxPKeJakWlWuhAeBRoXV7YLu+AY4RLUUTA/JTktU0y/sUI74jDjg/9FplJd8IfZhi
n7dSG8oqavg6IGQV19OlqBjyfYfljPRqFDAfJwV+vH81ZUSoLmJokFTlYpURGsNu4jlk0K7BIolf
dXN3KOAiqgmi/gy550DTqcjS4I05Ii7c3ltg91JEaV9y4bkXeHqtPMDGf7JoEDMhbd25aYeThYrU
l7BejqKkt5qO6PuoUeofmq9bZUVcC8Ia7WRCxGCqOmSJ1Gve5F+/wltWExEn10gpfxTPtQXRAJ4N
UNGzilO+UA3yK1Zp1YL3t2XXPc9d0aLBa8VtrZ4bVobswe5b1KMkvR6EvDQoLUAkzWDimFFU47n6
ARKD8zEF6ihLiXgOmeFiGEIWeJDiyG5yRAUhzpreEgZtK0mAHmwDA3bW65UnVtWIJ3BER7CR3DGD
jLIqI98HyXa+ARzxT5tT65TP4mZiKm6dKY9VYNjLBVpXgrzL0iy/Hs5b34vWXiSZY7urzUZP47BV
9CO0BHiLlsVQhorc3WbQEk4f43txoXUbyptv64mAsHeCHJxENoKkCZYjIICUuvecxr5FXCJT7f05
SqXn29Xvc/mBTDvc8yOqAB5KmJQE+yLP5lbmad9WbnoSP26Ub/mCtL8XYPtXnDAl6gwF/syMDuEf
rPXXY4UWjKFdEFbPETv/6ukFvAaH8kjeLgdDx5KqOA0JooHa7vI+NLW7Ca71F5KnjLF0rQEi3fX2
ol4Us6eimVJ+mLHk+0pcQeLpfbuRclZ4O311M0D4zsUlxrY2Kmy7OSSc18uil+IAoNbzKg0Cw75U
SD1QUFT9s5bSBVPDsyg9zRxi+JQV+dsaWMCD56VDW/3b/7z+XLaNn020ZngdE44xyDgxE+gmQOT7
lWxrlMV+v+lDgkgKvbaUPNg4Bp302GJasJclkVKqDfc4/pqzvf1YO+bKnUmYIaP93BAdpb6WdypS
Xm6UVlVreOpGDM9mNmQBwhfZENXCmeasqj30o2Jt+BrUt+Rhu8mHrFBIQW7+oIL5oeJ+JqYjbW3e
/dksHFoZYlBWHSdN/ypwMTP4sUJe50q86kJ1K2og2GLkcXstYtM1fP06wDl81J4Z7bdrAFCDBFol
ID/ev6QWnLdNx9/Dw1C+wnY/V1IJkCJqBWJeB+W3RiPAPWOFePZjGZ3BhuflBHEtdUukeIADJScw
MIeqrpuKYxXhVXK3QIxFCKmY1tzDfo80ik5/YyOzyWxhALlwPs8JbKV5VYZfQnOIMFzQGPF0Zsiq
DfDz1DUWvqgYSJZ7Nu1QBfxWf9TKntXPVVj4Ss8ikaty7tPQl/KqwTthSAxLZG/Tv9p65aP9r5vU
ti2XzxIb/uoJElWpu2MBecdJ4FmkXEdhWTWK6xc7eHc30khQI/ZyY8oNZeqBCELn58bJywqlbWoX
530zHCWAy2CFs+76pcYlZbaT8V/4UGhb+itmIdWWcGEtQqUmg9Jfdqq4uJAQqz827tiT18kiuRdV
PBPqjIdC18yNprNjnvGu8DAIbMkLWQ9xEFDbnwPeZ8QA+Awz+Otws/8lonLe4GKdAqcNX/qdD7CF
HuHhC1ZiC7hhRW8X3nutVvFAxamdm2Ha1ia5Hexcp2xF+Z5COnlTJlrdB4iy/2s2thVLGoL+BI2X
x5urVx84xtqwZQDVUUc2aNt/Q41xi3FI+6n/26F/C0LeioqOCtvlAW2co50zdmFyerwTLTpcP4Kr
O5KApgs5j6qr3+bZ2bhyW8kGd3mwjUKInrAWkwdiqIb3IfERIOU/5Yh8AQTCYpKY0iOOsr3EaPkV
Lr/FChVZTxj7r8IKSIv4osYHncDDLWVZ4YlX03462K8Gbk5Bih2JktmJtNy+AcdcjGOJ89hjil6r
zTk6VT4q3a2q7xE0X/ISgpnJRrFZ0SELlsMkbKFPknStLD7b87CJb0/1PC5tGAj7Hj61cNGJ7PWO
LRDyEDHCMWAPsqO/VTolxW8YB3QAzSzHlEctpgt5/8JWFdpICmd7pko/E9opho1LcLp+E08U9rzp
NEfaqnuCH/Vq88PXyScV2Sp2wFHzaaBWwo4gqdQdFVuP4Cckx37/8khDImbS2VzSMPjpwSFY17VU
hZit6yfKXtEficy4eFWLXgYE+0a4B2l94MyS3zfMRrXwYzR/WF3O0bVuHdwgMtaPgH9i5Q/tZOVB
UeMWht+mqikPwdrrhXJmZhe/E6AhVGi8DuDOPE5ofVQnpN0ST8hojhjOHMdfu/hFlfyiRBi9v6TE
EHHZF84QeV/fTBl3uv0f3xVoTQWGAUOpTTD3qDTuKWxOroE/f90IAHZKZ6qmCbpdBjQMz3FHhHbV
PUXsBymX5RmpeevAQx1m8hVHBiH4UwQ43ZXsHplbYmF6MvE02TcUpxOF9j9KMJenG/WDI8j49/Pn
P+BhrG0hfbdXdM2VKv0yt7eKVdGTmsyq58mqu4bgjqogoItcsXeUSsZ37lw92t09y9WJfiL61ZHL
fTEZLm3lqHc5SDFdJmgYTvApKcHo7tnpeQ2H4gnmBQWNR7/AjnwZQBVvZ7v546YErNSwL1O6N/dd
Xy+alMzJBhbZXqAuW/PNA3JhA3pB3f87i2m+MUf7k5T1S7VxFNTOtiB8SPjdopOkSQToVaymvQsl
WuItej9RIAP8oAwKLETvE2Ut3mrDtWHwMbJtkouG8ubbE+SW5vxT41h+kvfKpdtudkSCey8T8edK
giKFtUaT/5asy5dgmHFfKvZtI8We8sAD6JAUfd+H9tv043biveNWnkabw75G5keR9dutlF9Gb+Fv
lyhpU+oJOibHJ/7kO6nGSzDSm4Bsk3QPU6/SFjsHzrnCBxSBsu+nzXsbbrCbDw4zA6oRsrB0KCgw
3UBjNY0H3QLRV/VmuPCi/kmd63QZu1zDe5cIrWhPCeuOvxUfo3x6rdLhy8Po5fLDSidjh1jL6HjR
qMzSTSyskeqkO1TKBzDv46Q4Taq+AgCoPiJeOcH2hqYkg2O5EnpzpY2NYPO7SY3ufEBYebeEfPOG
Im8mmSOztIJkFCHG8UppMZeX778Kls8mqQECUEYLt/YQpIXlAc8elrdAVocNHzNk4e2MSPgSAGKn
/7dlZ6FjYthAIAyN37VUvaoyFv8E594c8AEHzcr6J2/pGcLLJn6v9z5k+0SiZTDj2pUDn4ZI9UZ3
9MiaWVj9A0kAUUgHK0ku0DzgpI/pqJaZ0Lx7Nb+gH8WVUaG2lAUdEPLnYFZkK1Zbcv9Vog==
`pragma protect end_protected
