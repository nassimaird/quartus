// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
djU8TwRwnRXe63oqiqqKeh0q5X7hq2nrg5YfMrTBwf2zbdabMW6jQPDEKQP/0tnUxzhdbyn0e/UM
jY0grtOMSE6Ilzfpu5Deam0evkxD4Qwo4SBqiYjTqF9PZeA7rZk1fSFfukQeKytBMwQjH3ZzD+Jq
/UX+8BrEzDTm/aHRae/RQCnVR2nX6yNHTS+HdWQItGi0kiWMP+tOZuy21JMrrUoRMcsk3RWCQN/o
chO5KgxM3OVPIXsM6Aa2Uy0k6Gx9ycHiufUW97ZcAyMhC5y76QRWDz10U0i0NknFLI/bSawRIcjL
nRujAGAiUPndmopluQfwYkxJY7EAxK7M9BiLsg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 39136)
Pw0cgKmrSCFTwXtSRUqo4kYuuFZDXwIb3mGrr0i1SIxQzj21yU4Bwkr4h8OkIoR6P51FHTqJRPQs
dPRnAfXYdkQZwae9lKvbcRBExRCRmavCGmA0hmkJJZszI7RGZ1xqMg8/JSvvEksxmPIS+3BpJI10
BwaND1b9VfCJ4w0Eup3/p/tuCwbnhQ+dGo7kwiWut7fGP+/jJtJqO1kwc8PZ4bFzg9PwlC6FIUIo
n1T+33DDAlmQbvN0dcECXP+1YHTLKDOqTZjYCh562ZFmrTftDZIzLqHehC3sfPZbk0kL5lYqLVWi
VDBNYTIndg5T37TRttk8Mon8a77ueEbvLm+EvopodNP/WZYEZNiBKOaj0FIYPuy94gULWD6StJnY
qrSmt2sdWC8WsuvzUs2qxh3lGLSIq8Usk6qXSYUOe24zL/YQv+c2pPnvwemU5chYJJ5z4O106uTi
y2SHfDJjS2ghMtP4L7UeslEPxZHVD7Xs46gFD9KqvUHiCKFHSzShqCLjSQ/e70A04a4Jx1w5tC84
7kJlUcezYL3Bkx5Ec+7lK7XH81e2N4wjDY+MhxZw7sTYYo2/OYtJoaY+OAxsg8WZBXabqk23m+cX
nxgf64XUnMpknS3cU+NDWcQeVh6NhY4uaxsht7dOzFXzTMR7sCZVoeZGPNMj6Uc8i7pgswVGpnpn
J22OJ9XUxPT5xoeVozIVbC32FyQXiyV5gysBST3sEEjY6CXDAHzt2CRaS+dJQyjMlWlBsd/r3Bqb
uj9S0CX7+MjUKdOr/pVLGUQst8H+hbJikpsPtMwHMF4oCzv9nJ1qOJGUorcYtSVaCI78VXiJD3Qk
YaIaZdmh3jBQpyATh7eTw9J8o/Q/XZE0HzTHsoPLfiUilpoLwRp7U3KqkzvkcKJLZysw9mte5IO9
nCJLgRneA+brNxznSu4FaQS2AKleOZrkJmHVNrJgExSvo5sPEafqHBx9J2UfPExdaUfRos7vyJ8h
bJwqiI9SSEgwFQZXqplGGikIqUQ9shqXcs618cYVAagFDhtIxcW+ImX/Kd6/WUfqjJWSy7rPUZxP
7McYmzWjRleIlujitseZ5d5p9RKFQRAI1waJHccpGt/r9RHaEabxRk9Z69eMUQD3sBeZ6V2MmvGA
sY2p5Ybu+UIBYyfRuk/Rzq3MhnJ6DUPezx/O4sdtEWXaGvua4gt9Mjc//z2Bm1XPYzhAwqpGw/vz
EhBwmzFUCq2jCpd2gmc0S3/WqdvVy9A6FDOnyJwfz2NEA5puOlU7Kqi3gqkB3HQk5xP6OneZsGuj
U6GYdkLI11tbmMu34r2emuusNyyIAXi4FxKr8BbMWUUgrtzZFs/X/E7UwTTqcfVwFv/eM8uKehNz
0rQsietRAr/iU3Z54oDew5e9iBpxJ2X5yTfIj8BCvSUTITmiUwe9gzoG5yfWP6haJZS+TD+RZ3dd
psv5INdQpI5knr6MTZdwWDVnYyAqVBqAe/jhQNs8wkr6bBTSVBpWhki1Nvl9TvpguGGatoUgtGMx
cFcL3TbHS8apVXVgpqzNKPo6k3yAPl/3Kd9rs25pGq6dszeqFi8XcWRnmLtBIEvHRiO6BAKEBg5V
SuluxToWODyKi+mUeVa7LeHk5yywjC0MxPaFVuGZFFyxa9fcKw9H4E/LxJlf0LJqopM7v/d1bd+M
kNYOgGD5Qym0Ai4cMMvqxIm9iugqNmNDaBzIns0v74vjAoLB2YnXnbIxt/fTQcaDwW0wJAT7DUZ6
AWvyXKR5Bw1fe1+hfvkXTXFPtyykycTZUP9COtf8Rr9RC4s4yz84QRVVGpvVMa/6Vj5rm9yXIf7S
VS/XS2pGppBE6sFzxqX4NSItrsS00i07lukQhsZvplvdyswvyGY03Oke3Imx7r5Hknva8uMO/CjB
UyEULa3NufN+CQJvjMluilPMNMWFL8UgKlb3dG/tKnLZbkQIzr+LuQhjod2QbdhLK5sSJhSH6Gfr
7H+EglsAotNb7vhy7t8Ubj0mforzvytYYCzsA/mGYPICkDWWWzoN8dutGfqoASGgosnU61UhsUBr
ZWkH8D5j4NnOSvq8f5b1IWtABedjijNSQxsqHY/k1cVn3lpMoKl+yCZUSUOTudF+56cGhb4aRhvh
G8Dr3b4pVXM8P0mYRhZ9AQsUkw6LggaH8H8SfVUMJmOtDc+P4aloO1IvyZBE7DsEoRNyVcpnblav
SptdNzxMmDxUaZpZ5h0KqdBAeOj9oCfJrtzz/WgEF6lmbv+7tfjiB7tJkt13SXYm5+acZKlOh4EJ
4WF8RMqsBrTYOBAM76w7Y1hNHxRmA9NEKG+uNTRdAKFvb+hIExsTMbwXvj13yRVnyCecvy8n0605
ddh5nZIsrfWpmbX4Zngczkz7JJVcoD18gH1dmWkajyNMlZYUJ/Ya7TwM6nYX1HYjYeKaBkfVIs7i
7fMQ5BAiZuOs/8EBqOJBIwrPPyGwn1iNPk4CLBzUhDmk4iW/xKtWYL2muE5ffM+BKRWkmP2CYGIX
eqKXULRdY/jXR9BGBMlb6xgWQdaYoYlNlsmt7hCWVdsQGtNVeAlIeBVxF90mqAMf/zr+MQB73/ex
Vwi6Tx8ArEYjOEijh0QexixSRzAWhks6GL5guUXSwOxL05Xvz6Yz9ORrgyN7+F8i4MN5ifj9RYEN
IuvEYkBg+ibLRQL3+wSvpSK2DS27ljJB0VIW1EwtiX1nRI33t0KQBxADSNoFf0rLliUpZLC3V5y/
BH2pfMcbhPRJrptHP0+4VpINaREll/KVHGJgQn+OYQsCDXsydfP1gbtW4zc18U9SpAmjHJ3c7obG
24mTDsiuiz8Oi/es9lyxhgTxC9+0CPB1ivmgbw6DQlDWAXLSWlhWbywnhF5QfZrDEyUFZAfB5UvD
N7kDt7svC8gyttzq54e0OlSizVoJDJVSmwunkxpDVnJZZaG1b9YZpI7/dG2s5sfhrvcginGRDoUU
N+Xq1wTkCLLWI6erRw9NJGCo7Lv3pfcqR1A+71oRV8/Nj7lUH4CI3Me0Gy6VrgPa7dXa+3GwHQab
yC/p26DMy4LoooEn3t79rYnpoUNA9Jw6heC1a3YSuMJYKFRDXQhAoC16nfSmBgqZ574/Hl2s8Lrp
V3HAjzdizN0ZM4lc7DYqK4GIZzD1+pybDkMah9kaWiFrCHvqQtrpSdk8mqqKJVqfWmkL6aEiwf2W
gkWUdoVsYoweMKlS4z6MBbwTBqVv8ZGJovCGsy04a74Ic1pvD2pt+OMIv69w1b8v552u0BqbFMgN
Ue+cP9hcpk2FmSfumAGeSBrM65gV+2TW84Fx+3aciZTSlQH35fzIbWwuVAZZDmNizIvoytc4XD68
YzN1KK/RpCHRh2z1BuYDED/UcgAOxeR/LhVs9ZYflgLswiKNzI+YzKlNQAqBGgKQB4fsgWjxDnp8
tlj53iBEPlTSb/ttvHouSpn12hjAssqYE6BfnO+vAb9qt5v2KifKWaSKKkKMbfJS52lan8JEawtT
ZT3rq9ETZq9p8/5JjPmrAztCcVV/0KyCVMeY+bAMwFQdotJrDUnolAFxEmC+N2KlzqgjqDJrzZTo
wnT8BzdCs/LCc7JNUJBrV+kpOYmPCsEb6QXaBrMEHDCAw48Z2bdLFTudlY9EU0XtIy/wrYBFGW5r
fhTqnM/jdUrNsJv/04r8urU52Xdg4fLzTeeQU9nAyE078h90T0rMKAwb2MNMuc3NLFbAEpgldOSp
boVTwl3M2Yrm8Nuxv+vZihqSHi2hBWcQzenB1yov1p3uP2TyqusDvRXd0ufTza+YFLC6fgQybhUj
9t5xn805o32qAI2DV141Ux+pRt9yfL53rSzaeeq+74l/ATkvW8ms3xb0AztgU4sHIcWcXYT5Z8mZ
gwwxLS2W/0RxytyNmFIJ3sZF0T6cfH0UDAFKraVfaV5GkiuIUzNSugNW8n55+eoqJOD9J75tdMJM
GqrItiavY0O5LbZGNOZrQoe4X8ETBXvMo0+pdeXCM/meQLJzvILMt60OULhAaf20jJc+VDY2deTH
6o4yefXzSpfFVEdGn6Sa0cgAkOKWdHhTnOXgilYMBOdS1zBGSlAMv4RBtDXRycG9Ckx00G3R/Rbg
LOupoF2KTuNgsthqWn7VCfbL2Kue9+99j93ZJiSedUXZz0q+htfNdaRHEZiw+8CHyBLEhbrSK+cn
zhElFGvxaIsif92AOAHOpp9l33QPb4vKwLykBOKZZmda4Ykr4DHiKcO38z780jxea+lvWQ3FK3+F
S5YvMKtrB4Ul8FAKyOVfWNTYZDeEVhN17gqlSFwWNQLHSTg0xLwf021yPHfsBkjAar4Bsb56BKBV
Z69E/tJz4UAGCIxWj8t+NuCbEQVMmK+cb9vjkbAnbOF6gc9gSkKA0z5ESHkv1wIbLB20Bw8SN4Mi
AYlMXeVuvjH3ZAzLPMgRjc48NeQoYWLMsLq5EwoUHRRM0/syb646dsy88iaixXVgEbWTOzqovHMT
qvLD5Cd5QxRWJiSbrlFywmWrmpNuhzejL6/uvbMWqpytMc5XIQCw3XeZhVevJ22sKpJEzMin+2RR
jJOTsspSepNaQCC3v0uNHSkHTq5ShhH5glS2qEbrqDwGHgGeLe1KNeLGwELGNA2Lxg63N+hqABX0
mk9Uswz+9XES9/n5GVuzEUpIyU36LfhE8hT0f4giORjXPAZB06n3ucVgr8kL4AIfRkeeqmuYX+qF
MIBKT1qcRgwvxFpBXFPcyEfFJjfDZtCTyloAiYN3MU75m0CCtjAbMRBfQf9lqjJbTlwWvYyF0LkT
CfQkD/C3d3MDykJ/Fy1y9BDQH9sVg98tQVQ4yc7s2t+MbSShHHXrpcuvoprgFj13FG54TjxTpFhB
0wBCZk5gstTf8sZgIJSW4GlgSc22/Z3G1sB3i/RnjhnLIrNEkP+0DzwRmIDEcbTHagKwYmH5bUjD
q3ooDmCor2vShShTXiHXfP9L12cTQ9YmcC4KEq+3ffncfNYJfOWPsB5EeiZGsRdagMwpLnVuxHi4
9m4ofC15OJBkQKe76ARbKG+V8cSalwaNBa6Xexuh3r9uJmF4kSy+fW1PyNjdSyDjHzaWyBWdV2kp
RjX2Ta5zaIKx3f1WrSXR/7DojE0zSfCO73hgwv0hztliahL5ipWd21xkO8NhAKvxawFs4b2zvrvC
ZEVuoy2tfRJ/iD6YHhm7MNwq/rtXk8oHDR4nOkO8IuTVpV0bK47jnxfE1gt4JTQ7y3wLqI+Xgcks
2FoVeJH8lVw4nTwrNiDaYAODSzP/SqALyICRVkau6f3EO6QNTo1cpD0a7uNwxLDCA7LlD1ZRtcIc
Nes3kQcvLILxstU26I8njkMa+QKtHSxGdjGHcZbr68/40hlJPo6v1dyA9brV6ycDHziAg1nFDfT7
XkhanLX6d66BnKZM/byZmdX1QcX618d+UODrZxWLAeHLdWdRw1hOcDo6lQrdMPtg9RxJt1KU9tv5
fGpizQtyAiHLvv27CRCqc7dfYukYeFIYh+H3i4+5PlxIAALNTpuqftv4PA5cUN+M81ARQqIDj6im
gcbtwz9AXtMfSvBTPjQ5/lVBLdtzzld5F7YNcOq2Yo9W0WiAuuAksff+VwagxLNVL5x8/XK+IBPs
C+GuJqDt2TMElSaXy+Vo2ff99YAwDHPwNdDOq0AOSG+wdf7uipOeSUXMMQahXJHTXjFkOkyzWG+h
54VDW906IKLN1xhXAQ3uWvs5Bip/Wrvy3i1xpM1Zh20QLvBFouX069XrqKYk/si50rfupWOrP1od
NbySF14X0uEiiZfQk+zPu9zLU//drnc8Fcdjf/RqHH6NJV227CN2I8INbl2WR4dzOtok/99eIUdO
eU6s9wjSVySv9d8F8ig0KfK+RjwcjmIsAAAS6PckocV290AF8uRikxLSPg+lv8l0+QklpBQb+gZY
bjmb2RST+EhEnbfAi2t7mvp1cxkHOf1YytbUKfrExVWpSWRiNQeXpEVldokGWBbyeEBcMTmjXF62
7JRdHykbIpnpryPpnQc7DWhETAQMTjtNh1TUnVrvgy0XKKkiXTOa868snhcEv9ZjdY53vhAi5b1O
zuEAAno2ziM/qeTrddi0QlPwneBBCGUU707CvjRdgF2hGrv9sXU7edHdpuI5eVVpW3E/ym/53UAP
FGxYjtH4BEMINu8wtOmHso/xppf7821/6Bn315VAmHtl6rqWJghTsKy2NMlPSCr38c5lUjnExZxn
CSZvq96c9qfmKt1vps2yNzEABPkwEYq2z8584/CD7S0/iywvN5ZOlpU8iZVAienWu7cezvaNd2s5
k5AGuFQQVrvsV3JgH3qZGgsDVSqFP/H2W4lDe9VeXUw/l5MwEqrHu5meWvc7sMl815ybMTXjmAs7
hIhW+eIalK6KHyX2t1MPz7u+U5JbOhh6tjideUoD0hgWxu2yZKFaC9+q4RRgZKh462PKN2VH4VU2
Qk+/u8TqHzEsGs/nRjGCQ7yuPSIDxgPcnq3QPKPAr0vAbSDhgJu1ABHnOEdTKBrpzIlOBCxmShCR
o1Ce8jGbNoREnOZFhlR4kelSjqoN+LmvGhrRLTNO9cFUO11cse8DIyvGESZgZTDTc8duCozu+8oY
H6gAwcbpKeYfYPFNGMreZrrDazNrVnjDYfC8nAyq9ja9q9xUcGMUXP058FC36iw3fnhR8HtOt2/7
Vclqv172ZEfI08VFO3wlTQGLzQEtSaJD3xrB1cm1H3rYKlrWBthrqk/7o5R/NSd0/ArF/WsVLBOz
D9jw/go/6kymnh8Rws3OFrZaMZW1W5LsZTu7RQ3aLsvD+dhPRVyslQHXPTcmN3XtlvaHsgIXxp/7
syUlNPmvLjnaGcC//7o22fbrmUn+Nb/Pml6dq+lYFaD0VpFhqOGClHHmaeJ56F+k+OsDLLwgHmhc
3tKuZ+M/dL4+lp1m1L9yAHygijmIqv644LyVHzrf1qxHtJw+EteWfHroIMPQC45l1oQFN978Kftp
BAJS+qcnYaupaUdE/Y/619pvugkq8VSj/e8iviPJYxfiY0J3tjYutpFa947rmr9MWckJW7eQQwD4
YhZ7TEEPdcnbR++/5A4KQufqsdknnsWg7hFFRDn9Ec2Vh77QC32Py6CJPlrEAJK8WhIUXA1+lanu
Dw7SkYpIn+QuqzlembpSFf8TFxPmCx+wDM3oATGX/WISqeO3kBrCF7n/JLCEtDLTD6j5VXaHtKm2
0pPAuxsyriaFtQ9v55FC0JDFYoLFfHkfFU2JIefM2A1zBX78nEJOJ3QUjP4LQTfG3uAWCiTjDeqU
xLdF2lA+qcVpOstC3f1yLvRTQ89pIoGjPXDlsBYDjaeTr/6CvQ3ocuZgoRf7ZCiolubYYQKStxZf
p9IppdZrZuqBd8pjfqiCG4z4VayWFCHhE1rPc0MKxOxS2yx7JrFxRHBde1zvzoEy6FN9vfVW4lqK
v3f07OXSytDiRRd2GXpF4oRP+kJ6hUhY4nIx+G75M1kdwxbez5V+l6Fp/alJSeEL9PruPAm7p7eo
CAW+qBB9sIbNSI3yLvCLMixAQ/XshBL0/pf62zB1z/iCQGi8cle/dzwA6xis25kTBcRuowYXCrLJ
nP+YUzyc9B3dCsHUOynPuwbqCxbvuLouJqNSoIyQzxPPuhwD8Ce/h6Y4vQVZOksXFSxjyllRGV+O
lDKIe/Z5dmjsYLuSGe9qnLqz3I21UF2zZTyuH5lHR8RtkL+AsWIS8M+C3ar+XiMcekeDnrzX6Qys
oAKbnEWegxKpk6rQ3j8fxedCUFQOP/eH1Cieh1qRDcq25S7J9Z/VIWOdnE+2DEDzEXIO0M5wP3RE
saBZ8GYEcuTRVO+bhr45vNteNXrdIj/GDuWRP67RpYROE6tB2eboVRnZZ62eah76dOhWHwHdKGcj
IzxwF+6w3TBgZwxoie0Qi46bNxzz5s9VSqartBZpjwTz7LuK4YbeF93hSyWLvvzwsT0mnEcTZSpH
KQpjG9KIQe5djoyG3RtBzpGYJC/xb/YtzKSaStDA6++BtYq77GtNmtyfkZWgraC/c/fxPgPnz8gV
+VI0ixS4OKuq5UoM13pkAfH1BYJ92Zd5RP9HR2oO/6KYE/AQkciu+1oNd7UyC4ySNneIkXBY1wjQ
3IH1WxtIPS7ivj4c3JVpIxxzwyrrwxR/QjbTgBHBHNg6ghZtwTBKNpzVdLTBJ7Z9xz033MTSNL0p
QmibdTDWIDvDTpdmzCs2DD82ryLuBKfcTE5gI/N27hmW8NOd/FHEKU6gCHDDOlMRn8XQoXaQZ/Lc
ekr9JhmDZ2hAbrvjYxs3LZpXZQNHxUOInLWGzlPEP4yGXGCyXuRDWhPbPdnfMmsJrkU6UJLBScjT
8t1ItdtuQvXPEdOT+JNa0Zq73FZTcWdCt4suMdM6fpiVIzvfboifuqJS+CsCNBiqw8MPfrpvPtz4
0BBSG8N4u6emxjf3k1bcltEeQdrJh5SHv5ziQ2CoRqNlQg6bsoEyd5EvDmLELkDDxnzYq/dceZaF
Dn6bEo6w8jF5lzjmIL+pjWM4kzeOGYhXTzYZVNzt0cViQo4Qe4Ywe0+zw7Eb9E9OHCNNy4Zos11R
kqDXATOCoy91Wzl3rDPnRTpg7GHWm4QUJ3YcC6WM3XXbCR0iQ8QMo3DAsMamixmodxWMX7QpwldA
lpgaUGRq63rIaw4mIRQC+7PRLFu6IvoWkybVaTx5lfAcwcrd7tLEPHay0j9mLs9zx/Gpz2WuqMHm
xD6OkYjgAh9YFYIrVErpr0CsGuxXDVA2S9zvKcxOaXcsbGdJ2yultrBlrwUzm8r9yPkGeYfphIQR
LCVbiNjZgvS6EerhvTNRaQV8Ke5A/+LVefHYpzzP6VVPXxKLU2WfE8bxWzlDDArWkpfMRiBvRVaA
ZGzZ6/ZwsYjdKAlauAfDxeuv3WsjMk8mMVn9JkihgxHjVvUSmSjcc1bIx4bUFT3G7ZWuS/edNszJ
p6gnJ3TeDOS+qW2GRoeDBQTeekRdCqUh9okFqQVkt2DN49JbdYMhMDVPH0Cy2z1IdIT5/8LBvPP9
6uiTk0w8AWHV9j7+Z/YWjkuxsSCB5rtBjlf0ruySb7iJTwgyOV+mf7P7iMsq/aab4yw95ehmUXAs
i4cNbKGjmMxs+GJtKE3JYQTJltIXm+ae6o96mB1NF0HmmgA34RpLA4SvjXyQ1vK0lkUHs3/48lyq
6gR2qSGikCGhVmO+DGuHVz8lkwbw7QOpptdO9xIzH4nn0twH4RxN932l54+YMIBeR7UyD+9bm/6d
qQ6iN2BRAZsL4YrQNCkAIwzv9TSXqAf9heeJYDi72UBSrX3Zi97zbkp3NPFQgC9bgSfDKMbKG3ra
Hlc+KFnEkEM6BNMI5JJLnfyJM8+Pe/f+GNHge04qt992CQD81iy5+TVDnutsFx3wdRHa592dojC1
VSlxx9BWY5S52dBtif6eVoFuTefN+0MSIoGaA2kdZRF5x+WJW7bR9kPuTHh2UKcqlVn14d3xl8qb
DhT6CnvG5nE5Tgm7fqWSSkpGyt96ZVSodzt3HDTyk/ARVKzbEoyyTO//8Mefz//Xqg5YexC2HPvR
723lCWyY0kj6Un9GPpkhfcktAzQSidHbnfe5iz5rO/oVxC/99+xclOyg0HhLYCnDD+MZSWCt69zV
qw006UkJXUKw6d09yEitOBdWWwRY2WZQGWg0NWo7Y2jUSgp02ljE8hVDXGINce26oURxPzCv8nES
BTgWpuDOvlwp+/PNBLyo57umxQsfMT6MbnTIm+Mf+3mI/qmY79cnykM7Coaioqc14FU1Igcue0WA
55BiBuHPBl8fBt7ot+ut89UBQTybmgByK40SugqPUNmt+QNcZPAxwZ4vV1c3U66P0jiWxoLRu+Ob
S6Lkio9VlEL+sj0MZsfIEaQcoW3OBeRY4VPXCLoHXiBlLBukNNtpvf8CT0vog2zz7TIPvsKie6M3
0E2oi85GQCWkS1o4RszQxdVrecL/dMqJzBHPF7WXKJn9d2dNTQPJoOS6Nixh//PI7RlJinjKrFMo
uWVGu43idTSaMVKfQHZL+jl4dBlUp7GXMEZ0Cxl/u4pCdqtRiIXf7WZWDNRLUfIjPA+3FFzCMBxj
Fg71r33oXycdXuyMyKouTVEsk5YD7+aysMAfCKD6Aso4DQ1BIib+r7Ae5CT/Um6o6x6SxUhuf5Ni
B2wPl28XZt0fg0K44dmbfQZ65E5vW46FgyrCTmdqnVmdSPI9UUyNJFV6zYAuXNL+xMcYhnmzxZBF
s0hrbF0vBlbobNXXM4AITfF0lBV/efByxo4ZWHDlTvKrum+LjiCEtyAlTlosiERAJ+9f5F+GSmKo
xkfWYQHrKVhCyv3jlPzR2pn07vssCvRGmhVu5YEIZRfpB20IfGwxja3lYzU3eX+dxmNRA9560evb
g7ZAz6iPKCszmlWdT2vPlDbAlhaSpFMYWCJe8/wlYjrmGqryn3JpELE10H3WNWb62xQCS8i4KWx3
mfBBXF3O3iNRS1wxhusnygi9O2rAAEkwDFz8/+vukmvGnwFPPEVfgdO3VVaLnBs8FArwC3Fk8vOe
B9A8LSAblcnMhs9phIxrcNDlmLskWFR+13rvJd+3IUs8wzovhc/HsMWMl1Wa6eVXAC5IRJmlSjvB
V4BABjHTdwuMyX8Q9zRNSPJl3Sf0iBTUgBixeT3pqpbZfssXoWVuoQtLZlkGMdT/0u4CxMzELHSW
8pQ3Yx+XaSs+hsoCJe3CBOS0GYIyaYgBa6TOI3WjVRwyLBjjGszTrcREM4xFyePeNzTQcqpfVUof
xvnrJ2GbmXH1dgMBwJDLe3CYvpJwJJNujeCtVILsf7asICdUPWlK4NhkDRbjy2AXmkd/Lj1abyYJ
2h/+rQzVMShQvjrKaYo3LqPOBYsyIHQ3vhylAfm7S5o5zWp8s/Ajh7FFoOtXC2EKssHQhl/NJqQ/
bcD7+7jWQRgu3RICq6HY8NiIrNV2Tw5xAdxsRBJ3abtFdazbUsBaEiVqw5g0zljm9EqVXot/fUFX
jTT+aGhb5lxMKi+TotJ57n9otK+GulI1cXkYe6YxysYDDNoV0AeKEd8Gt+Hrb5nGIHkDMiRLUPI1
MowP9hmK8gQpFE4uZN8Tk0rtmJHZJ1Vlo1aJqYcqgjlUgIPjF68rx4fRQpq3LSXLXtPSY3MMSMeI
he6stSnl4JQ8rCZdiT7FeuIUUCod/qvFmehsApi9pacyZ4nMfnUlAqQDeXagg73oSnBwrRLz87bZ
l/s5uoVvKY4i+nRSDydKG96Eke1rQURvLyR1rigm3pqTHTsLypAxTP6UvTiveVwG5cWHY829o5SH
C3LmoOMXFYZdIL5gY+WgPLjcjwVrl7M7A4X1q6XPH9lBXo0yyS3c4bBU74zjMJnfhSQHQ0whcO/6
LEub/g/MwG9NTA4lz4VnwWaDABSccXchhksEMyA/qmfXMxiHEe8mvBAxjh3WUpuE1yztcIMMm4xN
YtJdTNjJWXJj1szknXY5VPc42Rtsyt/ssYhSnvjll9YgAXx5/Mbrmnkep9qVOhF20d8BjPedUfrQ
tx82qvt1QVKqkYtQSqLt1F8k4FMDjx3SaizcJeB1LXkKI4KdOJY+SKEnRthA25ucbgB73JMK0mNc
tBWX5pSQj315SX1htDYPn+INu3yo7f25BWM8+i3PJ4rzjH+FuxC75crHMQ3BG4WREeKD9t52ni2x
Eah/Wn2QcHCQEf+gv+zlRKi1SaQW846/R7cqno/Tbf3Z+QCMRm7o3wIOo9wPCN/ROYXAdfqgRrsK
GFsPlPcpJiSMVHi2EmVRsOQiXx7PyClssjl1ClM8+SDV+Lf6bER/C309rID7XFg895gymnoabwnr
9Sfhy+f3jpEfwW2E/9lphbhLbMvIEFiSyLQMUrvr4Tt8DNB5J7nKtYMt4KZCJHC+6gzJ4DwTOJG6
nXudrAPzbw4IkBactFCcnDQpBn4HqTo+stCASD0H0o9EjHsaF+s7QVUkI3CdxkYFJv6QeK9b2W3m
AHXNWKtBFxvTlMGvnYHHvdpMFUxRrfOMQZKs61NG6FjI37S6NL8FUSz+iIPGnmIMVNK7mvW9Cufo
HeRuHRuwguZRmRq/MW9uAa3b4nY38gF9HdL4/t7SBwTFoPUj/SjXx+UVtkm9giXrAB8aTmfkGBVS
JILNjeSdtAvKYo5zlbGctZyvbfh1yrEr3TyHoXBa7Txs/bU4xiIqGMiAsARTNNyC6AY7zbh3nM+C
XSolVdv0XjzCnKMXiF4qlUuHOCHG0R8jAGciNrcUnYswMK0aQjjtZJ7yEBlR3jJiWoC4pKPDOPJM
A2ef/SHGt5BlTTJ0PJE3C4c3uxbUBVcsLnS8FVA8tByuBFZeepcLYhjJ+xtbB7zi2n0zrDUBykqy
0oh39YZK4PVsbLo+5kGEGNSMqjyic5dCMdI3id2QA2676WTXVs4jgBIzDgyPasAp+qL+b+w73JVp
JbGU+7pHQu8GnvqShg1UVdVT6TNR56acTWcWWEJsH2HHKu1EN4vDDOGkLw+/s3iIdwF6DNn+yXDc
mAS8awbKWjMplxXNxE5G5sWgZZpD/vGluHCD3EY8BnlDbzLhnkEtxudZvna/vW3HvWJ1dcdzt20p
XH0yPaO+hn6KqFeHRZ0p/BWqi3F3KfEtZrnlagYb+oLWhbEJjZ4qJrDDNxMNziNtZBZDwNQWPQDz
9wIzFZdnBAASruGPp6nINEFzOWbpBkrQCHlewwsuu0+B5taPvqKerAPPIL1ss/39Fo15eYonQ5cD
hTCpdR5vRHXqeP8klEaWSNd+0Oi/AJJ8Hnh4Q3mBu1CRoxcG/VHEwzR+rO+sNBx/dULHEFvGjrj4
Ywe7Zawjj9522s/Z6iSaykm7KpX0RD80ggPSblw35TjXHoVKRb2D0XZNJ/JLHdzKHATGr4ZaVGuu
yFzSXPDrQbJrm+TImYny82gpXvvLN4HrUOP8fDjeI7KzGXM9dklh2nMcUdH1M2tJzQvI9/kRLPSW
KfiyaWNMaLZdr3u0Qw+j5/QP3CQArw9zTia7+2m3tBky7dbavub6g3oWb1dDL+E0zcdfu9z3yDPq
v3f4BHPvxxzLGvwQU6Sm+fbXJebxWz7BT8MJy/BliMWP6A+QSecODeShgkOQdpcng06CxqVqF42P
ZkLHDcYigXeNjSGHbeuNaQopha9fgqpBoiJ9vhvUOIeaRvlhj9ayvT4dYl4p5RcnZhFCwfdM02iV
jyItHBm4uz0p3Nh9zKx/N8NDssIRheOJ51GjIpw5lFw3TMna+scHqscc5s62EM/kPMLW3vARhjRh
3FI2WPEwX5iUWB6daBuEv5/2yEGnhW3eejdV7yEmV0Maheynz0uPoQ8SoNtWuzRBFNFIBA64pRXb
9MW8fGoyLNpTTMyXPupMi/7pWtDBcdqoLiMqkyuA2GHybhO2h90/8PTLcuemtgXDTew0q8a42Uul
rn7vPIfDmHiPlnPSWT32yY5EJIC33vLp9wQJt+NrXaXCm0zP+MmdMx4qZQ53pdlFG8Vfwu88Ukqh
1xZqBMW8lD3QC9RE4IWADxLbIT08d9xNUaDkmajWUHeuRRkqoKpBV19/dO7pgoGReJebQMGmZUya
O/Ei6byHGGt1UuJqBut5E2yoqpsAU13v5ueVk7XP9KB/kuToJDOpOYjeVQ0psw48tTPQGrUx+vKO
aBJKg4oCzt0zWNm5EQlgUn6QtJwhAGAtmvvNgNjRUkslD4pL8kXSe4oYGAAayUB9V1pS0hqHJ/mJ
9CpUuh9ufOYgdTxnZIDtSpPtPE3B+9j4/rsoSxc0KyisfimAP+kUlqjwLnhOZ5R/rXDtqp7lUKui
UXJu+hhGMtdL6jlHabrEladsL9GRgAp7/tpxPTVCoMoMXUxp2zccFFYiqOc8vS//sD5AUARkyPVV
V8neYQvuGjYgsKMzqcbElv1g3f0gDW+6x35N4CX/AGmTFgaGYT0EIxyYFmVuBqBDSPmsUULHbAk6
nwzEMMMgfJcUgAG+7Ythzg+KeLL/9pX4SbgkrEzsGyLEuAwNRzohgG/Q8vQmHHsZXg5CgblrTiCq
RFles45XRv+vcKRgUMi0Yj67K3t4Sd90kZzO20Em5aRJqG73rpcApz6IvUzUM8DOWBKJFi++O0TV
y3AzayWdDptGFQaR6JoQblqeYjdkfnijlhB/utGpBgkVFhuUOqBjQg2TcDnFdsyWD03lZX+6GSBt
unAwGFBSCj4kFxXt2D/Xp3cHgNmT8DFw7AVD4XoWGg5zpqrO/j4fHAGTYXT3v8pPZ9RnaOJx97bz
dhaRLJ/vtBr6m0bT15LMlPKzVPYaZtKG5MdbnaYJJritsIYhJghseDELfMlI+msAHhY/BEGXOZ7T
XGok0RjhqtwBTSRKLveCAg/FlW/Kyta1bnKSenD+VtkXveeI1LTnhZYk1JqQ3YA+Y7uUwImZvorA
LcVBf/ZuAFIMgrHVBMwhD1ourbhlpBA6PRDoLoqTDIe0feJGi3FnkpKaaAAd4YaYIPoJA1QzwSd7
xsjUKqao6JZf6PhY76R4M0cP3cEUvU7joqyHWLLDdAsO2MN0EP/9JzdN5k+Rf8JwiaAgdAFVynKn
h3T+9VwnVl6egpX7Tk0hp//aOwy2rq2ghuIGDxOEAurH5cdoXYrbuT2jvnUb8fxfjh+BSwA0wvdG
BNuDBbY6MijDf2JS2InhdcxPFpR2qZnS4731UQ/2JPPdjK8dRIgsU7anDXykgsLwbZ0jaoiDAvDh
J1s67Vd04nazVWgzHbj1IdbCQgfPcgre1tpJCnqwiUUY5ooDMFer66oxzhpuzVHCxfv4J0o/TBwJ
xYvyUVS6WljWnisKGlqfvXrgpkoapHrCR5VN7veF8Ee/WB+Kw9ILX5rjjWbIBhZiRHYQx1BAH1j1
0WRw0m/16lOhoTId1EPsyx1/Shz9PbGDOn6PD/qwOhZIPXXjZrSnlZfwnwl1m066yw+MG5v+7/HI
cCoif3HyV3J345KkAKm7cdscHKumwyaAcbCoEmk9eyfEGcTTvNoi9C3htDuoH9b2NnslOpJngm5U
JbYw8CjnSOSaXS+rbwJg5lMExLXjUiiUwu+o0wxau1puk/qieREKUHM2JQ20edI6efUODQdRbsgj
gt6zEareMtsDGU+CCtPOTqYm7I4Py7AUEPP1HvIcw0FK5SmX9MsimT9dyMPYxh+gKG9WJJj0ACjk
2Jo1Gd16zxrPkaZL9rUEGPk00rX5oODGUQpGg+Qib5G2vbHNi7ENSnLlXi7+dH0NXLb2t3iXNsaP
5bQjXMqQ9jPxwPAvKiUOWC86UHAgwMMEUDiPDm1KZ6lPPJbU0XK83m9lBEIn6M80Rq5srYDqilvI
CqMMehCufh/kpnNS5XOotDxpmpAg7AAzh6QD6H+s5uLEQeq3SdQhH9xfA71Fs5T3jBx+NLdgABdH
QmieHYELKmxyBe4SssrnzYbPodlD1k0b6467ic8BSCNdwtSmfVhZAhpDQBv14IpnhT1yW5DSfLca
uDh9LoaGdoWKV5wpQSv4M9kXtE/ZwMJaTo35OIEBZ/uyv4/mCPj5QsGlKHGE1C+QeJEDPD555p+b
IeWMfJ0B3/83IBForS1/coOtDOuBcjvN6I7fBPPMzu3NRBNUgP/v3WAGBqt5jCGXgWuq7vMJPS5i
vZIQY2K6jVECPBSf/4EK4BSdbCjyfHIbSRfDrJiQrrAEFzuGMfMxlvolQQWlxUKvNVaNbsDfxJMj
sk+Vk+yl2dcOOvAM/Bv6UYBBAS1TsFoxJU4rl7oqOr6yu0vLnDx0UFNOK1V97nBdSL31XfKh1X8p
Qxp5S5c6LG5D7uKy1hT3AFOL2KTv3y4iHUWsodm3bDe2VHB9NYPJOmfv8mpVY+F27+FX9mK2rAzi
Adb0O1mHKBIquWwvG00LKyzqCWxQSPqWiBUfty4usy09v7L9Nw9tqF5FUNy1IrjrhRxiqWDAAt6O
PBATRdbbNvlkwLY3qbwpN6BYJxA/m1SCYH2tC7igVhDZc8OC6esupKYpN3U0oGkus0sQxXV+mY9I
sxKpNonzGYqx7IU3wk35V/IjgFMnNgo1ZrtELap4qcqlD8c23MvIGsuPxk3pUPlWPFdJ9MsTFvIL
AtMmAakeT6fTO/OqnMz1P/ovrnltSJAEl9RkAwFeuWpAFPGenQWR26alFgsDFRFllVsGfRcc2IBe
MZ98cwhAUK0r31YEDPBb3gzKg6GCFcLaOWLiiZPIswGh6oEmzK0BwT92GAcd7E4p2hO/6+9MMSuF
iyA/a3uvBm9DktYu0KIeAQjK+wb1BJ4oNwbVQI1Czb9apUS4GLMb1qQO+1eeHQ6Era+TUmHpt0QL
yQ2fEob0QbMwxG3tv9NWGH1kliOVzJrg3DWzImsAh/Q3SngkxZvJEVGFKAlR9zMLeqItak9XMYfr
BPiovnGVaedhDDpe2VdPpy6nNkn2yHw48Omw2f/FYCV7aVF/5mWi1ALwKHR57a9xeSodynCu1TrR
bEiLSwOx4jXP1JMg/RVy/ROXViQufrcqKKdCrIuFqRHoKVkWfJrBPY+rEdIR1U/bQSBigP6lFVM6
3telm/QWyK8S+NG/6Bo/N+bsLCuJVCRLd8xPRoUCk1tO7qyqXT4sO77xlx4kePmj8pvbCp/v9uIH
HpbNg3a1kyHap5V/uEfdCzW0ZoQHxDBMOThs/bdaQpxRtk0x+fS9XjMMyUAIkgikiWP8f9VcaPkz
qob3lPiGeIVHvpi9/lZrtfXOr8Fb55B1UHGub47WclCSvNcYX6Zs2Ep9sk62ORZfLgMVNKyfQdMJ
zDqRPE73/TObVNbeCT3RNqrf/YV0thDfrK99t394O443A8ZfHAUqLYhcaFI6IWuxhOUuQDkM1Z0e
CPHc42tTAnSAx0S84wTbDj9JJggeQX+dbdvvzeEh+J1HexzXRheWFlyoCINp0UHruAhO3Mpu/B8K
WTnYgeOKrLPJu2EJRtEttQOzGEAM+m9pgoRUpxmFqfFSr/iGU30y7kr/CCiGToXE+oNik1AleZNg
pv4yGMDXm8KnR29vhzUgZGikvhS1v7U/CZRtWEBlfz+0Km5w3Z8FiuDxqgMp2CX6XH5G2B5JvyIa
GZWFNmOC2dA21WT7K4O1HeRKq1soHwsgswmmL9Fc2kQiz/9x05X/cZZos9STsowGt7aCQxgoPvJi
hm9mZzaUTwawy+QnBiSZ90USik+dtkAuwGYMZpc3Bh5cSRcg5Oc4CVgTcCiaviZdSELyFTFUAhHY
kBCI2Cv81hAcPIsXVS/hO0a1+zY2/l2BgHHGchg28swllt4Oh5Z7qwPqUBADlccpd0aOn8220TKb
R23YlHQCRUB5c/KFfPeFRzu2nqlkUXa62w95/q+vzCIItwHDuuDUjY0tVdBn4CNcDQjSzIpNyx5z
nJRqEGwqalcyuw2Zl9qKcXD3IAHQYF9Z8JYUSNnTQUVKTJI7aBlXiIYXMk+wLJBbzLnMpqs5hiqk
mr85qpu/NWsjr5Ytrt20UuHThk03wN4ggaEhEi8UHsyCTqRBVRJ2Bb6lMND8enYT7JTPVqMoYa3t
yL6N/ZWT7rewmgDzssz1G8gcDBs1ixqdab9s8enCgznvx7bnI/w6wwMV5WFIOklvijXgObdJ39ae
YuDJxVW8M3XJnm2Bh5xbd+/7OTsMFlddnd9w9F8x3hDAd0JFmnqaYRLf3CPk0vsLCN8fnkrEK6VK
++FliNnrZRqWtIo2yoZuvcteLtEd8OEu0Ydkq0womq7xad3Y1myalKq2+9OupgDg/UWMGjwAQ3CV
K3tIcsKfY3OgPDXJDjAym5vk4eihrE9E8Yj3+ydXs8nxJcW/E51AHdvu/TNcIhMwdtlGW3EoMFYs
qvy5qvWb/0eduXykim510wOwgZ+whCMT1hI7cZDiW9O2c6RXUCZdnT8kmhkB8BqJRI+86Z5esGOH
tICu5zJCWDDsAkkGM3ip7t5Jkv4KaVMAYw20yPsrfdmbRt47+GQOu6gKRrZmVNLoSrRdBOG5qhjA
CQosVMClceXto8Rn9sc1Eo1hZtYE/3tA6+UvJrjxNWQ7adL/AH7EMLZJ9gmEblCa/+KKc1I0ZrT5
D5fC4Oc2OTNk2rS/KcieA0OhtHhz9eUK77DwwliPu6hZRqDdLca//6vG3GcwmNAO9E5Pojy4vx0p
2VH1wuFGgJzYyE6sj8gUgGPTpnqW4ec7Q2JymAOeEHROrxvr65GlP4kFYjll+pgbfPepKDDgMPRj
2fgIRc3O5j9GMeNiBGUhABIfARa3QUNTBqss1zsEPetxj4/O3ynC2em1Tjki16Zswa58FsRwADlQ
ta0WzLL3cC2eHSBQy/OvWvofPFURA92kXFygDatjJ3eu/cbg8GrxFG2m8gzVrFMzFKzdiyE2UyIE
kL3TimQ48xoeoWxEvb1paTyrhgsQH4H3D9kz1mL5hCktTcvywVdNzGtjQbeVpKx4VKhyY+VhaxXm
a8hHp8JyzrD9U0RgVrbOh2jTzyxIojy+jsitU+x+CqOjLopyOR5w5++56VIJ7Fev2KNpRA9yJarz
SZ/nGnEuBrSxU4iBluK0VhQhxc2NX0ZkNXgiXmz0bfnN0ul/qAejcjzmR+G53SsnEx/OW0WiaSrC
SNsK8GknkcqeaEyemCPNUDwZd37xrnwpqFb5paNqyNLz4WBr3ecjkGAmjLWFEeyO+kBM/Y6SRdUr
s8c8nCHwGA3Mk+zjgDgaOSHz68NDKazXGToz8CTgLAkyBh5MYl4jw+/WXlY20J3Nj011k8/lhS/3
3MmOx7x0zQ90rNZwc4MO6Iinnu9GD+DSAGc/tnwx289a4x2AfHL/VirhPqR3QrGLipNbvdmX0yXS
p44BkI2ySIiIqn5QqGWgDNcxtpaWRVxXrF639bpu2J9qTUFo6+19B+sAnq1ejLu+VHQONkHGXT1k
jQ+FJ0XvmB4jsNMOJDfgGiD4upVtqz2QxjtAJcsayaZYBALzOACUmG6VorTwOESJS2ONg5E34hf/
KLVeXzXOHR3VQlfojHr3NMwWZzuFQoBlZ7OHL2BfsST1UGat79a/UKmBrP2xK/bbIca6gIaIMJoU
f2PU0zcOxvD6YBrvA8+cPuTZT7JyBH9LM9DoGvznlDLJAAgpdZIR3PHsrBAL/5/HHLZS1qjw2ByJ
3k0LT1f4vTRtrjwAnq2CBVEwEmkgNMkeGUunmORHanLpVls6qf2QHJCh9Jtrk/rGs5TS0tBTZ0+B
IxZ35ExuaCvhI0+8OnQxM7ydETq0OrKZkQEIlpgje5IjM+MwLMvzk0GAQ7R5138rmTDC7sASbpIH
B0EOjnkhtjNgjpmHuny89jWrLGkPZyDU9fgCVrOd8hpJev1BJVZVUUun9gi1sykKDE6SKbO4iYXA
DSjbunzx7pQBio/NHMQ2vp/v957POIWmMR514pAIHA62YtBInLsCwMM2bYlMg26lIvAstb7FMfFJ
DTHJP7BvmvRGqaHm2TznXJ6zxuZxr9TB7Ey/vSm/cNT0Fd42GeRj2nZ30ABTTgLnAe4YgKnr5Kll
KA5M04y8sSQtCzNZTJ1FO6XZQPF3/+rN5JQ9jPUB8GYxKYleH6q32cINIxvBsr/i4+8FX+h+FH70
Dd1NqFJWE4SZcYjzpkCAy7outxLjmlLK/mdtLuPxM7XMb/gIad/OFZmVOb/K525+Sr02RV1EXROK
Wj7tTTY+QlAyWTVK9fB8YoetALi3bmq6y4zNT20pwAFM/IgrrAAsdgLHU6yGWMeO0xA1eVZeVkrA
80FT5LXR/8moqN/898b+df7z84ZdIue/qmzKL64/eugh8QB2YLdRk7vvH0IwIuSXLgPHWEOuas5/
YqfDZX+fC1TsWAAtbm6wjjtl4qvuuS1D0lnf5MJUMXdDo7OZZ7z9GStGlmUYHCETFzWDdFmaQH/8
X8yS6LQKaE0X9VT5ygKAaj0xWayo6ijEjlOXgQIgTXJARRrlJPyvRBd9kHQ8zlC4Ux21iVqSR5qL
C6qL75C2iVo/iVGsM0GzGurKHrmMJH+0JzcP0nMdxSR3ur5/nWsapUWZ+mr17PmYJUTRvsQjIdNk
eIlPuwaWBGIqu+uE1LrVfZEDqVVKDH6U6Jfy+Fm3Uyi/FupEcnOTSFgMlWpQzodhygOfCONSB4qX
pW5y938Vf2y+811tUoi1T++owT63O09Ab7cgHXghTtZC6Xmq8Shm5k8FXDLgKpwmG6s/hnh4Dq50
2CBFKmH0DJhdw94lLIwKJwwJA/nluCOCWljHSutnmrED4XAOFMY0mJpti1rVjaCeEf7ytlg+bbWN
eE9sZqt/BBNU3IR/geaRFxTj3zUhBlQ+Pu0qSCUYqNsErLGJHV1nTJyFzZP+omX8xgQRS2O2j7Up
ZEuQSmVAtfzIuQ8cW2ngAn9OX0CKh5kIE3kfkPvTYMNeh1tIVWPuSBHQQZYy1Z/h135TCjMCwuBc
AR/JFIzNy68MWk7nerWRcitMzDlMaK9EgkEGabKYd1Mo6rfI6uAkPA76IkfQrq3G2Bc49g3t7Dxr
Z3GVr5gNOZL2pdJszEIUuP08hf92RV8ZVKN+9paiP1gY7JBmy0uRHkop3HZN4t1TIOrai3Ew9GTT
dmmzdLEIwS7frbwVC/GhcYqZ6RCDAG2knvhtRXNDT10974poBU8dPOlT4GLuEKyI6fNTEBTp+ptE
pPsKTimKYHfMNg0CzxhJnxzuj/qKrLHnxX9WOcLcPumPYoe97lycfGs66CMqgM8Gbw5iwosneZ2E
aBhThoBClc6EPM76pig4UoIcLBaezaTSLQvgJItR1/hEIy6T0xR2yheUxXLcsWmaN3jyuZaWfORC
JVoMz0bpanKgW2qhhvtRbTLGaMgdl6h0CJjBmKRHXr40mYx2y9CHPPZAi1xKjjG/sDvdhrv7AVGc
hkqpxDM0OgwYWPV3sdyMKF7WlrGItX+c8zB583cT1A7+gR2zcSQe2tYOX3i4E9FAm+10fsQN/uxg
sZjolzsLnO8h257kOv379/VWsSrgzkt5yfebQXB3aNQNkuu92cewfK0yK7MhAo+wMPEt+evE0fbq
uAi7aaH8bwPrCgIe1zoWwz0degl1hf+etx+Js5Q1t3Vx0Frvd1BH349Us7vduprBMHBA1nSm2FJr
EqTmsP3hSgLvHR2N8+Rad3uG1kOO0a65LRVX8TWGk2n4s/XrGwZ5OCi/2aWVSt8io9d7NWMmKvKX
t6m/zK0+k4j5Qsm5vj0b2mEYt6nubnvpgHs9a5dXHtUEk7Oxp51+DRtgTPnPU4DlLkkzma6B2c2c
Dw3H54RUGgQ4Scr4YwIkDadDcgOEM0Gc8+grTWzmgkPzOmr/ngQubdgBzvLmrUQpZ8MJEjFq1CCI
Cp5UApWxKK+1tFyv0SSeDCzMIeG+xNBRYTFJWKYLCjUsDmARgfUb1QQN54wSwZ3g0tTxxEULVakM
TIsInnZwdCUI7HXKmd8epan55a1qeKiYyyYi7QD/KQI4ratA6fOwgtm7C1JBBIJtuskMMsSeBLpJ
yBjK2YdrmNxDY8ER5/gsTbwdZahTTQjWsq8DjF/my3V5vAJnzDSqScTE/8reo2x8YOGoIQbsBulM
PdYgiTCAcnkcZTAoWgejFKKQLOZDlOaz5z2de5keiMwb8rRu48Ql/h33HjXh7cDHKpbeoZWdiuhO
gTsO5hy3sY5EYgsPWbUWmrtEgFXq+mb7/HyM1pcXfVG+NAYyz+5SaniHbHenWU/aqAy64aQtd+vh
Ksh0yC16UaAZB3gOAqjSJoNEG5/Swb29AvWfg9GFEU4z+Sd/JXPHGRRJPlHQPjbuK776Jl4LNQzm
C/NHMXsw4NPIAG2tPkCzljrZ3HkEPTyz+P3OIOuU0HlLLXgZXeoh4Hf9/qHfxR98p+I+JQMBrxwA
mqFLqer4XxutRDIsV1O+s2X0lfa0WU4AQ5itXfkdIICDLiiGVcRomBlPFSeUIouyKgccRKMLgL07
jblQBsp6wFZ3o1G+aq7wfT9FU63pzyB2EevfAwx2If56d8o4e6X9c+ZFhU+eX6MDlEdgy6ECfZ9h
ezQh+UJx55NrwIVMYrA43myC/PKnazED3sb12i2YxZPJ5HYWmUZHC6kaDiASRPCQxUiSR1fqspDP
datGZxA4bR/8wXGJ9+sp3PLDpfID/kSEcOqrIHOov4M4saRF/BC9kHOXALTrrhsX3k/fYiRKDpqG
XDJp7IRxHXL/lKxhAeX742dR4blG6hXIN6yiG97hIg6IH0HOByTMVxwRpVGSEC28ZIbhNCCRW2/E
NGV2WoZEoLziGoGoeBRNiPsl5nT1GHHgEHX8QwGclpc1qMiMGgBNhuNm2ejd/rDYwZHaTRlcDKpU
Q/1YTxeZh7wF10oYSOwAC9ZBTDVQYG1fHCyNDP/lLpF2YF9+kxWxf0YpS65gSIpAr2PdfxFrQLuO
CEq7GAGYeYPaKmHYpQAwPLAt0sH01WWHoQNR20o/eeW9b10Y3tDPZzlgBJlu+G/Z8PjjES1jRhQO
Ltfl4GCMg6+h2QSfGE2xKkqfP5K3jaVOBZ390oikLbgz/2lwU+T00bJSJ16hKzLH8uEtvt2Pxzz8
jKKJuWiBVQ9+Ypzt9umVHJiJrp64bVHfyFpo7+JTT6YsUSYG4jIY7MyjXb0PUz2z9QipxeAkkTXt
BEaGPt7lWQdAdPWls/9v4OrZ9wjFF2krbo2IzQjChqGIrRyybvCNfrxQX++0v8fOI4ciCgnPCZWB
tINZf6TnbQV8hEjf9Kew6Vi97VdbOhvSRjRHlpHId48/eL7g2wGxp+SkgS9XDd/hCOOZsbL41wLJ
JpOr/yquEVkVHQh8UkXBGh3XcNmrRZ54Pt0qv73aFPbecqwitSRqIXrvOTR8fCZGgoYLx90YWMaV
ZGkEAIUPheKIWwGXopRhM56Kr3NjE6dFlp+7MWLrvw19GvJwwnkn2JX17jaFrvImA/TmX0y3SCor
m7vZnmQBMepgAAIV83Q2Z2aCm4i7va5URByqW+Jsj5oAbPVWiqIBz46U1Id+wakEpVF41O4InkkE
R2F2qmUMqlcwEJPp7jJd8Uye5l4HgindKFauwF6Epaai8ROsb4CInB2cgbxONflJKunvtcGlpu9s
wgAmP7xoER3capas1CoyRM30+zwnAzS7YFz2G9lCrUAubrAibmjjHyxeYC2gN8tIbFoAEkOI+gmK
tbN18ywEzhTmDGJT88h31IBHUGY9Z2hRlFdCSjy8JgSlCDm3oiiWH5n2pmLPySuGx3fAVYuHpGjh
qsqBkvXenAMnrRr/FmJfx15eQriT3dFp/Eo58XyCFQSne+1huQC3Um5kRoX46FSOOnm31+YY+VkT
UKL3IUQK19V2J9aZB1FNLyQnRo6FRtCRDXdsEbL6UrDhL1gSYdyGQ11or4BfYQyFHxFstmTaByrV
OW/0TZhMk7Sec/x33N0FuEOfp+RBjO/SVQ12agKKbAQXVrQdUTGexyNvle5mqbpAsboCcWrc6Bgz
tDTEPrLeazLbF+BCWDA+YAJdpufo/+kCHdvVohdC4A9wwtAI3GjD77UNxz+6p2mAKXkpRLUAXNAs
Vj0YyPifMDMmtU0+cEXicOHjTGIFcQu/sk8vF79fKVDSAGdMlydvNwoX5BWhBo+M2ADc6Od/c1Kc
YLDDEyzdvcsslAYn1WiXo+cTJiRqbY37+sqUZs8I5aomrChWW7BQSke5exX9rkH+2S1j5ZA7SKp+
2XQLaZnZZrGUaiycCNX5q+2P0e6Z0R8nJCoy7F8rUsSY250lBAdNZfaBnaN8wDh5XbIbqL8A8eBE
yutMslbmtNdm8EFF4VEOtY0lsOqtyJgofTAJvUhCmrjPLc6DAEu+qfnlDa+VzpENRCY6wtdEcs6c
366vKWUB5FJW0Z1U8Yji0Z6DzTd49MjZXoMDtE2V+HpZArf5y1mrdclIGRONh2+Ab70aiyxyXwmZ
meRlcfyUVCN6r7pVXnztSSCAOM5OmBOuGqZNSwA4VC4Di/NLGCAlUSTFxFb4RsF8W3yMiXSvYwEA
ns17rHvVCsHoUo/EyauRQ2bOE9023as/B3TlFxwG4bpgZXT36RGn3X77tvHQ3x3WAsuJ/elb7lsa
RnZhyuTun0/o9ZruWL7z2KGyLbSdm630i4VM+Ltz1Nl4Y7GMs/6IGVK4BCgvz8gm4kKq/eZkxTey
7cahX+9EoKtYIJKUFOapJMmFy1BNcfRPqkw4JSLPnHmIev6OS46QQRw1Gol07wWCaeWtP2vOlg7d
haZiM5HFJVGu5033OUN8wu3SppLoAjqnQWLJ6NVKm1BeO/Cpyy3iymUe/h2rDlMnCya7w/pxK1Iy
35R1YZgRfFrvg5/lod/UJAbxrcv+/xcQmox2D9HUjjLutDnpw1O/jtCQGmw/vjBaoDPvECyAt6RW
mw/qqEX4X1rdBVpW2165bb8vwaT25LktarSwbp8Rb8NT8UPfs5aFDLBZruVn4eN4OSjGVfV5rL0u
+v/xOR6iS0H9WZmEf6FQRniZRWRiLGOupVGG8w6eQJ4HW3Aq+yBhzpxlKDZsAPdZ/LYDOCRtJi2p
eB7LYgxCs87Nw93E55OMGuAd1RWSuBKFsIRkSRN03fNQ7oBi2xx1u9Rd0Pj3P6HplR/9W3VwujYS
KBZK6LxuGdLgnyamWyzZrOl2Y9jU3GbVrq68jH7F/xlNIbvb3A5E/sEHTLaX/Yv4kHSe7K20fVLt
XOKwzLxbJEL3QVal3dVSQC8Gl4O7ty2eNZAUiK0xAudUCFRKTWsd4bz2bfTIu7saBAgMurwoopI1
2NUu+yvnxSVwdYTeWy78myopSOMYC/3MK3iUK8po+BfgU9dPBe17G1PMEGCXoIvtEnOhQP49Q4cY
sEzacE0uu/YiLo/JnztGsjcdjMFyCRyC7vfM9CEN9CYgvUeFxrqo+RWYnvLh4Ec8kgGSyO1PRIMJ
sclCcFtxmfgIHJoOyMRu7v8AEOfI+B8OtvSj9MoU8gC1zDW9F7LAx+PLKlxl512UJ+/EY/sHLts9
udBdpiqS9tX8EKsj0mkvXZsJU02s4fDKFqHyn2E5B4zRyjY5khWaGC+vJ6/TVZMbEoYyrJZM1tBA
IpPrRmWwMudVEr5G2+5X8ObWikY6xDkxKX5XU2zyxL4U8aCl7vraC6XU/MG1hJjwm1Tr+5bxhyTv
I36kopKfvBJnuXDjtHww6fPnoNvYmQ/szxorTQPe/flR/UQDOu9Bk+34LRBQG7gAzS76FYkxqP6v
4uqvXQ8nf3rLDG1eNzkfmhXh1siVRly03ipBdqXXTI1KsWwQP375SxIBnSAFoDazuW5MRu+NKL5E
MGOGaIGmyPOnJA693UJ4bhU/wPulKE/wzWD0mamCGVbmGPcDiHp1KCViVYY1oGZFA+FPYE+sIWkn
lopqFrpwHvZQQB8BukxgEpGysuQVlYCOfjk+DICUuI4R9NLQFaRw3gnbiy8kkonMeuogp11UM73F
Vy1sNEcAxMRSGcCf2WkChbsju1dSfvIg1984wU5znkpGr+g1MTS7RdUC00hxsbPPSU/Y6vrdSFGk
SNtMFOeZT9Uyp2BXwgFJfpJd7rI4n055O1Tz5K665UMIjc9/vBoea+YvoOkpBYx11tcoJRGk2+4o
amrVirapyKy5gvDSjG2wdxUJGkFH/1HYtPlfHia5y0RTBBaG+Z0Tm14wwwCqv+wPK8qimnHKKJQW
FR2VrMcPjEB3xj8bJkAy6zaEQ+e8kS9rcIMs+r4ewzmM1ZVYBxcoaqdzkp+NXahAwLZeSbDXs/mA
fckD6AaVQ7aLFo21TuKuV5Ci1HYq2cCs6iL+OA/E2tBo0qXOqHqsy8OgjLC6PyywrSM/84gEmIZz
jho0o6n9BEMq6Rb0z4LtufSdd0BxxIZGG3hjO080TSXl73PbXwGflXyuEdqT8PYBBbn/z+zck7fR
7IZmdRVjAyZ/RTgCsQYo/F/mvXvevWyLGaBGUXWFl/n7ZOPreHwPVBGOPprlxy0fnt7mo5Z3wjZ+
3VV+FT55/Ktwn39rWpjDW+wH7lbzqsq3eaOY4rDEBL15M4P3nW+4APA3i0kG7al3wM0eGSAlX/fA
kZm7W20nGjLWiwBDwb12IEGYwdeY9lrG5K1tRLN8eZzi10UdmdclGBzW33Ld+HMTNSBphN9eX9Y2
lpyVLs+s3sd46oCYevGCaonen7kTXvmoydTih2UivTKP4Q9rQ+Ovi5X+yZfaS+zokPSIHJPdq+Fl
xQYtA5cCui0+kGgeIkHQ7IZqXIq+ftj4NoYC/yUqrAKvWPoonTkim7lHTMO3+gXFLMPWVgVruX74
2jthqqSX98FHO6hVmRwqY7D409kKnws62hR0BE/vsWp0VIIpVGl9kkuS/c+fRex3EG10zuDwZizF
4rTdMgCHZ4B1awHmwYD8kgnCYFbbZNJA29VFFMSSKhCr2S5mbkl8hE5k8DhaIfPQx90ouiHQIuX7
NI3ONW+pS6/o61EGv3PQhJ5oC18Vv3Xg20cf1GOg2r0Lqd95Ero9TtDYCCEr7ObBqDeEG5bAL6mm
FTOiINbFf/Wokr3s3E0rQBDd84z0ASZlG/+6pQvzAnydh195TcA+h1lAUoapDI9ZUhtvjCs8eBfZ
gY3Pr16xe9k15Wej8cAgxJxDfgvYSrTlUu+lv6XKQ5yvQ3NIM9F8ke4uUzWfB6W7uyaiKU8vz+Nj
prKOiv7E9kg9MchQU8tRZVx7zxp9CWLkoeF0NEcpn0AJtplWWM+MDSqj0G6KptvByKUXGKkWdJ4N
rLEB1ZONZbNnWdzhHMQF7T/DjIKFsOIu3Gv56efmxFRtTdvizfNYy+Z4Qu+vHybK/G8CVdia6rMM
dd+K+hV9+J1SyNE4hEic9lDFcyyhZZw5eTk2VJiwoSweoJ3AUZs56Qt3x/08oIbRFpC6gxxi/b3t
PMjy6rYuYss/pPs7+UM1FLG6jVw2qYGY0tGEYCaIOe8JijiBLRGb7I3OJqvdu2lUJmYAGgbt2xuW
MPrlIPpdZLyLJuf2zgmmEiiMnnheRGw0ng89QbrDDC6Gnaay06OuXNb7P+k7gbAAueI+LJf1v94q
qydt/xIPMVGZRdWXNotnfUepq3axtOgnueorLA9wV8953b35OH1RpjIL2Ie58Bk9xnmFoGTrsZP5
xNn2DlxCYm2bFN5xv0eji2yyU5C6jDvC4eCBrL/CWyeA96uIn53Ztkd9t2vp9qLqAgATqFeHfEbA
YH312a/F6gbaoOjT4vR8b9t0MC5IE2ZmVgexMnO0jQUlKdMBvLKdvGA4zD+JynP73+yEC08iipgC
ZxUfEtj4XvhEM/lir7gyMHJ4pc3wz9f58HsM6tiG8uWcVqkejOn8XlO3RQ2Dt0+6jTZ8yzY/BZnV
KXqd084rWXQO2bUtxgL2GPKWpCRRf06Jw9pnBzwXxcWmk5YKkmfMW6OymZ2qTBs46JAsrxKH5zWl
FBqmurPNSvq77I9MGq6f3nyadOZwGAEA5wzVl4ZOIy9csKtYSnk4lV2v5yNJvB8orq6MVcPjYKx6
ypXg/XFST/ukxMlfVFbmGxHCSBto1csba3C/lf6K9FQOWmJXLc6antKqPiQWE54B3dBx1DzbyZBX
07eg0Dydy0TjShiqCAuM1cEOD3ZjzHwGcZjlybfKfxEMv8KTirI2l4NoYOOmQ1I9cseay7ItGsRB
8V9lT2pWgmUr1FkM09IeGjPsQaGQIwRCuHAsZ4lJGDfvpnwUHb0OvA3+0r91sa+ZfjWFRJuJr44X
J8tHFs3HNiE/PM80AJmczXxypkN692lpFEnVAS6Kfs6UicZNacg83ib9vfoEI47oTfb4tPkwQ3Ii
maqXadNc4NNu07WVyJ/kiCku1kVKABAbVKbDCeXx+F4Djb6OEo2tWyB9lrpa4Y+FVC2xuMhuO7+o
d5cnCOWwFyPEsSRld/Y6fJ5YdpWfPkTbKFLfnol/1uVw4b4unEU55ii+UUgZuBXRdtL+RJqXJkEN
JxMAGYL6kwTr+sg96+QNUqnkiaI6j05mND3zKTOu9HH9w2Mr+1QlFcqIy1nWU7Or5sK5Jxtu7ApF
Oi4hTYpnfUQ50RFH+VA2pr+fYYilsMAiMXMGGmhlySynmzzW2lcqzVaZKzOa4/jrGBe55xvX+ipp
9EoXinmnTBbzwixGrdBs8D78llf8SvN0xQI8Obd6WDYn0rGiZH/PuQLDkL8myyfd2yXoW5N1szdV
+FGULq2QSJgp1lS4tJpHWb0xjRu7zCNWOiN4knERpiAHr0zcKDSLqu1N0BqoDC58F++XYfGS8/Dv
I+1genfxoj1RiL/Eruz2WwUGbAFCf05EZbuBAJxBzv/e9XUPnrvaiTvOYY8JSsHGGErIXQYItY7o
W+NIofH77e5fLgKcfUUCgknidqPVoQ9DtW5+6Gfn2FqIo0k/KL7yT/gi+FquQr0lxPnbtlrD73pQ
2sNuZK0VhtLOg7PN0xUg5p0b4qV0ilu9UJNKoadRXxO8YuuvmozE0p2Qsr3wJTrhAkiDVLZP6ASD
Z/j4i/a6Kfg5bWqy+A8gwHL7aT33OkVoqnmS1JFcCnj9XEM42wDvH5QMBasOie2K4tp6J7ReasCF
Y6NN9uqQG/o6B0TRCBvDWmOxIFw9UHn+ZpdILgcdLEwMTDOyPe3JYZ4V7AoHM2TPMm3whJL1riq1
+MZwsquz8dqjuNJCf9HtE014tcDH3ZA9u5aXU7aFl5R0Uzao5jqPyXogMXLZeMezObKAbktEEJX7
iScvWrqDwr+qOQzfJpjsqHEUi9NAhYdAeNrirG2jUbV+i0rEM4UufvEeAY2kcMFzK7AxsiykVgGE
kejS54YYwt8OtwoD/IEnBvGowDGu//CIreUo9Fnxe1qdVV9letQYus+gfDe1vW2G1AyWMtsgPZ2n
qG0fWOcSne0HAWuqBzpA7O0NaZyinsS/0qktJ82pkLGuAnsoenVS+s3JB+QWW2jpaVQKWo65adGB
BTkxNnKm5JeX0xsVARd9vG6XGZytb8hu0LMJOaB+IKZaLq4EvDaX2FCXeexXaER1DcpsuEd2d6kJ
DqNAmgjy/KnE5UNJWhd9mJg/1SlSvgZ0dtlSCmUZXACxu0ERj/NTYW1lO84gknlmqo7OuafEiWzk
Hn+xTswWtKj0k3ut6mDaGX5R2u+adotz8MNcIz9JEYQ5BJclwprx2luF1lBME4y3ftpu7Jzh0uQA
doFm7OnX7YhiFgB7/WEp30Z2RYzAoZtqJrP61e5dpfqY62h2BFCQEKZkewY0wv9n4aUFzpqBOnME
Jel+9m3vByu+903WSXioEIlofenpppJG/q5cUC4DO6jqL9FUTEeOLxlzloGe4vUoBHQbS40Y+Nlz
xiqji1gH97p1Yn+duR97byQNViSmjr1Gn7vM0rIjYWwox3JpcJ1LdEabWPWJpBaDRgLWhd6cVA4O
HOthn6c/zQMfxwpid+cNF8YX5aZjLafMTX0hnhbGTBXPrGyqXjXbmJU/6MlOjhio3t+0RAvrO7Dg
OEX9ridmTk8XnrRWNZk9RQ5H3AOlwjAQyilSKgNchDcBTA8LnZg+O708SGst+yplhKm8/g526L22
4QnG+t9rsXcFGMlgdtaZ07+HYcJGzi6pEIJxpPcy/XaGsk+Q94I5fb+ewWh/LM2k7exX3L590M2G
KtT8Zxy4qRoFEhKleuj1nSrNvP+QEpNJaC+NnBNDCtkmd/CH2gntr73cZyEK2k8GKcIgHibEFC+c
Qxabm81rd+0j1MJZZjAQRyUHv8NQRcPLzYuqb3jlgWVEisEF/6+NF5X0CKnVabA2Tv26U3goXUcU
B+stYFO+SkbkOhAd2urrmgF9Ru8Ege/24bSGHOFVqReJtFx8reMEqFCtxX9I7/RZZNmY6VWkRRtA
edhgIxyCz0Y2RDRBOud6GD5B/IsM5w7EMAiG1BwS6rYgaUjL3vdK9t05o4r3VO/I7VVdGCck/lRH
b23J7/D9krjqlHy2SvzYwDw6cac7y1QRoEOYVkG5h6FDm+aMbfbvS8Ad4hsxbVJ+iFz7/JHC7OWx
Gpm+J2kzbE+tLDXihWUCg35uyiFe9RYFxmBd62HCEPzSRO0M4462Mq3oUeiK5YTLXOZC2Bn4hnrx
vxWKf30Klx6SJ3vv3dTz4jpM5/gehbqqPv0vtxAN+7lasoGnoTy6SyQYEvT6tASmUUA+Tj6R9HAO
7Noz0Jn2TYEi/OqxKEmYZR9tJtTJWn7dGLLD2FiBJme9uHWvZGasdvdw6sF/mfP+AQ60+rhCP6br
EIyYp63goj9hld7MyGqYF5Z2UNCW3KlHGKzm0D3N0phnvaach7pa5iGt4s31LnapQzvLRwrFX7Ku
jZgIFocreG1L2lCCF/tgnAiRONxAoGtP66hXr7/7Up50++2pM2ETKrlOwcrhAILWWzmgmuknJuuZ
8DMWeyWyjLXYOQbc8+2Nd+WceoZ/zg6+GKJXVbGRAE/e9tPVsvsoiai7GIsxz9p22zxlC4HoBidP
DJqoVdOlNndrwfbNi7q17PSFRj+giYslLwdoKAO5jdWZS3wnWIp1tEfWsya+/WbwJbMsY+BS6oP+
fptVVo2sbMqDSezn9zIAG0lbrgGXBnYeNrh4H5aw3dp07n7yMhTSyTnSvAV8lXNZWEDR6xNVJlNB
BlQ0OoAELrnVv34eTvS99+dtAgpkEkPGfKiAPeK44F8AOb8smY/3NbPv7Yd5f0U/b0OaUWU7PuST
kyuFpd0ZCK6NhxQFXF2ibgJqNUrjvr5DdgIous5e9izJZYTEs5JDea9yTe9QPDQLCdR3SeheD1WZ
d3w4NTPsaftV24X7soz7uh3c06198HwqGAgFEcM+pdLF+kyOqqoelllFY3LOjRzrkTx2/Wb7/3K4
rpR6pvpqmBPCP7tyHGFpZ0QQVZcC7V53Sqr+qQmWm0Zbqt7z0DkViy8nRJveSMA73Cu+iB7EFGZl
fcuA/THZ6QwVFuVoG66F9HHOAzpfpBboMS14MzZuL/fSLARkowdUpb2Jsnjo6rcGDiiUsbLf+GVm
4/7pn8/8cTGU+CwFvPofg0TZwtf9O0k7i2PjmBa1JCsPkOQmfL7qISH9i+Ztm8H4u/WT8nbaG1Ho
kt9IPPfva1c3U+y18DUy39PCU8sjypYiHoBJIgXnI56EfD3ugCaGVmUgS8YBJqBPM0nGWsQpCmrh
oPGqq2phuSmBlt5LBMGH6WoAJy7KfSl8gVCGQ0dJKVehTE4KknO8Lfs97ANrQ5zmvAibeOwDgSjF
R/aNon/uCgoRKWarCIt6UjqhadLeHqUYEYytVpmeqeRFvKyHhco+VCmW1koygeNfPuvC9N8vHWk6
imgR8I+4ppbHK+o5UIuk3enfjdcZrP67Zu+SrMXbxmQnCb0kpDiMLd2VX5Nq7xf2095g8+Qa0FVZ
VsDXPTZnaX1m09dE8pNmMVwuQMfetUF+MfcAWGlIYow/+nMBIpbA2zJaoqF0kgi6St0dnUcLPJkZ
420CB04m58mROu56VuQP3eu6zpyckjfyKQk2zQ35AFJcoK5VLT3XshDkdufGIt6cBtYzcJyJAVXG
oXf/RIVxxmPM2G/M5Si/KYIfeyM2aj7x5R2ULzHR69mSR0blDQfO7NFwz7HI55fZt8sHNuVC5Xds
6yehkRTSfZtL0rrl1wNmkYj9rtQzSOhz1ROS0cH3t5t+jYh2v4iIYyUFNEJPQn95wKCpIIX/zcN/
t3r6jCD2hzLH9hxBV/zFZplQCkcBLECCzg2RUpS5XneUC6K2FTkLfFbTw8fFABfWZxinh28ov6nq
HG6h0+Jxg/+jqPcfTdpq03n1qPoM6ZzteAwrp6j+Brp5BRLrcH57I/q2Sv1/onACqzi/Lm4TEp1g
K3jOymA/y4f4CcvUaeizb1q7NI9Iozl420JMjlX/sXh0lEx7S3+7briuUtZI2hXKaY1JbCmTGI3I
0X51C12b5hc9Mf+bEGEpy0Ui9ABfwgCuVJzeQEPoUYrul2eXJkI/FnBuRupJYzl2fJCZbX/W/3sz
xJIs2j7WWzlsPiSORExjtKOxNdJXZto3ZjM4ko4Jy/6F60pVIzml+IqnlsSvl9N9/x2kfWLfaNTQ
aDJfFBOyw0n9LnKeR4jkEA+fylXSSvNWsBmzuzfvqP11quGrLDnOLHey4lNMnmZNTPAz2Pliup9e
9ONMpv9PEzgnBqCsh/28v7FWi2xGYg7y5+Ze8cM/qlJf7bKLJbvyAmLtYH1k5mrcj4EdFKeABta8
StUcWf7brOgJJATVvRQyQJy7nFshe41GeTNym9RF1PSiDoIyDy1ZBbBnZczUQ7/F/wl5sBubWk1r
T/iibyYLt0sR6zyL1zbIZdF594LzLb2XVeAjt1tWjjaVozrucHQNnrle20/1v8i7EUZ7dZwGjt2G
V8xEtOzef+u+VbwMhhKAg/dZme7ehgRs8GoFfSKYOKHc/SI89hxSwdbwWgRnu/TI1SnknkCrWgh7
YwCVZab/MCyxd+0Un5IIY1PylhsuLAbOK5+mvUw0kO+bAU9+iihKc90cqavRVF2SvQLKOl7tpEJP
0y7RfquFbgwgI13mx9YRNk04BvcpoukpJ680PWHGIk3NJlhQEdYSSjT3Pc1ClsLA0Cnaott2nvhe
4wEclJh/haTLsV9OVw45LpzvgY17TfHm/KjOvzAsskCCc2GPAh+YFWTbAwr6vpYNX/zsHg6JYwrZ
WPp3vjejBa9S6njcXHucSFz7+6rzgkMMm1d0ckP1bk3Rzolt57lpHDBx4cHlM3FQlYIeY31WT5vo
mwnxLSsn5snTBKLKMZSC4HRNy1KJ7s+j2WxaJ7l4fHoXncuKDsik8WXhiA4+IkHvwdassHRX6MSi
TiMkAvhYK5x5W6IHR3gZ6XyJERaXv+MfJfkV5GLQEwU2bghdW6f8aTlMva5d3kWBiEp++6dO3XWc
tgMP4+UlncINUtj2/IyXooawutHO6c945eQW62e9LFACyZH37gTBdVGYz3SJFA/l5MoO2/RDyR0g
Yd1rpZpFyQ98kP/GMOZ/CL2qxLjHoQoXUtvc7LrAEHbJxi1U2JLppQ28dyuALU0jxu280qjdxgVL
oeE3GGa+YwQYtb/FtwSrKmTovXpbwjG7NZpoxmN3+4dAZbbPOuPUXLQppIToriSSb4mB6UCaNXnF
EMbz/BN+O6irbwpSh1IddNMhr/QOQ74H2/QFqQbA1120RRDKltUQo4oGHmRgBbfcr2bV5e8g8Axe
V1IFoRMv0GPwn3s5m2VhclV+BJQiqh+F3QahKtscLfw89Z0fgyMTKQBGG/e03fkuTe51Gh2gXSEs
bfWTNq6QiMRY+fYK5Ib5OEu+gEDuensgAVE9+igW/iRpfSr33M56cfyuXzN+FybuzLD5dkQjc/nh
HmJkkNeDad2Vx1UH/shx1Bs/R+6MmMAssSks+bmCUIhAgp1egTrwr1L93lWqnnHSlZw276hq//pr
n6YMZCvnWldrZW9T/pkp+PjWySC3Be4DeaXI2A65B31/3GiAK5SccHtO+w7OtOGBX4cip+ustZw2
g5894q7cwc8GyYUI8XSuxeuj2J1QQEQW0sUSLNaVWOO97nJGFThS37OOWRl1RhhpFyVltCFztUdM
CXIiY+qd6LeLhO9omz85OAimY0M3Ht6nz9+szWjHAFmJDJV1/MDMj/Ci8wFzuIsFrTUFOuo2YvO9
drzAQKjG5uQsgnCzxNzIud1RxBLmLHsX6BuBEpHUDqHH28zf4BWl69NgdcVV+WMAqOeziAoxBcWq
7SckwPQqarqCLCq5Z/usQVSgtT0JbjtDEugzCcdX6/c/+kCtCOin8mrYhsmcuSBwKixSSPRyXpoK
kx1g5NMv7W+1SFdfbyrq0at1Nek8bvcmrRWuqLkfDsTtl3HxmayGW8xyHCJvc9dhCu+Bd+W3zC0z
Urw74p5QcNLzW26pfxPWBpdg59SNt+U5zg93yb65vfWqoJGr1OYU03SiQAbfsIidgR3/NdIVCgJc
uGlQcnPz5VR92d4qD/KTUo/qpYE4up+X6w9/+YJ67iXle5IvinmXYQLHjlJR5Fugm10SGcRMgyk5
t1Uvwj4xj5uh+j7dwoDDzuIDDN2PHHZrdC9ae5CbLBoZdm8fpHx6D6aoFgPzDjzlJ89jbNP9nX+W
s8teOlDoS5vc+5ZIXEJv8dgndRVddH9MZ+txJJRW7sHd3BKIcA+URC6uNvoJkoD3w4zob5vmN6n/
r8bOm+ZbjVFz9k9Ie/e3fNSwUj7kk+SFIGVR3WN6mkACd4/0FI0dJznCu+2VZHekQ0Xmblbio2/t
UK2UsQCjaZQEILUEzqJ6p0rh8b6ZHA8HsgagF0pA0uROg4wZQ2zyTrbGbDWNkIZtDGtAtvsfT60J
jBrokj8Bt1OTCkYarzO4oDWaEKII9wYw1WPiG8dMNgI20L7YK+x83g+rREo3aE5uxo97v2a4ysNv
IVmak7SnnCVYUT4aBrxRqgHkdMLpDVbu1Taj1QTkIxV1JT0xkV314xwP9gD5AgWBL4WM7aUiHVqf
O8Qf7XVFAdpDM2UGbtY+RMQUhSBr7jImHRPSwU3Wc1tBwqjTi/ph4HhvQK4OZoMLqncAJZ8x9FuV
c2j7OfiS0GZ04se27cg8+GH69LtqaCI639spUAQeJv4gzdGQOUaBMO4Ls7vgY0OfYekMh1JQNsI0
orV4Cai8v97KNVfuiWuUCoWV1FAHsVaGNf+LkQLs4UmtVaYs7RiCOrrwS8EE/KpwAufoZWnfNN4K
irwiI7cv/i1zX2GkneJmqU4oOz4YxtbgtWj6OipzLcoQGuxblDVnCt6L+l8v1pvY2aUVMoASNJ8W
Yhfj/vl1mdPiQSJ0EMl8mCxPh6Qa7XAnd1qjv12nbKUaM5BpAc4kDHoYWn4QEvgOMWF6cZ2tNnKL
snsiyTKMXR1ijiwqJVCR9rvThu+3N4+xfyFo13tROb7pbOIHODrMc8phenxQBDl3xhL8YR4tgUJh
ZBwC/P4QWGIVFIqo72uiT+OsifyqdkeuRTKt9Ahtr3lRRN6Y7j/cLeiXSz4ihfKTLw0CGWWGhwHN
58F3AMKUGPSqT5HvYAF2SJuYrjY+0xXQUcXlNzNdMxJniKGSyl4mXipbIqwBD9Rvb+Df2O7p0SBz
jAOVZXrymln0q88wWZ7QYpS1h2QpV8A4VW06m728tRAQ2Fc17fR0uK3oblNgfeXiFuMzqDsNhZ4J
luohHhml4SZsQYesBaP0r69SFp7TBraV/I6lYIkQ/52OCNBBOUGzGPrVHF0WFoOsPkDWpiizUI9S
2FFxsg9lQfguysL+OSsn5DvhyfonGoE2G7u3jFqylfDDYK8E7fvx+VyvdPURzlMF+ozC4W1wEqQf
fmjp2ip0h/aqcs2I0X2rJGTVQdxATdL8XOpo+mmo86uOgDsvxRUrqJqFgY4OnAB2T2XT15+iJqDM
L+2Sf9juaCeYdKdwXMAt/m7F+HUvjJZXjtqvzcEKucorCPdovUT5MMsTjblxHQ42GtSYhdaUUf+1
cOBfYFzG4znVmUv7JOIokpOnXcwZkpny86ZPeE1iZpBUKjYuDmQgyIJugCZp8yd0CNweh2Bwyr6y
yjvEK6aqdyFO70M3ffimitw1r8afKH4FYe+fahkXUH05cOVMeA+kIe0+DbfxlRM9zfrXcjp3UTl9
SusfMvMbTpDe2cJhsFRvDXOzd7qVCwrBIlXZyNbjwWbc8RoBxLDHTOqK1iFGawkeILMPkjaXNhf4
8bk8KKCo9/gcukLHS4FXj+dtegyuq8oxWERZGmKpGZ4nDg6wafFDmvpBwAmBH2E50nPRtq5NtzTL
Nu/MLFPp6l8RyctNDvnM2KcmFskIGGm5X8QAlJDIHPpK9erxWGpZQWIWtMdsld8JLFmHD80y/a4h
/813llH0/WuLbjtVrs0aB91hikfEt9jI52qGwcnVOx9g/Gj5sg2kKEhTQ8Rk/+zYNYQOiuaJvi/C
Sm7iD2BCnxnlZMNFs5ZMf9s+HCsomFgIFCDA+kKqkkk636IlRIDnA9q5djKGyjpMZAxWzQTCeHiC
6EKu8xSGku46hv3MDmvoPiwksEEQ0tW7HgjWxXg/iRDX3HbaYpgPjynqsKYST1ydDLkeIK5ORbti
E91r98O9e0f/685gSBhllrZG9dk8OQ/SmD6nrbXgOar6eTKhtX21iHYo44KA0BDA3QU+PX5aV4Tu
0fxnlY3rxcjcJm+b+66y+rVWE9qO+46CAMFK1riYCnQId5gMwAd/cNeHgy6KEV0VC8cId4outEvt
3kHkb4U5BOmN0HksHcRkubbZGH4Va30iBbIK5sitxVxxkEfdRtnGu5vopwhO7TcPLEK6Bah1ySTk
hr0KufuggM9k/mpGfhLobGi4fKq8ZcT1TJed5vfSn+NpkVoE5mZV+MTF6dhylRkZ0DtUe/nUNKcY
X2uuktEXQqvmiZIzIQNb7EoRRYfRGbY2a18PpXlYTnmpNaCn0W1zOwRAwaRmRbSBmMz+k8N3cEVx
WjHxdhbcxamyTWWv7CjFdG4qIdRTUXhyyL5H9Fh3CbAFd6n6X0M4iIOq7czP9P6ptrgBRP8n8ver
4eVaSHA7Lipwv5Avywsl/hjNoR4vVyfC9UjLL+WVHMABhGNtNCN+DhQFYhK5MonamDAFXmLRjHh4
oLn5N5Gv5SLgl1QqJ9Y8epXFYjZDorfTmUAON/bewURezKbo7782i6L7Osv+gDwbe89Dc9BHmeiW
6XAJHPpaVgkZST29yDGmfpbSY63pVpxQfmmvyOcTbMBNHkcLOg3+pHltelkFdfvja+MKP4wgQ6+k
D1ohbE/adfEpzZqBb0zbUn3PrczdoyI3VxMmDaCgwHMVd0cYVzTEwMzrFyvpRrgDdXvCDAFQqN4f
u2w5wf9S9K9Vi8iEKoZlxRfHXwQ0tfOE8nmAjODcQHhxZYVaoaGLxZFzzCt9Z4ndkiq20nYmcLBX
0hYhwnDmrmU6dWI+Ud4xwDd+tmkFYPV3OVjhBb//WNf+ZU8MZF1UWmMt9ZQReVrjBQQFvXoqtw1a
ZW7a66yxfhBoIdWS7Dw4oZGpgty1knt+tZplQI8wHGv17lp8Hw+KXSVSA6eQI0+6ml7aJSihbUkd
1sSBJGsJ29ViM9CeREn3MA+4Rw5JTjWs+kPIEOlrqWY0BISCUFSzD3JSwmyZWqJvrv+NQZCi8AXB
ETvJYR4ETcNGKRRwKNRfjrX8n9coC9cTs9O/L9hHIyozlfQw3ORh0HZUopcbRcnQLIls82uy5t9g
F0Lk2ZGPVg4exnxj3BRc0xq9F2pQdJk6fopj2vTPkAnFCV0B1YTpaxEuRRt1V9PpSmGnk+9CwWcy
vBcRmHyjZQc+dGdATzJA1cXwUl27QV87a8m+26bsCLlc3Kw2SPs2DkiWGfm6GxeVfv9KvybNCl3S
4kyZw7XBwaHKuI3IX/p/GNZXNPh77P96zyudBBqjGOWkKnDOVcaMbXOqPdVKnIBdSV3dT8v4nkrF
gFKffibNpOiRgduzFAM0dxKdPl0oZwB9cDyY8i/ca72KUoFDOTVj3CkFTcp1JfJ7xrzln7iD4/BD
1fyIw5o78k/vqpvodprPihfE8PH1zpSW75Jm0DkC3CqbO9GpbcJbUXfT3uijWOqmNU909DyXdzJM
ZeJ87Q3hv8XppohhrAmIeHHsMQvKifRKrgQxfY9m3ODfZeEqikEoYk9XtD3sCt/8xEF8cjBXivjy
IGZFdCxEx+jP7zdcUTR05H/s7Oh8i9hYHSUE/oZ0jCHr/p89k635buECRjYxc/1DQzPTolbS19pK
Upi50dI0gq4AP87o03HA0bcopMh9p+3O4e+G3Q4RZoJN2nlEn26hLfrcwJbgZVhSrUOOAs4BuJQE
Fq48tmL9O1KjH9Dn3Jpp9wYu4Ijo8RaAYMW+d8T3MEkKnIIbpD1mNXyGVPr7aEZVYgAyMXQSgzX9
q6HyUPRrTUPZaonuNvrG5l9mFtAXN1GVH3zoiP5BOyEEcyRQR7sGiQbdgNmAWWscFs5swKHDFFLw
eFoLTKyKVUltydAEc1V62T6MHqs0xqd9OUJIwixlAaimSqqC4OqONiFfqVrEgSNK/+2sx4/0HOrO
IgrJT1UUSgevWWd5UDXMwAEH/O/qU0eDQCbJjaqRS9+zSaIOXWc5900GyJublG4b+Vfv7b7w+m0k
4H0tw3Y3cTvVif/MTqY39aVcfmZQLOBpEwo0Mg6rzfkhgR5oZH+4BRAcGEddY3N9/etbQz/P1ZPf
ZOBnM0HPzwA6zufZRGy1QQguVPTF4Zc1joq9glVFkHNYbygzyLXl5yvGKdGNriBozcNjzNIJKFpO
lM/XYgG9vFjgLWsa+O8mlImhTZAo1XZ2C4NuSXXpsilxMvTunFLxWT4nrq/Usmrquto2JpDKzbbi
R0SXpt82LoCPvlyFQ3DFBBnM3cl8LjE3rSyn8PtgSW4ApHSYVZsQQZMMwryc7JXkC+/5v4EAnDNz
PKmgEu5Ieeqn3QQ59CT0C/Io+n+dezIHbKF3w0r8jZNvt0xBKFRzncl+xv6OTVdiCwtv/Ty8U1j1
dHz1tU//M3eNIAtt0HEZVVfDah4lN649ylwrh7UxQCkHvpan7/DURVMzgaNkjYoeR1Wmaq2F7xps
rg6+EB/cEo0iKcrCqV4vH0Uxebk7BoNEw+zP9fP3WU4Vl7v4qjRsHiXPXS8udxyQFfeFiIkttNqu
t/XfJJBd4ymtvneMYpkfViYGfaituO8pn/VDK6skieZhlS26Q50/m84k0d4rFbjyYSgu+nN6hVZN
LzBhXbs0MQbcAJwO700rY7TTWNeehF6sfKbRszRoR/PHoj8TqeBCMNnAJsnD61AIraizqKduKIxX
QyLtl8EdbJSOPfK1Qran2jJZkEJm3nnWRPwwH1dScR9/k7RTgdZer1xM2kFwStN3oI5A8Nuv+3N6
UwYfsU/fQ27Q2HNwz0zsJAFgLyTVC7003JAl3TEFeOxgrZbyIYm3QDzo58ol2u3AHUanDX3ANln7
RyfSpNsbpAr+BL5rm+85jRHJRz4eN8rwpBGOwMf975e8vgLaxA9ACvlQOWCUQC+J2G0InE0OWxZz
g+O1+iN5bwfzyVaVMvfJIvl6YFQokMVNexaD83z77x/gYPO8F9rQhNfWKnFvQOWUBezqYG8JLvaP
3O2FXnD3f+uf9UYsntwEd/Or38r8lGIJsszqTWwORBpPahPF8ySRuuwxEbXw/nnskwRtX8i0DtxY
ML7LXYxnExnKg6mU5OmagjT2x8FNrdvXtuGRgHQtjD0JaTjxf3/UEIq2GFeNnimqb5zYlirs1bNc
FudxNQloac9rAvn/5avd3WNMsdx1c6nQZkx89xEedTfg97uV2n2itvrM0OLDbBWGpEPCeeKqRqgO
k7xgzqFXHxEDVDzurA0Jts4G0h+UJ4hnc083f9jIoKAFn8mt+SoSt3VpLbsSOSdD3/qfXZeWlc7P
2qxKdtcvLqQB/cPtta+Knc2BJJCGmTx/zE/yTEONRokAKikrrvWeCg2KiPVV/nLTZHWpxAn11upm
Ay4aCMNGLbv8MIhyXAV3SE5uFy4lhOeiBAkUzNVO0tXryiQjdFwtPWPbXbvK7tqVK8Lc35Zz9Ud2
DW+Ji0mLlNaPi2g40UtA8RyYqqOeHBl7fPB0vuZ/o2dZv1CN6ZGRrwmLMNb/kXhb+XK48FWNd103
p0hKvtT0HIrz52TDJig6PVGNhfiRggrNvfmNiT4FIlXNDeySQsJMSM93gxdfNcn88N2PbbuPZiz+
ivMJX7x/dFCwe/v6W2SbNUci6T0PkC6W/J0P2dHzmoJYX9BFwa0c89hYuP7gr9UJsxDDT0AmfxSz
kXucSg/ibj+nQV/ww0H7seBNw0LQRrl86JgsZttiXoWSfOAVWTKc52HVj9Dl98boQXR4UqlgHEev
pz7wU27nY2W6Ac19hcWbmiIZcEvWM9DHxeTtlfsvTieiTlxZrxfvJRMtx8o1Ri2BWcDNie1UmKPV
mVipSZlQsmCfgFi1HDzYrgT29CalvIa5RtKMC28KG6Mu8ZnNgoh7b69dccQpV1CkI2QDg5he2cnF
5SBMi1MOkAwsSugWC56GESu69CwJ4jjDShencHBcxJiF6MVhlYIB+Cth0FOp8fRCQflAUFwHGsBV
3Ip7ydTgLJQjVhzRPug4ixwqArC3ZCzYC+cN7LDIOFt6txgTGSMloEmfzuiWxJ1768k0DkI5b/I1
O0UEjY2q80sgAurEWzUphNlrOm6raMaj+wq3rn4PM7U+30Hfw375N9+1kudRXyr1CTFLE9pU4y4d
3RwarGdhi4wSWvzXmb+SAsWRo16OrAbDsNLN725iSjdMbUdVoxpJ1tyD75MYmWvnWPQt5io2MGpU
Xg4io22w0YB3wVFF8cOyTvof6VPNHJeDb1Pt18gRH+MadJK9fc5WztY+GRxHV4YiGC54VZzD2DLa
KblwLSmpcge5jt0YzwhxuxF0AnU5bkdnEhNpkAbF9h/e6vzflpZucuU5gLp8Opifm6MOfjWTQb2B
nz+IuafAEFFMW7WsLXiIhaWHBlpjH3wAPtby5FAEmTch1BkgOmbNotitBLE1lmM5SWcKms5oMZyJ
XDD5bYOqz+DUnfSknj9nrT6LuyuVwnOPuPKxskKiuul4JqFP4eJ16ae9nsDm6t0ZttGAvZRAI8ff
LkRmSHZrf6dQlZ2yP5i1DqPaVFT0lcllZO6pOsY67a/2p8nE0teqKCzk7ssfZQPvW8j5bTEBhPkg
WPjaiKXMOwBCJU/qpHWRsawfFmvJMh/jGfizGTEeZbbkflNPrOOytu9NExZGoIlEo3KvkIjNQTo5
N81ZYQzG3Aop63aEBtglpe/72KjFx2mEIiHH6Y65pPm5AVcShK+DfSehinql/9G85IzNUM4wpNFB
yhwz4JX4daQXEWBMQzZQM0+J12fVxSs0dQcf5QCpc1c2pbTSk1Tq9pwbN9k/0gkvZnTDhFLLJddy
KtF9e112YO4wcRmPdZttPFUezuAha1zNORdJidj4+CPHMtzsvzojIu0xqAOj/R/B9MjUjtLMzSWD
0zCDVWmA5diliBIXeRHMgvIV1pXcbDlrN50YiGWU+oN7jB9FJC1LVbSGxUdJ17AKcsjO4a4EvWDK
tsIIFpatF7SfY+Yo6sRlo1q5pXBSS4WEoUUzM60nu2H2Wjl3L6YVzH5erP5B7hwatGKzX2guy1Nj
cYixncINvufkv+xwEbmwcb6O+zxJOrS2g5Jyd5Fr0tDlHfcAbOIxIoizdGfNFh98qO4x+v5WmnIi
MLFR3dKWSdimTZmpq4rJRj/TKqj1D/9dTQhN3PMY3pcS4kvnWKyMwjaFwNSzDt6RZqV8umhqSf/Z
xQgJiOpxJmNRXgQmV6YzLm+UJzDpem4vINLutqZMUL/HEfVUpMrRgDlgDDnQ1NxAjFAp/2hJze8Q
1s3BIPkKVpw2Rl7uFmJ9J8qRmYLDAN07z+htafG51NnYycy2n3PInNR+OT1MnTLZO3q4K6uZU4GC
R/bbtmZjcubqneo+RvCfN26INea+lOIzqCu7A7sqJ6+OzHhpD0Qx207pLXuxEfJ6jfhmYrh5ovQK
6ncc2h98lB0eJkdoSds9yAJQkWy6eyp4h1M4w8I4evWr6UTC+G2K/pov0lJy5eJ6uKbLceg4CJwi
qtcuWcU80/dsDMwaZueUcq2XQcYWSPienWm14DFAYzmjo6CgwxOlBph9WIcuPVeO+ZfNGUG5apZz
/dpqEC4ykMHlZZcWPnP12QQwb9KH17iT9Bci4XT3RS1+63wYxn52h4Xl/OkY1WtnSRclNglbI1h+
VoFhF1Mei1Juv3vTJaLx3/oVPhMLJXfEbNektTK++vcocoUC5+Y5kfqKBVA4Pn604B1oTRLBk93+
nJBMRf8/7fMRg9X8p8BpIm6T5jB68lhI75LYp3Q5KMXWVFx20A4F/POQddAG/xs0ujn10REBHRYT
B2+U4OHS8Cs8q26noSYNH5cqEqKn/Toc85jwNnOkskPsjhYXoqQbtcqpYA4aPyyIAtvKqF3bNnGf
Hz6xHHrm8agqpu0N5uEnJJ+04b+YDn+JPB/rEYuIXnySa05Gz0zVuLfstIvqahegm4YsO6VEi7VP
YYUVWi9L98CM4vZuTmIKknpW2A/XfBY3B1aRUBtYP+JAktn/3+vI5g9sRk1c0OwOFzE98W1sOsUS
CaOahFOrQQEh9R8xaGsjsx9fvYjWvCoh25j90KIHxe6iVOlm9AeCgy5+thHOwm+pyVAJuEcU5/0l
r3i2OGVSb+SgwU8ktkh6oY8l3og0E4wntyJOBR2hYIrsJXbF5cdb41RcbSWAa8Ub0yL8B60CezCP
kDngS5BLB9Q440OtX9lj0xZGeOhZ2IMJDEgciR2V3E50QyPtzrsl+fxfRmId/58rDo4VNd+BIg3E
dPIvpXDXs3CgIEGutqkXagKzu4+1aTLlNGGYRRRNM1nv2oo9RwpvdMuLIbkHcGxliy9xxGYCwYBh
nVeBKEry0Uuw/qY5Ll9C0H21BlMl7EcR2ZZPGlaz5KihHpWcVNjxYO2Wx3RP3NQR8jI/IlNLUI56
sNpCjbmM8mC4A9E6iFrVNjql11xqErgeiGLPlm8H2fug+MHN/rolZxV/990IgYZ/63V+Rgx05k1Q
akTPvVUz4yUQ4EA284kKx0OflcOEDfWKZGpBVCS9tJuDi8ppepeyITphKhdgrfnwkz3M19/sTKME
uejfvlAXK+3d+hTVAPG+sko/osKKFQMYGJ/6YS7j6b2rMwmMPPoDNLZVmhNY2484g7pYNezy9gQA
T7YbyVlX/R+KjKESTbPTQgX/cIYqfg7aVPO9rkX1BE/a1mEWdeFkPKxls7PnUAoqDSpX6Ba7Zvp7
YSEePg13qq6A69FPc7LWTSARkylDzjOnLgVOcTFHYnY3MhiZlqkEzvrYrdVOnTH3GUKRWbijQKtX
edU/4T2nqFWtGybwf/HZ4kJk3QBeNiP/wqQdqOTwMf6MR7WdkBEWTSU45n8NTssGBIjbWXr6FJT5
jn9/v9KPzJUyD7uj3QtTw76mHXwVJ5l5zPBp3p8ramBFCGLcE7PT+ydqcME+/TqOUat+zzu5o5qa
CL7pN9ps+KYXnMf296JWgPrRJwyptuk7kBGoqISNj+zeJBtgcqQbffM7AQLXjH3MrTFqye/WGLhX
JLIKTI4InDI+7Tj/3P/cEoa2aalykBnoquQKJsUsdbbq1cxfcDzkxwCxCbb/iNNs4KEjW9Twpp99
lngNTFEJfWrJxHy2txfl4m4iS1sEqZdOcO5x9IU8Esnuz2Xj8OfzRY3yg9C7AKgau4u+DN178gSw
L1/xpdqbamEy1ZbprYsmIyEhtPEv8eMN/ciCJs37FzkzVBQ2J98UUHhyaLCS/CA8rAgEuDiOYHF0
+NxELA/wFAr1NPdEEp3OUhmdWQU8Od+haQnsl/nD+fVzUEsd93YoiA5w+eBULq0LBneTyA1H3xjj
tBDkxjddzbYIEVrgT1YdPqW4PQXdiplU808RrEAb4NDV0PxVvIqqg66Lytr+2aR2L5TCVl0c9S1m
uLHfA8yIZpifu5bLbm02aJ7rTwMugbbxU4nvwhR5qVAw6+mqB38Pe4t/2XYQwLresJTTztST8fnp
dnnii9QrVCLyLGEgaJTjMp0h0HtAqX1frAZd/zoxS3BCyW2Q2ptNSMtM7DbkozbCLoBIstggLXYp
Bzzl4/uvOlbr/wdSm6QPiDOdJz8gf0o++QPGX7ngOg2+rbGlBINiM8tbmoPRXia3kUbaQhNyrJ61
c6JNxXf0rwYh0vdeU7yAR8vlwP6cdpdNQ/4nV0hth8OT4i/Ln7jbEU4KA9o3KhMT9Zr1qFL67bex
pZnkLbMnkTcyV49TBbvEpG5uYCIN4wX2daI51L9bn0iTNW/HLVUbRPgKHeY2SMalZ5Cm4kjX2td5
RIFY3rOtTTDBF7ITOebLNEP26IM/jyvWHXvcUbH6ta96xTpcuf76UNsz5BJ7KFwKogQIUl2Y2jRx
q0c69egBgH9M7LU7YU6qmVMK8bFbgW3BYCIKOLwki1HH6B7C57fQ13KELtxCf+yheUGMRXye7EHI
aNpI+Fxf+pjz5RczfVF07oFdFgPovjkHVOT47NbWt2H8Lh6XVoID8ePlUOKLadWh/h7+uOE+oL5E
08ziYXeRnxsO6g6uHb4UgLAu5sPCL8WUOh0PmG16nN5AIpL2SjszMDOS75HP0dp608vHklZL13aK
q/xlWUU49yeFQg6kSKIDpD/8PTkctpFPXEnRcKjhijK6SXGnaFl5XrByZOyVIlQZ1QHhA6yQvRNx
2ICdv+wPcAUGkU3907thEaY3NLrjoetnz2Kbbr5xqEZGlLW/DtsEhZLWxUrlYblT+Nt+66p8hojD
LIBalKHZvNL1NEihwkznnVm1bqKq3mKQXxfd4uP3uFaMa6UqOJpevQPTqp+9AJZXeB2pd2oRwAee
Fd8UBbSjHbYrISeoaT6Z135wyAeIWBzIbqmi4/4UYB48ygb8y7fv4uXrlGOnm9Baq7DQ5uzjlXOU
deF1/MNTsi0IruJ4Zvya9u4KpS2cW2HwplyD1Ak2OYlklvSR7kHQK1h43kiFBv8cKfycDzhxVuty
a1xt0L+QoAU+S+OH0Sz0JR3/06PVmpZMhSAhVq/WOojkKQVMbVtjhodotLPoXWvTXrPzMYDRqFd6
tuZcQfsSDhcxwcLZayslalGtH7XKs7QoxFckBQ+j1+shub02FN6bSCVOGtINUePxQYLx3SST5XVp
wKdmzSVrN3m096prpCFBENV96lVjVyp9YATyaSbV/sIVplrBRJksDtWRF+cz8NsivkCQDWODaEJ0
GhJ2zkXB3d9UnbcYv4R1KadM8BM6Us9Xz1Huc6FW82QQ79tDyQp5uiiZRJth7jMDqtvYOttvgIY/
c9WKzK60nm3cUo4c7bizH+JLeWyQwZyz8wAamAa52i/eYJo6Alem2n7r021lFORvCsa4htn+upiM
C7K9WDaMuZVA1jzk9cQP8O07xCKSkIVi4zC6zGceK8FcsEpPXGCTePtGnn+bJUknE+8PV2358S2g
DXfXVovY6nraNPD4uX2pdeJ3jvFDmemR7xnCVfbvI/rv1/u7swOB8CUu6f/F6RxYSlHjlrHu7oSM
gVvofUp6+DgNbu/vZmDWQOFzU9i4u9zh2UcyHTUu9ZG/2bhsJkTCaTbPDsNpQ4/fRXyeOAbSdZ15
jvCKJQfjby/OxupUeIcM7ReDD4Hansof0M1I6lkpW/xioj8E0S9nEgMG9T2pakXosuemBuBQ6Tci
K0TMrq9krtXD1DIk0tmK6zGEg2inCzaXE2v7jfwlr/xbONd0X541f3hiIQd0OHKLh3bCMVNERB2t
l2OkLy1OyH8vAa4mEM/r0cAm7YdA2pra48t+IPNz2aLKfiuab3PEYbI0AQ1iT0hCpuoDnBHO1ib2
gQ5sIJvzK+1eG2j8mKR2imUY391IwDlM7IxOfXm0OSMp6dRP17jKfizXmwdarcdeW2OIOplCHcRw
fPa2xqTGEHhjRyIrHGssHWQfSH3WqvJZdMkRxMywkpVcaQUQPywd3RwMEHGVQj54iuUpCsnkQ7g4
PUwDDgib2mKdW8LK5NvRLODK/jLD1bks0g4T6T6MoYQ/ie5NKILQlVoVONA0pCBK+KgYbRocn69v
kE+KL8vhUnTWmxN+OIm4Yv8rNJ3vZUxNFjauYIH9/w55LnDBa9Ghne0SQV+ufWei3UfMd91E08ZW
6xqGeF0A5B2Ds2sVZaL3YzW14XWsdstUDVkKjiTSIEAEA6odMTNKXA4N0pUX1elDOhEuVcigBKsP
N2CKMwURYZqDzJ7ILTZh/74e6kGmvpcxNawhwI80Ra97OZrJyAg90bsDOoE7E+FhXd/oIPupdwmN
tujobK9ptN5HmfMfH3HrW0na7d4P7+kQCa72naXiictz4aCeOLtr73iDxx9xJYBw4X/i3LX4FClJ
mBdTRvx0Izh2zfRvr7A+XYmAQR7/umnpP3+ORv4AFvJrK6WWRF0Fq7dGNQKVH8FKftvkNAGpGbNe
787gx4tdECdoVCQLNxCibMM+rnx3YxmaTAULgFw24J3vbqSl07QhuhU2BSJ6TGHoy7An3Czw/lke
DizTguVfSGidOk14k7SZb6Mf0CIqPUTmq/jlIJGCCx/yEqL7b8rmAsydPyNMb6R5/dbnXFCDyxjp
545Wi52AZ7TPgN+jihUeNFhGWU1x1AFU6JosNM4dVlwVmZsX1hsZALUVaujWDbg7cO/A4SroLnwd
9MEHxtk7/7/hyEvwty6YMj8g1UM6kOxqHoLkk+vycaEiWICIzGm8MQ/+qfLfVVpquMVdD3cz78DC
in9OzFDnECMgQBDLrhN6dYDhf9y3oE3nONkneCqR8UJBBwXghRYM4Axs/GqMSZ4E+BVylQWcnkkP
bhPGPwCZVKXzETPMLyJHqurqiQac+Rxcm5/A7F8cqgNtUoKOfnz/TDno3Yz+NbMz/fTm8H2YBI1b
mqHh0I16CIfI8hlK6coQ/ky1hpyx2cYnK7wY3pDDM7oX0Ten/IKyPRtsodApNRDcbFja+p385hD3
pVy5BT8SujMgLTgzROCmjEm5Jj7wszkP3ywGtCmoi7ad+pfvAZ7LvNHB2wFk0Kk4PrXr1eLl+reg
VpzagRNDHmKNNd4I7olc2CP9pCFtZ1k3xXj94tZ0H5oeSgdd+9H5NtWEUQdQX6bolf6ZnAVT66vj
gVjIjMLC34lXoV0FgPkOKBIL1JsAC220Lwo4VBXZOEbxJx9hjFh3U1i/1vb7VyJ45HBYifX30kWz
nx4Ww57+5DE9L3CqEvq7LhSJhQjNe7HcxoF8gsf+n6I6OGkFSegt0tblY+gVLwVQgNWdUh/Ea+R5
1zPN9bIZjGbE8tLJ4C83o+cq3JiI+BZB20lbYcZQv/sHBbBImv2ZDsIcwmfisxvcEvXs8qxezGhz
M3ZcfvouwrlN+RUxyxQxgGy53jRPlse7qcjNT9TDpxyHcDBOhkpPMtnuvOoPM/nSzTMEu+chlHYa
Iv9qQzhvJqw2qTtbyX3/3opZSJhiK2P55hvrwDfojW4q4zJz7d4lUziyaRA9xvmLBn4BNv8o3k9U
4PASYDTY2AI0Y8wCEEVJ554h+4Dg7qm3Q1k9yRo7kLog88md9YBJTT6S7Se386SV+anELd6eNQT2
L2yTfuR5lseaag/Q72ggJDwXmB0L+kcNgjXJKIVZTLjZZtiEfOT9W4dvpJAmlWdqse9nDLvsQ1Jx
WifbbSFIOO3y1Mtp6Ggen921twLyDp86j4byQUJf9sWwYVW0/aBUC11zKGygNEv7T6Tja8du2IyJ
GWTOdSQz1zygE1mG0mv/bVZXiPHO1rZ95fRFegHvDM9Ku9n2Kn6oDcSD0VeMW/vCAJ+8Bsn1CgP0
l/kRMuTQ4n3lEr7aywneF/PGD8hDO3VyrUm5vjQDn7J6I/KozxcLhXgXjpoA99EXD6gvZiUdYoRo
NVVDoPmRgUuO4NtRUr4g8wyPyjqJDCV5tQA9+WcryPaT01o540mBpdqZqSb45KHSZ214R/To0aQq
/TgTqnchM+FGYwtJOKKyaRGa9FegJdtzOhm7Q9NxKO9WR9vBlBbzUcRSHambf/9rwhcvxajruFqQ
tQM/WifQewgTiDE22lcIA0MvBvhM+r06nkwH7u7rHFR1lBU8IIWX4sbFyj3IuG/2B3eOQ/ie00nG
1jkBfYdYSFkS0Akz5b4bPRNspBz385H3Z3uEgZmRif235Zqf66WTcDQnh7Ml7+EhiOwHltacNHYY
MHBTAO4/3HAfhu8FnA0TqFdpqWcl4B+ty7oZRWcL2tgNeZotJ+t0DaB278dvqdR2Bl+0QHM8WtxT
lfTVxTMfXt9zNw+usOemf91QPGrvFLoqzrgTmzCh0Yg+nhjtyoHmM7nflghPYTTT35nKfjzKLyOt
SMOqSVtZs8rBbNmBRTDg6YTwTyeRMQjV9YLuT7Kaw+avBm4I/ZcPYCzHBJ+josDveazmGr5FlT+R
wHt8nEWTyRTiAp2+fV+6z4ewx1/iUV/hQSK6Oipm9A6VapiC0dcEcrBw2JI3n7MBV1H1yOL9sddu
A0tDGOxSHUl8JVPqzgbLB29HSZvFxBNCuCff2ZwaaiaQ4wUc9P8q/51YiSvjSgZs+Tj9TZa0LD9y
b0pIHjvmj23F2+O+XMPEYx45QOT5+k/JFqqNe03YA0o12FtKDeOZivhuzjLiaUbDzBfwJ+6tq1Up
g25tZZgUD8kTdhu/S/YEJckUxMTuJd0yVMr88kk0ZLPzkLpFHkLno3ROqS9SwHM/+7w1ue8/eji1
gfWZWMVqnXhpAwbmg8VSFRVS9S2K24rFduS8LTOxARMxgSFEJUWqFYxWTrVwCpY7h1GphkJzAUJT
09d9UPdLNLn3URiMISlrO/6nWR7JBRRV8vQjcgs2jWUrlXyvDOkM2xJYzDVlwbDMhq7Arj8AfXt6
k6WMeOhDPABuInMnXWOXceWvUGdP/sfLjlKXnVDlmumwc9FCel02LmKWfXGPuNrIBJ2vgyex9RBa
vcLgI8OeVM4tI+xGTkqF3xt9T9323Rcg19IflfNu3ekWrKRVTtSObAAJ5zktIIusS0noMxCDQHK8
w0ouQgKrV6UXkr3aDbog+dpgodtJWbMp76BP9JFs+lJWYsWTgq7271XeREO5LmLsFqNlCdD5NBnQ
4j7eiBmSsVP4iYaxzbuAiBli96nozyLHNv/rTtgknYzCa+HOlvz9lKdvgfpfoJGZbiXiwMQd4+8o
8B/mA7N0VCxZNyKFDwKPygOlEjRLtjpXT838u4RR7VsjDJ2JI/HsBU/5U8/xTD4sSnl3PJqFmRno
WmAFsdXQfu9ukEj9G6/8jFb9GaxunkaclslCEZJ0C0ep/XLGcziJW7yStfvj3vOf2pbWHev6Jsg4
qabooGoOrR1U4L2i2MW7qmBpQ1q+soh6W0jLNFJ/rFeyQHR3TWKsmn0i2b9F9Dbmh4wV18TAnZ2w
sXE7x8uXTzALPwhks0w1U/yyFGR8VLiW1BeZEzUad7dGNP4OxhZO+1hUKGtpGYYqh/MoS3EhrpQI
QKAxblerx0m0fWXJyLL1b/TVR1rgbzfbiVqi4mOBImQEPZpCi7ZJOB0it4uiIvs6Y0jMcUUNxhCW
PbDi3rYuGILZLjOHL6offyGnFbrk8f3nngYplqmqVj04ssXelgymTdhoMGDQFjKkhiurSC+/0HmL
DyE9apEeZIAz45QJsWeXICwbBmYZDw6cQBS6HdHe2L+15io5g1bDIbRqyXRMvgjuET2x37l51DPE
sDxXRFfYoH8Yra5xiZM4LxhJ9NRUndxyUMGpPGhvdb0kLEcFm7+r13mwmqPSwVpQo8tqnB3c2/LV
W0iTnT6tALUV1CmcdoP4gl9F9t8o4+Tocr8AkZaN2HQBfbKZezunHWurMD2UdgpcmfcU/of7S+Ca
l2MXedwsb+TmJ6J7EcYFLX/iBHfnyYW3DX86XjaRX9bPNQF6B4gr0ajIqdjBFUx1zjt34Q2Zsy6t
bcWff1c6mqGhqvIBQUinTf3so5PzsBKxEn2YdkrJ5NLw41E7xN9nciq899HrCj/QLXmsxAqiOnek
0sS20CYygikT01ei8q+npEF0DXJa+3/JK2G9zTAt8FPn8zikxXXLH9FQDohh5VsrvPbZ+mCoAyyt
+aAqfsrt/FlHQ7dECi61iYpPOn0ZuMkn4ipUMgjmGPKE5sSQc4KFF0CsxWW/UAxY8hj1W2LuyYpG
zTAhPgceegVP1L9SuRavLDMRW/fHDpW7LH4RLYNg64josn5gz368r9JuIXMhf+XAPabM6By0h55I
biizJTtW2en672/p0JbyIJnbkNbomtgf8y7Pq5Eu1zy2+Y4RAHsK/aBeVIGx25ZwPrmj1y9TCoq5
Ou99KNd+JGnIFJJs0jnUtiUNJz/NIgqpvp90kfYasyMduoFpjWglie1ZYqtLEVXSyb5pvKfgX1lh
fJxJCVCMmVMH6+UHB8Csca6k1dfd8ctNSOSNKwBrhrUzr+lf/MmCGXLVrFfgYxbAASeVn+HXrfQQ
RsAuQVREDl14DUMj2jZNRGTCTZr74Kzr0AsDUuBgSAfRW1tlY2NYFlOoTEwdrl+ULhXCWcOuc57+
y6Y8ugtrnwiBEwpw+Zjkgl38eyCcmSuGrRSjqbRuMYOSU+V9crfbnaR1dV4GEuaZYuZkz/he33mJ
G2f8PypAY0wcUIh6TEaNprw7dsp0kFHjjeJMm/pQ6EDgAMne082RI3+/VdsWxxG6J5kDJW1sJzZi
8OlCdN8o0Bfr6AxcEruMsk6PaiclJicd94VnEJWt1CXUDrlEnf0dC1dw7H/rdI/bx9nqyJMkmSHi
8jpEKPRX7zgEy/iVrT21yrDgMtlmBUgq2TPEzoe/+12GiH9KdmsBbpEumP7FzgEbVEehweWSLcL7
4mIt8vxhQfBpR7jwx/WoP3o84HL7Hbt2a7lebV2OvCA+rb8GZIsdvKyGaa0Ey0J9814j6rtSTt7D
N5Yj3tmBUQHJPLNsqH2iEM2vy6VBxWX1NAVub7ebV28LzOIZmEDnpzXDVP1vQ75uLxOTyeIPfTuV
/KlOnQ/i3kxjcGosouTD5uFJTZ83+jaqTk1uQ78kDI7D6JKzgsiopffG24gXmICOisL7vhiJDHXc
6HTrrSznalwpXQl9R4y6bmhFA1SJwPRavZCeoStLfsNg3IYQmfkQGHbNo3nZkubKXNL93Pj7JW34
orzwG6T2O7jKWL1MJy5wbDzhieD7+RxD4jEkeCD0aV+TAs93FYD8KMLiYUiTImJCHoKcAp8mLIlX
axnwjZ/EYkOYHVW2p1MdrrFidlrA+cABZDQUg35o8H1fo0H93DzlIQZ24eY7wJkQ89zIe2ADTlSu
1QNDulpU6fVPLoNsClO7AETN0wmrMePspAX50x/nIa9/qP3RMJClE+qbG57H+EG292RS6TU+1Vmq
aspMJzRHVf3VNwpNnib1UAbnhgs2jaGtzBLl1P/V8PpSnLxAbDGas+YHBW9kOyPXzrh6e9N8UWe/
ksdxMMT3gGjJC2y2KCsKbCrcNjalLlGfBJTZ9+7Mkp6/CAmMJqxHg70NGzJKq6eRqVLlHI43f/69
9/8MgZwjl1meeTTNn7l+r6bOMPLhR2SE10tkN3nm24br/Qq9vP85f8phD5CuSYo7L+se6ZZDiOqO
ppp21nXr3MA34Chg35Rq3RrJnmM8YXYv+ETfBnpf4+aIEigoTRb9ZXUlgZNqFA/cBOKY9qwfzQUD
4bNnN20PnCJW2Y5HKknnA8B/l1YJUuB3tuLhoNHtfmI26mMVUj78y2VuDeXyghCqzPaTWTEZdGl9
Y5PEbndUsMuU152YhKX9biv5TAlkz8To/bub4z4fmw19HLXNQFr3lJHbXS52AKj6UWYr84vbuvtl
uLd6XrcGHt4knTWcr5IRiSu9vgyaKWqIrgDe8RtUjeWaYrXV7IUxoGQ8b9OOaWrzKHT7ov5/Fb15
qbeea0AGNWLdFSuKS98mkxwoi0qdnW6KtKVz7ieH9xToV4IxrEAp0qebbnAXqFqsTBydi/g5ZuSr
TcMtINLcHdmqGnlRmMbQ+iljUShQxCIVOl9OkWiUmJDNi3qgjbcmlbwDQnzGSaxp3IdiGkF8iBR+
2RL4+8p1ghVxOKjjSrW0Pt14zxbRVX6NWaU+WFVOnsS/bORss7YMTsQTQJcr7kNETA8yiSwC0NGT
WeiW3qlthrvEt8Ghg2k2Xhs2IPFooEN6sm0CTF4zENAjj+IqhQb4bnIJ/QMlhHUpVf9WdLpoapu8
L+iLvkENvBQPz8Nxd/jYN953AiupBgDe/YL39JuZUuNiV3pATcZWYzTVBEcUptHR3C7yKrPhxM4n
WjgGXY9xy25sntXTBHSa0J2v+IHhIvRbTuPceLVO20tkx9gkAzAlHcH9gt/NMGyLQqY7gMrnbg+W
MJbuLhMXfZCpVvEkRIBkWIaQdIPy+RdeQwG+JdirEhvcqzsviXNh/ZcAG/GxL6On39gHu1vLlB05
529O9XNp55cpUE8i/ej/bBi7VX/cOGPT2pnPWkeyreV7z1Wt4i38Z0/LKWJVEZcrzLQ1H7+NzVz6
qW3P63/QEUGUHfQQfvkMbkEt0+xVK0pinjNgx1irR2tF8Q==
`pragma protect end_protected
