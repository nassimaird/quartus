��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_p�x0S��=d8�F�y�"��s��	*i4��j?�A5���n),z@�7L*��b�;Q�{Z�òs�x%�Z��g�CSH����l�D3���٦B_���pR%i�/�eP@�}9�@H�̱��u��q��^�Ol�H��G� q��|ީ�DJ�]�Q�;�B��f�'�X�tz�*�%^��}we#à_]>.�)kqN*�|��"�����z�rB�D�O����R�M���Cem��q.lL��4)��(�H.;>�$.�^��'D3
tc����Ԏ+*���=_�?�86�/���*Z,�>D�;�F�M$8�s�`M3�s�E�XZ���MPP0��v��0�T9j�r��ߺ��WI[�ɛO�^ܱ���3�BH��a8y�R��4r$����^�~W��)d\�!�U�8�� �©�(��d{��$|k�G;� 6�3�����5�%�9lp�EmB���t�u,��Dmh�O��`��|q���q]���i�S��K�T� ��1$��)D�>$���7>��h�0ڄ�<�&��u�����_d�>����)oW�N��T�=��m=ȑ5�����?�8�� �2�>�i�E;A �e֭<��.8E���O�+����2��x��H���7���ΪR�m(?���v�^A�6����o�-�f=A�
 @ӽ`66��������V�7���TC�3>����yTĎg���|��Uz�b?�ZE}�9�a����N}[��a�Z*]ci���æQRW�h��Њ{��6��>�q�v��-����S�i�_	�<-��4���BȆ	���s�]Y'2;��*��d����(zpWi���)����V�n�����n�K��A1�h��
Ք�6�2���ǋ�Jx�;\àJ�L�u�<��r�����|)� D�1�b[u�0(�˹�2�Vm�kս/��.pw�,��aaK�0�+�����/{]�bfn�1a/#��!�?$�6I�M���mrt`��t��g@�6t��|b��s�d,d�e�ϻ�z*n�.wQB���n��s��L�#c���V��a�g��M	�:�Q`��o-��+��Q�&�y��Ŧ
�B�~�-�V��l%0��V�C�����7�U�ҫ�?}����P)�?�.A7{��K@��]+���>�	��O��>�����H�� ����X�A�*b��@��蒈俳��������bo�$"9N��c��"��*"�D�4�1��6�������US��=h��o"N���V���?��qg&��7�;����|!�v������� P\Ь
����FA���x2�������{���ͥK���S�e��t��^<-A"���̮wVb�.��	Ke��Qe.4�N!�$D�-Ԟ�����M�8?��s[��,�@k�/���E�޶[9��E~GOq3C̦O��!�Q�<�Nۜ���b�Ny�@����"G܉R���&H�F�z�0(T�ߐ�i�4�-���/V-�Gqp�_Ӌ��V�=�yw
��;�����V��h�}��h�����}Ysޔ�A��N�m�CE�wu��5@��Gـ�ɹbǬ�+i�#��G?#:�	�2?�$/P*ۢ)���$xhH�5.2�^���K  ޛ��j`�{T��fc6�s�b���d!�3aAF��R�6IG������n��=���Y��/�Y\j�6Y���[%�g����x��і�_����u�v:�]>�[�	�{"	Kx�G�'��Ȏx�6����>j��Vf�;e����i��T6��N����&��i�3J	9cu�1�݀|<H��/�w'�:����U�;b�)�W��6|x�s3��w��˺L!kouC���5�7\���
��5��O���%,����~���H�h��h�ݛ�2�IQ���6��@1a�7���6�B�.����Qr�py>o#
�B�^�͛~�i`�м;i۵��:��?:�ʌ�;Krݴ�C״.�f(w���.���!iB�v�h�7;P��UWG*P�T�_��m�E�#	�"�޴�6�HN�$$�\�'�[>Q��rkp��3:EF��?l�adロ���b���`1:�[�ȢϮD�s��/c�\Ʉ�� �r~&5�p����K�P���}�W�5	�>FP&�¦��m ��H0�
[�5W�ՈLTv��?���L0�����|�^�"G���x'�N :��`4s[A�����>������3;+M���I<aęъ�K��8V_<S�Tg�:4�+�0x���ɺ���s0$T�R�*4o8f86�h�ȩ��м��'��!�l\�N�krZ7L����M��v�z�5h�2o��m��p�J�� �2���V")	�&<i��u��G%&�3��;��ؙ��14Q� f�����k��+�#(H�'������0���� �FYl��hw�2�i�"�*�d�0V��8Z���CW~�w
����n��"����݊i���J�1,����N�:�~ڻp'��⳧;%;���*`����R�
�}�ܭ�%�M�W���6G���l����α��)M/�}.�VXwF�d���F������l�{H+�7��5�=�g,��Q���yY�����g����\g�P��8�������.$>���Y�";�Co�����2��՝px�3�,t�J6֜�U�9������Z�|�:LM�w��!M-�$���a^r�i�mt�@����}ݩ�^ͫ�7�~Ww�T������E!d��,��7m�9�oΦ��X'c��~��}.O2VD(l���\��xPm���l0 g�N+����4M�`�)t��ۭ��t���K ޽���Ax>��@{�G#�F�QD����"F�w��m�I7l��O%�n�%~~Y`�ң����K�0�tJ^4�*�i���
��Z$ ������d���Y-�as�p/���(�%=�w?���g�}HD<t��hw��%��mh�|uYޣ*Il�Ee�';�4�X�����LYnz�X��a��B����aL��U�
k�r��)�~�a^16W����0�;�j�D���Ջ����6ü̱/��-��	�Ko,��:�~���{RD+�";�|�@��{Y?�j�_z�QFd��rt]�别��\y��vW�A��j����G�έ��ٝi�iߑT6];��T��*�DEd�{����>��M=�&d1p���)QN<���~�B`O��j�S'c�":���ȅ�!���v�;�UWXv��Oe8�!x�-�F������ER�_�)p�^�xۺ ���<#n�7���4�V��O�g��0;ܨ04"ئŨ������4���%�#~t"���)l���&�o@�j �r�IV$pPaϋ�tµ#>$`ʱ|`jOvG��_F!���0�l���|�1�~;Y)����ć�%sQ�P����f��(�~!>1�O���>�{i)|-i�#�Y�A�p� /�)"դu�s�����p�[ώ�Rp"m׾��
yJğ���r�4�F����:���?������({��iޏ��)ڒ��o�S;��I6�P�&����-P�ʰJ�W�*��0/�TO�}�HT#��u!;��N9!(����rw�F��(~��*2�}"m�4�Й�.@A�e�P��Ӊ�hڰ	��>U��]�����j� ���o��K+����Ylt�����
9�یK���r�fT(s"/�a�쮠��N������g���9^��|..�KPR���Q�g/4PdI�]q���->��m�i��#���zQ�L��ak;��GJ6��.|J0ƻt�z�@����٣�?�;C~Tvn00�7r2�h#�l��?}x$Ş,�o(Xǃg�v/C�S�
�~Nf 1B����E�$2�Ϫ��R�X����ˉ仮�(�bG����uQ���)KMZ����řd~1�ϕƋB�vQ�`���є�צ~͵M�L�6]a�S�x����m�_?S4	D� v��3@aUw?��4�j�g񸙞�wm��f����l�]+%�_& Z�Ɖ���J���Ük�4I$�U��ɺf,�k��P�F*�WKT\�Ϥ�p���:+m�_y�W�=`2��hKت�f_�����9'u�9 ��)�	��1a���]]���p���$L��C��N���>).��^p���I��k�r��r� "9\����A5�.�Ky�g�z�Z��w&��f���������iy��i���2��u��GtU�w�/�/��:9���1y���F2�PQ??Ί�n��M$[���K�q�����4
��,�T����lY��o��⟓1��7��B��ַI��-q��s�77|@�IEv�꘻f9�P��T�b��8�V���n�������\RV���U �z��Y���n|.�H)����`d������xJ���