`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RbDDDJXosE1MH9k9SrACWqen+JHJgvffijY8aoyuhutnyQlfHHsRyiJK8y+U8774
CwsunxM5598+eRtrmw9uWCGwUsLJLGL4BFVD2QRB6cm7bT8FpzY980gy/E6dzaB+
bn0Cx8gyF6zhvG4m8WUWgyiBbII/j6eSL3I+2zGNQ1k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50800)
ZctGPsrtD/BOBeSv2+DKchto60SRgjsEAqJkLH7vDkn8GxtKe/o0WbRg54ND4Md3
wFRjWWJCqXg5KEb/B1Ex2A1Rp18t5wFz6oXjyd/tP4UMfLTRk8mApEI8v/irsTjV
2DwKUWIAQR7GOTo7XrMorWMEAMZ1ch4Azo0gEMUebJ7f3MtBkvJJFWSqmlwQQ8//
amsFDwiIfdnNsV76ZDZNcQnYgKTru0FaAeUke7IhGJiYHR00tU6bhZEgxWnL3Ec2
xKg5SAU7ObPD/L7k0G+rznFGVPEzOYIwSRMrnGKd9hwDlQJB2iMt9Sgn5QyspP0c
/K1WcywlXdlGnepSAaVd+bqMDtL3T5kacMeSn3/VWVnzRs6E+BT69Nv5vthdn7jc
XPfYvKFsxL4+p8YD79wAGt8F9O8U0VwrQbCgoui6Br1TzKDRTIvHcHJNhb6c6QZS
haKohXx55qqIsI5UWkH8mDwCBz9kcVsNs1ycS6cHgL2GjVt+3ORNy3E/j3pnPAWl
Ny/ARyW0487YLl+KVwFh1K2B8EaU8tEB74a0cr4mYRc3uWepuVLOlPPLdrmSpmsn
lxPNTO9fLQ+EVjuJHXoXZQ3NWAVysxABuBaTjHokscI2TqvDQMwCe+Fkaee7c/a8
NXAfSRTjk9bIBeMJwoUGE+s7KdVaWs1cY+wNj1ns1/F/BWrtBU0LZrKIP3ZyQRWl
6l++fhmskK626uGLSxTCzWvBWbxJo1yXUiuAiVOF4RiMEm3NPa1ZtDN9IuOHsZ+A
5XVAzPhW+IcNeghLn64zF8wNzEEfMAnuPAP6lQtNWc4FGVr0v6iDWZ3pAeGBf0QY
bAexTzBET6qDqnWCEUPmmi0ln/H+DW8Lvr5n5QzZs2EkDYGo6zT3jsZGFgjW5s89
riQQ4M8tkgCCaMwVy3bOaQoT3aQ/QuY+HY/TH4YRGHYDy5/z+9eMxlDtzj3HYOKX
CliA9CvJBwF1/TyqWaYVx2NN71yWLriUSNSOfi8g1jMDFAKtGsfvQox9IoY3kxH9
ggWwEGaN0ojlgjUPoexAq4EwrHZ6CmQnrWFM+t8ytNxiTF37mbe8PS3RZdmU8zkL
FmmDTtXOCZ0CpSms1THKCNp9ENsZcGLDPTYew4G12R9f6ZAZQ/UUGBDQ8UflLbed
TpNq2/OBpM7TgYTNB9VPPy8z+NvNcfAaEt/7xCq6CVJrryvKKiCiU0kKXfJ/xGvm
MoU4fBBaxrmukL146b35aPF5JfY5sqnPnupXdkDJ6XsUlFx3SQUje8zYPt60aezD
Mh0oIPfCy9v2+MjhhXx5NzamBoNc7C0KH66VMy8HAyxUwN1oahlCL4+bEMM4ewW+
DydsRti+mvd4rT41tKXlxqwPXFksmQifc9JB6bWiGk0UT1IQr4Vki8ctO0S7kdSV
BvCXaTwiIcDBxu09m565shLQf6DaguqB5aiIEXYDWWCmVstcJh8bP3PwRBSdgIMm
lXIScc7/J6g6y0ifzUg1qJlkySDTAAEWq4yBXKzdQRzEpC2wT2zR8+dY83ZIDeOz
o/tYPcRmjj9vgPSPzLv1W79PkKCyYFfX4T4AMYewo3+xYdyUOM1EgELefcTb2aeM
Dh/B96RP2htJ1aycyFH5XM7H2vT4lVcVNBYLmszBZeiFVYmDYb2YNp9O79qpfWpM
I1YP/blW3R+ePrYwqOSkpI3m3zz8tfvBhNtgdb+fF722v05jiHIS/cF60mNJiXcK
UdveqJMWKcFGfV20vw2i23fusXErLE3PxIDqfg9fWWAhwnIhz3QBomzldOnOMtKC
FxB4VR6ROoewwd9n9zLNXKGwTJnkTtiHx5CBDlhC+XtfMDMUrFeRPvQCcXu9NgYh
2lbx5zIPl/cFN/Gjr63RtLe+WQCWNTBsJYh9ckYjhuoLnwufFv5t1gXvqAHFlWyh
mpo80O+ddKV+C+QW52J6xVIbqudDpQ9AKapHk14TtmutJc9ArUlPsDo8dfZUtSOb
Ruhs0sNKRXsLCgXq1YNwMZBwmIDTxUggIuo1AT4jxxEhOFNqIl6QFfR0A/HU8Zxt
d5NMNtVeKUkiNJZqlLeAKcwP5SyNzSaJHhB8SO9OhnPxvqGP4ssoh6EjzOgx1W3T
pZjfsnjUMfDADr45GjC89dhBn7XoB7ay+1HJmmLomE2+xZy57k4CCepuJGM3W8jX
8FXmfE0ATdWK9Ftzk2upf4xlI27YviC/8fd0Bqe3SanyYLQgfGHzux2Fzwfp22rV
TGnxsjK3oomC5eVORmjcF1u16MWliF8qCx4ZVvfnc9b9MXHaQJck/LVV8QR4ySpf
TI7VLKJ4SnHjnK+Mu6ifaC7uOM9tACTLH9dmVhpgTFzmXP4XjmIto2QmBh5nhF17
ZpCz3XX5da/ORLH0DeAVn6Xzer5eduHTyuZ3GXR6WZ5KjqH0+MVDcla9lcS4LmxA
dqelr/WfQZqdLc2dYAUCDNk3mLHVgvJ9fxrouLm0g6Ih7CrNsCffeBVxMwWAgBht
DhshnvQSg3zGs44VB9Q+FN/d9ghF6GnAvGFQjS7LyueonWrIu7Mi973wzvUCIuDt
pE6Mq2xyqzI1+gJD+7dOYILrNZ87LfRq7HozaGLeyE1itngZx5BL5SDZ3ZzpUtcm
wOOH6Flpl0Hg5GFCU+nBYX4u2u76BCu5YFl0zVWE+qAn4DEhrCy/RNL+b6pzUecB
ffGhJ3tHcpJPUP5CwiFWNkQnp8wVnVxTPV5xa1JCK1lXmzj1TDPNUkzgSVZdtic4
12guRQxAuFLr1Mf1r+h6teoHRRz0oqxMyxOzOAVl7yYaAGU12IdH6WiWscPJbMiN
janFnu4l8rR2w1ZRVVauEQEmXJ7Dd6ZoA7TQHYosOLjpOeD1egS7nSHepVx4KE4R
mdqpsZjFA0KQc+tYqAboxyFDuA6eETE7O0eAi+inS8lWghBqN9uUnx4VW9PGuKHw
fTxvLnJitMA4n+ufgjW8ihyFPJPmgExSPJ8DVkdjaTf/GrUV4EDRv22wj0F6/Yhf
i2urRd8UU4eVHis1Zgg+w0YWKXbLpJe0+OQJIZm94R+L22QqZQGHwQeHoHJo1jAG
WRtOEvYxqXdHdFLnNCitTT5fhVu5CHePFcvnENXSyKXgkZZkCenMtBYsItxhbFOR
K3Bc1MoVjlw2dU6tGcH1kHO4AAzojatLnwT6nNHgRKjXoB2yecLTPuBcxKqLk2Ew
0MlWPbs3DJdnMO2kzwr4K78WojmtSyLYNv/4CQd6J3KrXJin0wQGUPTo3ikDlmEi
3Qody97DOlcm7Nk3n66I7PfT/P5GjGFLs7AeAI1s1b61dE6BheibMwRHVzNYWa2F
f2nDeFUB63oMEQLLgC5Xa7u058oLkqMyTrSXTpgDHcqYZreHFveTKvcz2N/T85G2
oWktN9R66SsoBaysVljlq+Cm9gClykFLzK60ktALjHS/1QZprJa1ufE6kgMoRUKT
bv9hAz9RBm34CYVAGZOd/Xc4PRCOSF+XyuLiM7yjIcLXIOfZbQmZ7GHOS56EvESM
MO/pMAqAI/oAM6XGxklPYnZNdmdWORHPe1f9YGBNYebOu1tUiIWCxhRpFcmpw7vW
RTn6z/6/nSFMPHhwgFmP9Rgf2PCQGlLckP/I4t2JEsrZbal37doL/Lf0V+B3eCVE
IRSkYolSQ4q/a5RlpXyeLjnb7ZSrvKzEQCB58Hk92rFH0UGM3jp6OSIjtVJSQ5Xg
HY9OCGUFMxZTHC9juIMNYKtJJaon4XLFQ2bjBxlNIYht+ZwLp+ZuIsMyeJbTXSG3
dov0rZM64Kj46a3xsJ2tF0t8RZ7iU3nAyAn6dXhYpbqjMHdv1Ba74Xckc8yVbU2x
ydt2Xs87hTjvqQTMru12S9IoBfg78ce1u4oAI3tn2qyhsm0kw8ucJ9LcXsFXlXba
h45SkISaxQ/ug86A2vWyQQmNSt3b+CDzXR0cOH1WbM/kTONxJvHSEGdmBQy0Pd5u
bq4Wb+9HRnbaicOds+ddvNXUSYq4Ym5kmyheiKp17BF30nPw+PQl2m/unENWfsgU
wWSxpnniNAJpa1afLoWzTY170J5chBs8/CFWyG1cgY8tD00jqH9COfn+SJTTZolI
blbLgft8HNVA2yyJx5Rt1YdbYackUev0N2AzMHMEI1cytlj3oidJSACn5n6muFYA
Shpuet7XIFBqZnlgOfhydhSUv/qVzMdQoIeyeF3Wkxt3Tpne5Z0IXfuc40jAHJyc
MSTaHvWD6H4FUXV6C8NaNy9LQDhWRctDpN4H1joCg1ymFRgoC1K7B6iRUESFMQsC
f2sI6eQIxKolzCatrcdw38SV5Xdvt2+54FoLLPiv6wij6AHg3V7DImEQU13AYfw3
gc55hblHVQ0FmtAQEBIf1fYDuc3cPAvM9zHH2k8TYmb/RvAkl5qT2tQQE5ykMLSq
PfEcXpOeUl3+Lto2SYQu7uNqX39I4fnwao7mwAqWH8LJ06nUn6O2xswKKO8dy64z
DrTyCy4N8p/ZyxDAMUNKADL1UIBl/EaUhOIk2FMBg82aB0OnOIGZH3ALTLmoZsUs
OwQewJKGzCuIyro1RwPO988OYugXtPcqiNMiYDZ3GnaldKiuurbuXWQUM49NCsez
p4piE3xPfWfgHcH0iTPCgNu9N+JHMYvtRHr5ffmxf8volbZqMdINc5DSZtnv6fPS
fi4auEwgtLApU/gL++9H5QCoFvtcBIJi2FpjrhT/ngnys6i6bPE7lz0qlBS9BfP8
6TtZd5X26UTCvtvR0ZB1zT+/1IY5h7+ggz8Xf54sppSp1Qe/dBCRuRY3bKmH0EG8
p67YRXzfORv57WEPoKM4CQ+td//yjh1+mJgrMPszUwuxZ9/w9ET1qHfmpo4Vcgsh
fzKz2sD6StMPsd4GD5kHQzG5fxLij0jCM0bX2g3oZveVML0Lyzlcfy+hSKsouKbP
SMT0G0szgnJvPLwhBjGmr7VeKlXeMMmjLb8HuVRCGQfmk4/zZ3Y3T0wGfD6a1bNq
RCT2ZboXIFxnema6N+v0YxLIBAzWfZ61aG6GU/HGrI6l4Fg3DfUExDYJ3GN57gv8
DaMysjtX8hmcPyh+T9tjnRfUN4w0tGe/qKDAV1VZer+u0ppj5GFfESSgpEnhkgwp
D0g4YPrv7X8GyC+qLAw9DOo8pB+Z438y2rbQFWjowdHBsdJTPmKujSHiQ8lu8cfe
lbaC2lJlxH6FHKMe0D9cCyoMO/SnOZEXnfj4N+8LCm/ADtX1If3ay006QO/oMJIo
PMoXRcxNn2pOegg8y/8HHLp/4iVII11Zy7EqWq5x4fhGUHyTeSyvmPA6qpCn/Eux
7p3wuuXEhK/Ea0nb7GPkj20DV1xFPMUH/6zAY4F9e7cF8jv0Jlg/LcTMXOdZMi1I
qjEFVrGX5j4D1vcM3GSC8wCLgywbt3rz/fYWnMTsSvERZVTUOJS0avv+HgHwH8dA
KeOU8bonv8lb8I9N6TvZHQgP4uUzVX/md2QrDnOsLcWkPr6NpGLmm3b/Qv1UNT5q
S2CWWM7ozlcopP2l4DGvEFYGOqthoVrNmW7M1M4TLCIXbbd78vy2QUfg0mhYtocX
or+1Obk2n44s28YwdF1gEUaJ/oJRG6r0hIvdSaJ/3Vd8xC5gXlB9OM/jvPeyjb5a
F+YLrb6UCESLvFJK2o4mCWCjsgIUU0BLVECkXWsCKlUjBqiUlWbue0lZWEmKGHhs
WUS8oaIcqjQWQvWbkf6DQJ9hsXTCqbu1jQgzy+meiT1gixjlIStX36g8U+WD64bh
IDjq4uLmnCh9uekPO+mGRBLg3MHgIeP79ckoL4OIzr3aphJof0ciw2lMc2VdDGLw
V6Ypf1nE9XRVBYA5yCV6Fx2D53ZIIp1PDPPzLDcSw7Kmj/UpelrthGHbwgnExX67
GsSskGo9GO3m5JTRpfe2wyZy/8dvLHzP/ckgYLqi4BbDVyjTfkSowG/90F52iyQX
RD8ckgEZ+kUEM8OJgsZvwGsGvN2Bj2T8J2ELvrAOaLy9/bjFuIERgYvKSUS26zm9
qdw653OYRB7Xp3ldDp7x+jUmA+aoR98/jMy7RzFoAgTfOccxAXRjs/JOmczInT8O
6PRocJ72VMElvC8dpsPii7eEvDqwVu8zvS7OVECNmuq1gp0DhkuJBoQGdqT1C3wY
ncpJe0/tWyN0qmfJDX+DbRc3NWEX3YsKAqzwfo6zcqLlrgt97qil67xn3rIAy0to
ZACYxUlJSIqR1cz/JmU7DslIkJ5ALov03fbUx4trqZQr2gmsJhKlwcC3mlNk5cW/
MTZ4XEjBSRrYMho59a1JcgJBADolHZi9leHLrfZe8z4Hgh0JBAg5bMFuXhsLGQDa
HBS8OHFKaYjHCX0Qo4oiRPmQPHSMg32yzgTjMYiUUMQEd8PvnEzL4GWD20hsfZVe
R++ohWX/VH4i1Qwef9Np0MWTyyGDcvQ7Zbt+uWaGSm9XNjV8jWt2odPiMF/HP+IH
4xRadTCkctL7FWH5dSkv+33eZPEkazm1dDG9r447xTPS5EmnsJTLsaG29qZ1wEVq
1jkGH/nzx8mwaJ7VLshF5KDEvwF/thteJjC6zLRLRRBeq9Rr9B/SQBZ/PP7gKCsn
ityGyG6dipnUxYBhb4ZTlfCtrMChcrFzsNWa9zpQQj99yE9CmVKYCnUjCAdj7f9v
XI3CdFR/XUJ9fYaTlQFRvuYtSZQ72LVnkZ1rudyv40MKviJ3OtvJ3P7sVO7uDV/C
dQfDFei7uSOjx0WP96kH3iKV+Tnr0km7lDzgMvHz6b6ElONhmkn07Ba1XvtLi/lw
fTa9QsRmqFGzEAeDZmw9KmNxkN+QjlLb3SmlSfF15pbu0xW8gaeMjDEfVGjv6ten
c7ksvOz10xjHWLSOOokOT5g7GDpbHoJNmM7Tkluoy/6/Oij7m07r5jfjpwG5/XTb
M1VZJUfDTBfFEhpj2OF3EwMIEu9KD8xFCQnb+uIyk9J1XowwpBnAmto8j/YVDTTi
hmk8IfNIWiIND29YKFdRs4A8u6V1sF7LH5L2Fhe/7C9jLdkLXTzXR33eV0DN+JYv
+ZoFBy1SBuyhAjmRRl8f6STBeJsSzYPYnBLAROb8kcKoj74BDL+y0lWstXf6z8lJ
xqcRsLVmXm+DRkcrL7jgyLc9HbB0r4YoPDG0C1e1lavfTvHaZjkPzHnBS6WlBJCl
Eah1Zf18JEUzi6jFE1tBsOMRJYeHrT19Ict5x/jz79CIdfTmcb9OIyHetGTQu9g5
TUe0ho6WsbKB5jXSMl1M5Wg/sZZ7lgURB6w+O4mCY4DM8RBiKcZT8EliW+XFEH8K
rto+BhFitwrG88Y7ErMm2CCyUs0zhdH8quEN9DqFG3bac2LQ7GjU05ZOt4R9IemO
QwidnFuF7XoUWi+EDsxsVoIPQxBkP4QIzcfLtxQo80KoToP/GDRG4LgOWU6yWKLE
2VaEjBZEX7HVRdAs+3Zy7KDlHRoZtiVIT800gu5VUL5ITnr+Dw9mEAcH04F3vEaz
dYZvzcnilsUSKO0O6y4wXLcrK+H6G4NV+0lmUEW/bhE/zPDffMkaHgLYf1wIfSEO
sz4FI21kxU2dfjJtsOBGtaux2Q5xW/qQwbg/2H0hdPZV2uWZcxTLATEwiIXGyQpG
2SVmu7ysj+dAYec2v4T9iENgr8UlPsLSlg/OVTNNklg+0dmCBruXcOc0cUVussK8
SgHoZT56UCdV81CTlUmHBU5eNHfDYAYIdLr/+gs0CijY0wi0FQjmCarNbbKSGG+Y
2ouZnzLhnGP1HhSt03OXWd/2LER5wUFmIYUcwZOOQdzZIUxvH8D6obw6AUaphGOw
0LZFalIesWdJf9i/xu3725af2Ho11X8r8DzaOBy7SRaMnVdMJ9y4ipsYxmO4wp73
1/rrdNvgrhKylLL9y1XU1hQpogvoaozJ39Bq5XzO1fdG+tNvkjHA9LMcU+Ewheog
cuJKEQsRIwC00yx7Sf5nyuSfI1XsUYHUc4XEVQ9YN1zC/xulkTzgrmhHy+EkfPy+
j3JAnTyfmJMUrNT0tbBLdc0p9wGw6GBYsQADh/mcGZ90T/LCdAcq75O41/fdvvyy
Cvk/+Y3zq6yP2S/lktZqCTHSoYiyT3QkZ15PzQbsgGFdvErS26G4v+XYtRJWc0pC
oB+sv9l568Dh0sr13hyB9BRWG6ZtuG0VYqPUAEUT1pFLKUKke5PWS6DkXaP8PRyO
rmgmDaPM/j5OOFwOQ3cEo6h+SRda10AAkVknwXoAoU5VMwpeuv86Ieyyz0Eg2VnC
PcpVyyUQSit+DCrtCfjoxG0/jmlVce0wcuGMPaBlzk/qDOp4J/uBQYi/sEGdpGkw
uo4v/zWuTPXC6Lu2OEQ4C4HudwbVFilkzyRHnheLHeV9heiowEp7vRFhr0LK3WzR
vkdgnE86syHfszowiKKnUM5n3KtRgqTjQb78osNLjFzsXiWPBevL3ikQg4LnQ4uD
T1N9HDJan0/viY0w4BhrXPGkz8toncgwqyyuz54FWnGYjXPtzG7pYA86wSfcyMgo
Nr5eKV2xn+DQ2rSoOGpMPf+k8YmsBpoh9s/WFLlLdH9NvrtrZPTNOLIByGct+BcJ
lBRvRQQyEAg25IMtlQAnTEHyXT6OLXmfj6WDpqvZa7lZ4Ruxlp6fy/9vELU8f2OL
RfvgPCv/Nwb0SEGURaEpE2wgLap0oCR1rfGD0zrSSZIiOSZnu9F7NB2LujvzN7LF
mAZDIWrH68pBuynr6+lN/1xPYg8IWDHCqlwL1kQTww5Q8nmOsScZ4pcBfId9/29T
PDJ4zN3JpD3rFaHyL//1S4sXgRyfbmxlMnjx1KKgR4ADSMqhh5vS6hRWm/P9cfMo
TIsKLoiUM7SmxCSY3CP8iVO/dJy6UF/ZIbeN0myDp7VoCGYBWRMlMJ7Lgfl3MIzJ
BnxG7nAEva22o/LYQsFBfvkTeC3AR2YiW7yH8f+TZakMhjAvU+K0k0MvOndcXoGU
T195PLJ00bVfQ/g4F1PlfuqVkkBBN0Yunvqmo1qX2XQtw6RijYdwI+XTuLaNmVmC
CibHZkiBdsWo24VcmbWcm2ZkHqW3uqarLwEUC2KJvqzNbI2uVRKQ4Cus2JWOwqly
RlwPi9IwHsV7lLstYE280bxy4NvEY/pS2gVFQs9VzZUL8yTJUYp73YIB3ZWD3wID
aE9Zs6zunDv/MI1WxlFlArSrjhwmHq3EI8VWZQ4Yj9mHqh9ByH/e+p2zIp7EPRWo
T/FJDKPocr20+vx5wJOGLOzQ2mMq/WcTLpt4zp0jwE7WX4hhHmMlWyU34insJtEL
B+Op+3XO3Oc1puhJ6Gt/vvf4pe0apzuplDwmHu+tik3GYA5nEH6uAGAB44lsNmey
0NwSdJnEw9EYfHVWCRdrKrZRkizY4LLV5mIE+YVu4hQ1nl7uBrB7KQEZotiQlM8v
DCwnmnSIK4aMB9sGmFq7eGvkpAvsokQvmuJ6tzTh2B0M58rPuv19e+gmvGxrWjIz
iz/jdSpKMaJQc/sFsGoD+hW3KaInNEjVg8Jih6j5Gr5sPV5p/mchenCAclL3KAFx
RtijujF5Nr2Vwyf1yd1KfjdnrifCyqDh5A6jdqaibaAovQoxsjum1JyQ5aTzJocO
WnAZHLbR9vgVwrpvoxt3RUqrkr6qYnR6lO7FpSaVioL4GxhfZ41fOpyIhwTHyOfC
UdTcdboeNgjbdVSRYp9XuSSCuaUeSwUkiKgMKSX4CAihfXGzjJ21YmsheNS3Le07
cdIndEyAuiZ7cgcbSFr3WstRQwBDY/FcUZT4eoTDA1rRHbNOfAkWQKoQ0cWpwjGI
rqe6v5M1auEKyW1lyt5fhrU+x03Cm39/qZZ7CrzrbhDdlMy4PH9aig6FIfxUcTZr
/F7yn2vfQVMTpJMsW78Ye2Q6bujeUL7fZQntkw9+FPC3tyVZruUP1SFJcMwX3n84
hawcxkr6X5vi5+L0LQBYn/LNU4DlO4ViZWKxJcLAKJa0YmlKFBIpxVdBQcVWvXKi
mkXVol72VndNWzKPccWW+7TI6khPICZ3TZJ+Q7QB52GwN9g3updGKFk967AxFvZw
qn+im9+74QCtRe3IX38oTGbjKhiyIB71EeAwEYHynyVcOAXPQHTXHxBPZ2Z/tEJo
evVF47h3zhA7daCGUGgSwEGA/cs55pAy5DNjQ1LjgbNj/0yMQimEN1cADgBxo4Qk
jED7ZVOp0FMPOVc5yRX5cJlnRiYZ32QjRAwahFVZQ+Ycd3HsoHt/+WFAi1X2F68j
ruMJTlG02eG6DOJSp/YV6X0HU5Q2MMk7ETe0hUqmdxiH7Chm8KcnYY4JjCOxpzq1
2G69HrdcPPmiu4zcGOna9u9iQrlTZw/ALYr2Me361zStfL3NG615lH0hp0FbXUK6
zPUGTFk++8nOmp9RoO3S0KVgRTVROQ/b6x3bcj4K41VqfMdJJZkjr+vM+eiExeE6
etXotqQm3DF9BQKB2TYAy0M8dE9I1Fe+JlTF3B8dPywO6Zqw8TUdBAx1kEgH8Wgw
MunzZEk4T/PPqXm4COUb9zPvvwUN+pDSV6BUIbHaCtrhXeieOAhRRW0620uq0RSU
L0NpzhlJENecR2XKqj3k8+xn5Fc+0+zqaguJ1aL2TGrXTyxeTDWVk61RYivzKLkQ
qRO69/mKuCCxHO+dLWKb2jJ0v2Y9xwrFaHprHablBXGZG0+hreJJqFXaHf6+zTnn
VjrrwoE0G67nojydpeg6tNMrbZOBLlPIRvYMMfBhUBpQGhbrMKufu1tBuefs5Mw4
r9GHQD/VPZhXMgnz9Qxii3AH9Tl4poCZ0p3RxfkVUa4YdXGL3m5Tq8rtiaVVMBUE
xhN5ZNF94FWW5sh/IAdUmSFPDYk1ClGORlX8t6NcXoRpOi8TivplLrRH2sTnkQFE
aDpN8d2ukaX6poxq4lXFkuSIiBpBYqd/sQnawC1CWT6sch0Xofhq6rTCShUCsfUC
kDe0bV1qhs2ONBYakcGHy2JxN6JSNQJ1i5zJUt7Q9tqzr3WJVEBLUbl6pZogKWG8
oUHVmSFNtiW/KZpkPvzV1DWzZAZKZ0oCYLudCWPBkWAZKuzECNXdvt5LtIMCnOU6
r8SXp3PZ1zek79m2eSTFiV5HHw6kS/Tf9SyAekcNVYpDNAxwaMKORUN9ad8O8CBp
9YINZEuJBvcIs+0hTZgNCYIFyE3duNDGX2u4hD68uqPqKUspb2Li+IQR5XeQfha9
FtAiaAIPlLUyKzpUa1wSCp4p3FEOI/7fc53n+xCgSDqoyrgA5ixoxxUG4c0y9x1w
h9Tuwla/Tv7jvLNUsGF/d5a4JxhijkQFcIPUhAAYAl3kRUtJGWsTX1toFEzvTuhv
GRDVoqrj7zlmer+kaTT9XxXV+kEI8QUVX7nnA6sQWDJHCSlzBXOABidwtOU1uM59
2aopaIQAP2Hi5p9sJwEZo5nzbc+CA14uOGCD2UGBuHRB9g6jPQMhFPCEUnPCW58F
b2qyvmdvKuPgzMBpsM1VdeM8hVbShlwv+soZwII/37tvouZaMXlxq+ALjjPwiMM4
kiUg8AKs3zTeJc+kc6ob242OA3MmBXxdIolm7hXTJcxAh7ZO8cUo4x+ZYvPHBZCV
gYnO5dQm8KD03yYHvurxUDBy73KW3uycXNiKqaJp1LJnuEhlXsjRl3irSQmoIghc
Z0FI9RK29fPy9kla+W4Fsg8dhw7xTcNj77W+dro3LIdPFGtBBfMMi89RObZqpXH0
6D6/xOLbPVZc2iX/1XELkR8tWNpvBae/684kgwxv7MthHJHWgf47V7f0nEk4cZ8s
yFSuW12uqLZU2X4aDyPsdMO7XdyxaEpIawooCmqG3f2PU90mGSVp06FIOmAmXFFZ
g8qitW4CNabe2rKayta2/vpUWRfqTTh/Odud1MErH5aKyC/L5rDPSKfEgsLYhcM3
zt3sxKuDZGn+gPL1QpFNWYhzt4ag56JrlNbjNXQxOXRTXZJgPbZ3pvdCMbnnPvWR
OVltfoUKYFGUUyVXwGN7GRtQaf7Y/f7ikEhfxzgdnuE4U2aii/XI0OaAPcBqbKH8
oGb/eSV7e7e27bhz1gaQ8sAaFdX7NNEH/0x75beY/J/FusFtKeUxSfAQm2QyWvwu
TE70Tucmq5NFGtFH79uOGdMyXEdBiw+lqutFbXHXzdWWIY5d+umKxgs4HkjEi3rb
b4DmpsY+X2Qq4EUPutw0TF8Zt6wH7xCPMzcXu4gNU+/f6yUapVpNTwB4U5xbfM8Z
cTHe1+6w7RoqLOVoQeZ3n7Iw/lTPSJmlEfGEUnXLmbZOEF+R15xxFY+7Ogq5/Il9
USql7BYcUXo3p8dAK17SvXBup25r4JEFhKgRVyTXK6XS2VdAagRickLX9q9ErF+U
8Wbh0QlqMkoK328jwUJHwH3q0HHLxt5kv/P1GNLfNgZaTHNK5lPW319K+kYtP/+z
lRutzXovQImuRaLqa4LfDVg3BemEz/J43MD6ixYEf/vAPQmeaC2LBg8ERL3rWgde
6e6AJNHpJeLfUdms6cegQXSraMgw6oxK+vLOyASXO0ib1KZlHzrkq3QFjNb5Nt5y
xT5TdC88x51kNvQg/vdlRUr72cPeMgXr5Rtn6Ukq62bysSnnXqMNbZjPOAXeH54u
nGSdckzRxro+jFT2LTTtke7bA5qNlR3bhnZ9tpQCXevnYku5ejsBLhTDhyJtZQdJ
CwphAjJYCuWCl8IuquWhdyJORXMGP9RUjJnaaqIrX/VKdCsop7ZVQgjMxIWUYOOQ
lZoXGXxtk4Nnx1l/VevQlO/f1UBG3tKsC0UFS1xnECTGYHwlyRohHLGsXEUp9Tw4
qfP8P4mbb3Wg2I/PwsF4rKSOcRuX1nm/VkQStSAKCFUYw1QrU5XZkLAyaXw5c6x+
XNYky2/6H4773H1Wk+badaDFVa0D69tXrV1DHd4MuvIV5JAXho+4qt6X5SyX2kTE
LLbpw1s7XvXyslAKS8hUo75+4FbHPeMU86h3LxuYuw/0ydw9GygSiryPbWz4gjcy
ceP0KHQorXgPAWWJM4QaxGWm9JlqB0tu77qsG/H2xbYrCxoyzK9c8VHsuNFUVHSM
EKnMV7om872CYkf2ESG6NdsILGOsbiceLCBiuytoluM3AkcUDgTt/rBtD47cojhf
tFf5rmDDOw+70y2Gf6F9L3R3RMdCWKxwCdjzs3zWYFmgdK7kVbjo/mkRztzkhqOY
aWT//oTSWqbIUGJCpM59PSTk6vElIwTVWzr6mGJbgJzntIG7GvjzILXHoCtAxi8N
wrI+QTk6GR4mwxULzB4zbg/n/IFPS74yMK+ZnTKjLmQXE/xIEepZ16eMSgBQVpH2
0XUENtISkp0yKaJgYxo4Vv8f/ZrUtRBiWKHqITC0ZktBi3BWDeXVoPDEljZdrrGQ
eEThdmVqeds25avgkcumLfwuIO7s32+WbYXw5kumNEAsWdFKlTHD3bHcewXZfwgk
/VCzyyp5Lh2Z19TeCwtGwRMqxyvvOOSG0PeUKJN3Wy7y8NXshsEU0xhHf00qW9l8
QW1pUPC1ne8WE1lzy/yiYQGFRoOPnW1LRdxKW6TuGLlmT2SMX4ZzAsBzfgdmAzG3
LHEarNucQXz4WEGSZZ+bHWfniUMFmyWqnMs4XUCg/QjDwzg1oiI2M7g9CwUztGq7
AK0QaJ/p40PF9rbeuE6H9yklqcI4BZsm8oo1xLhWicfP2y0pHseNM4Lr3QADGoSE
0HOK2QyvffNVbtm2ZdEYG0+ekcv729Hk06EhKKZ93pyGkmANI+6t2DASc9FO/QJW
u19QVBTh53/UrZ1TaE5k93u1sgjVltphOX3IQQ+zlBpTIAzc5Rv/yBiAob/v1QsM
OjucJIzCIKVizhKXkz1vlKXGbpF6tTR9oEUKzCikAkkLEjQzq3tPP/TaPnLa44ds
fWB+sN/uEI8o3NLqPBvZFCOoth2c3qBHy1oeeIzgp7ZGBT/F3p2De2tkT4Vc3KPQ
X8kc0XOUboTwrgwKNS8hFhvqCVhBygY8CtWuKwkmzJEbMFs3AZYTykIWqZ5/tuka
GdUJJADxi1zDOI5a5shCv9FQD/C5mE+l46+7/iL/9bgPoqOJepy3jE7RRl4AmYAC
qwt+qpqqFR9T+hBWOMLyWNrhZpOTfO+OE1Bnl2kGT4pJAejE/Sj6Hc3tq9GGAr4/
QzRCKgLLwhH4KQKInZKRB6ANLsfaEZwOuunFSKU49+vnRUx+RyB6ZYAnjoMQNRvX
QHdSuPOPIn51sJXe31ajKJnw4MGiBF6UbRvbApegIL2Qss7sCmmv423iObZcTQLa
KCZpvI1oI+oqE0jOrVoWoeLaxXHO7QQOpMedKDbBAhdcbf0c2JEIzl/uF6OWewOz
Mv5xL2wRjvleNInkRzSmTFwiSqZ/pkOo5C7wcm/ZIqSaNf05PsMYqTi7zf0AZX20
5eamWQKIyM3Vdzo2Gp47p++hI83Vb4TBNQL5C9l7ofmc3sVlji1T9IDacE35xVaO
GSFGnMLEVYp2712AP+KFty4yGCM2YrruFoEFrpJr1SNAF8zAtMRFDeM3wBlULx/t
grXMseiF7wVIypeK0Xg6CuEFTncojvVUpoB5yS3OXzqUkm1gGevA4rIolGKePUwu
sMxSqY9jng1WBjaT8AfszQLYycv5aWko3O6YZe4o/IhgLFz6iAlGvdGYUqpU/jP3
rfy2cZkEB9dXVSbkTJt6ggai4i3I9orrK4L5wnYqkf7ovbmcjQeJcdcExEXxL0t4
NrYJlyu23TO0Q/kUaplDMBIN6haNAmQBffGjQi0vEFWEDT/SC0rW468ROnTUFkdn
/NnUdBvf93TG1zin6jeRVk064jtxew7Ne+n0MNZiXtqlY4N5okzNppIIOLdnD6Lr
WQSc5i+ssLK3NGXw0VHHDNTAZV/NgU/jdHvls6WT16kPbTVMineCHnQfhCghVFHE
m+vOk/lnOKj8oPKBPGeTIL5X/Y0TZTqAmeAtuwidJDsCrdA5T6nqLhEyojZQ1u2d
frRBnPIoonGI1HFg5KzQXnEz6HgVj56xHPtfIR87KMKXDOnIhb41nd2Tp3ZjnaHE
3N1xXYgqNKWT0W+OlWaamRTWPwb5NxJU9He9WB0tARJwa3jxRO7sAlcvwVBQwJ97
rMNN0Oz5i9U7RE6hoAFNijDEPEC6xDR979+5dPXqISADPj7qLCVYpo7c0Iz7pH/Y
Bf/lEngVKKJhDxFJvmzHk83HWNrNB+Y/Oc/4WEpF3KokDndXaef2UN9I4tiK8jA1
N/HV1FR44HbtSAPUN66WrEoRyJUYcm/Ypm/k+2xXouPPztqcaFBXguqp682sTKZB
Q+UkoItXtXYcdT5NFCNT+qta30yMseOH4Oku5J4a5f6huq3Zoo6e/rwm6P86vCD2
t/C/4JMiesMdYvH5SRVmZXZLK0b8PnX+eAyqRwxI4tk/1au/lXjMA6Cib3R8rb4w
HI6ER8mPTVMrG9xQJK8fzCJNwC6SI6aShrmP9MxBouYmyxHDKT0TlyQWOdR23RkV
iZQLaPGT9PtKNg3OwnLFKrdHYv4pBdNgOOqeWR/Gw/LpeIP69zBocaxkaj++oAeZ
7BEYXJeYfmzsCeXTN59bT/T3UQsCULmyfrJzGgWZm838fuYmy6LDXtfYlgzi0c9T
0n1Jx0LSY10qRnmucbWWd5Xgod85T8hzU0oqdJ32nbTk6ztFeWBVLPkbCCcsDZ1/
3ZsjkePrYCyEZ6QBT8oG3VashZ70DFutQmd1vxYk2ls4UDiBLqKXqjC7nS1Daw4w
S2hlNxqu33CMX7QgC52yRpYdZw73BHARLSZy7J/UfsRL9Hsj0tUw4tjwuU9m3RXG
H6KRRNAAu4A6tE/28vH8u62FoDx2p6GXyO8c5DM2JDDtPAPIb0vA3kTiZy+v1aIr
0gwszPdwb11WMeN9IZWLw4Ze8xy6bCj0yWsf9Hwn1j2KyuNj/Z9NeHeM6ecA2cTx
T6OF8vWg7abf5cx9sB6+OsdJ6xQt2hY5UKi0J2gBxtme4paFAGqL9Z8vlS0peanq
fwnv6+h1M9T3uS8DjeeoPIrNM93I/Sz4PK/QjpnY2xi5DVEDutfgCJuYZiqCQDnH
Hng4yzxrdzISsHgNCptnYCF79BemCwztquxD7CJxHjkIV35SRLhBvi3te482i2Nx
EPXD6rTuigOM25KiIHYae46ETitSJ02dz3suN6Ozf39jC2uVi0NnvfpYwp5CAA2l
f/JT4DZtLH2bW39+vMeHivzt2pueg/SzxwxRj16lZfIDIGRoaSTO+ksZ/86RiIKp
TfTkejYb+myaHdL3ILL/q429tTZDqAPDUdW+9T95dNsgP9JZAwhAirQZQEt2cxjh
Ji92Me4LJcTy43/00vqQaZJqj9Z2QytDaNg88dKtPxff9KZMtlGZ0l/8+A2Be3qt
oo3josJKV9Ob4eHIXOrV0GyCJ7l5W2S73rqPgA0xVSnckGdbu2cR4Fi8xn+ZnWrN
3RdLHt713bK8OEFJcOGAxnaWL6d56gYoByymjE1A0KGG/UA46hmOXw5rskGwF5kq
/gojX4b3oA04nJTbf5l+HdLGF0VaylsDesePn9WGe7wjmW1OeDR6OdjJUmaodN4Y
yY0J93FmswK+wPXkf83HDn28+n+v4IdhmeKwyWvONqgy6qzqCR/vRUUGGiKWzSNT
Sh422SWzx5jlFARpfC3/OowVyoXYZlvxhTfiklrGdO3hrAb9A9N1VwJryWE7AXid
PyyOmVzsfvrx8SW0s/TrTLYBRYtFLFOGnmPccBNDnEjhGlbs0RdcVJtUJiXSKtAa
ESCK4/67J+5oBJxBtsTYcfzBPHxNBlbhgSBA8p7Ruj+I9Mo+eCEx47mQHbqAE5cU
1+u/kT6+enCCBprT6uHjJ4MdwNwEmq0/hx6Ho4ms5VngWkFB4ZvC/1QKAz+i6Fq7
40BGJh67zXdQqmk2wqfQoKiyzQe0FDa1jAYr+uHoDRw6zupm4pmo+wyiGS9z31lq
PDEuQ3G6HEBuaysKBDjLnVDMIsGUaW/B2J7pl1FeYzpL8IchZfaLWvPhO1w4W5FV
PbUcpjcxL3kNVkP0X35mcSveGaPydax6M3/5yWoJ8WPWZkx8dPvB9+6YWASOYzbt
HUyIrJm7/c5ZsOX2GHeJ+FFUygeGD4/mc9P5Hjj4dv9Y3wR3PWsb5h6VBontTK9c
MvsYHL0jFK1uI/c/ff2Y3PfdQXdie38yBDFRWqnMYO48DFUjbrPs5BAgln1RCSPQ
rR6Zl6u67VtCaqcrcGwRSdZZ0EG5rvuFLKbonQYX7sc1uANiVj2LdefLkpiyR8Bq
6YAqz7+l7xKy9d4C8ZUN3TsNqWUSBBEZw0Vh7LVxm11zyKBpFyahv3JK0QpiR6Qb
Kl/JSEyISbOlZder7CoZM/ntJLR0DwSpQ5WyT9Gdlx4WJCl5F0vjd2pCvS60iYN/
JZ9UX39D5Inu2PHx4YdSOQy2SnwlnZoJoTl51aFRtHqBlV5yMjwRkJGpUayQkNw3
cylXkOEyAGZwTpzr0SpyhMhBIe4dn6p1mQgQwhv+4LYKAaZrItEz4Yaq7C+AHv56
l48i0IJLmlARvJnptc+0kap5eShVJt1mLAmNlNjt1rOrg/mQ2djC3MO5Jgrs3UcQ
S7XPrV0tztlCFgI2ZzpJyR9jGVwC7MyxERuFUf9f67gZpSAJKId5zW3dreWGCWws
AbtKCPo5qlgWdflvc0IPAx7qIBXTLNhtCn+wQyeLUsN/NBAaL/fAa4QbXOn3+NF7
VCirn0xhhtdSaL38Wq5Y5TfVTSn/KjvNHhbEaRF8h4ai2YrP5TUBMfJa3rekdKsq
dhXtBGm1MJrI37OD6ZhEjur8O09K3SYAy9MOuDjszINduzdLPZhTMU4A56fSpMjQ
QIDiyO3PXgnUSFeoady47OXwD4sHSYWftpltHNBP+Hlxg2gKCxXK1A55eDAYiwmh
qztpaC6lGueiDNOL08ac6ggLuKETzZicH8auOjqGokRs7E1Znhbj0QP75UwAFmcC
wEgemqwE+28WsExcv+vYllznVs1jlDn0nhH9aZyNOH68PHXxdgFFrIS76h/ahy74
fa7pbpsCfqNQ5jdgpAcT7WbrEOPTdqGpMZEj28HCgyRQ6bg4O5pK/lQgEhUGdUvz
Ico2yAAn9YFhAyilo3+4uqllzjhU9jPuefOlU+ShrUDVe9uyTxzpb29snhIH81/M
s9/b6JgbMFpTEpPLp+HQHSIJh9bBE24l7kbbcCFJE2dTKuLuo2cEPnaxizNUQ8DE
Ls8P10VoH5fWCfWA6LA4vbj8MqIHZnPyTCYnCmjoJ0fGoGPZhjHtYfF0vpJoaWVT
eboDnEytN5EkyuspGgmGympgRVIJgsedCmCUudkoPVULj0iloJfV8j2HwM4wkNAC
tMVka95wbXrPqx/kHRnMZVJRkDK0ZeOdK4qslUGrV9EyIX0J/C7MnqmE+WTddYBa
+T8a5MTULVu9loYoLCNYsX5SvesAH2yZP9MOiD8Tx1huQGaKL1xXv4VLTDIrzgYv
XzAfaYldwrTEN7t2D5Z3dgzrsqFuWcYRbgEZixDHG6RYjrVI/moGX0D0YnXVmIiR
1y8tW7YvoN2xbbKh0VyrmnkdmeH0LZyGn5QqKMSHBehzG7/epLhOAvXpqQVOFrif
PCJGHC8+Q5TGqZFgnN3rn2WDhZIEs71qyjtREzFgUSz1L3hPYRmg/7A/gf1Eo/hP
zPNCMbS2WvNC/9XdGlvokXCp/k7GcGpcUCP4kyBgmEUO3arYRFIgCl5ThgIm8OVs
S8f28mM4x2Pv1Tn8Ixy7eJogL2p0d1VWmqHcHvAy3a3EN9QbK/e3SUMS2wyKeJEt
gDYvoyKTa/dfQqNgcxQBKovk0E9EauC7bKISmq0oxUjrWrL7mVJ7YhIEWP3LwEyq
TJzs+nN0KpUwzakeOWb3Op0cUPN7ef7o9jx2W1+xf1QR8zQDQMWj0e0G6YvAMPDb
f+TaB9CsQBmMpZpB838APM+rF0ePLBupYZj1RWXDH8wyRsr2DxiCKMEPWTeEkARy
pL9nnBmFM1Qvkinq+Ndtiug1Xr8iWMUwyYwL48a41DvsT6jhjSYTxiO8h0aIKo7W
FgfCJlKRwI/k2ZbS7HdLM5ii9Ao7S8qPwW4pFydJu/5AR5Hb1RzHWj2Rs+ekwWw4
x4YgCpORDMfKbokZMEM4NhZCtG8u6Kqg6tnLlJwDWWPSsfOXaUUHMd27k3+FIaCc
N+/H+PjWpmyYCP5aZ8uNNL6FVJfZx8Jy6ysJ5GwgtYIqv0mIguLGlX9MF6Xs9BEm
hIouV4/gjpQJOCJHMtZlVupIVNZRgJDV9nLTv0F9sfPOZoZzL8eApPXJcMF/dXlJ
PtztcE/JvIO128nKumrSWkE5lwAxyX1Ez6Bpj/1TahnFL+BIu5rPY4wL/Cr9i46S
XO5yNuTkoccegnZNu0PQkOP0pviASbZuXE04ApvXbkrxMKUjmN3BV5+GcjgZu2tY
reeKML/W2p5ukOGKANBl3lDDubZei1JJcUs8tLMSD+slodwTCfe5gJG/NhyT7FXc
LLDMItsxO2YI6lLv4x7Oonl61z3ZwzkeMUGaEg6hSEe3u1wZABLF5E4Gz27xQBT+
y/1k1No/yd7WOVu5NLT9i+x1gIjh+5L87mcUEB/HNZ+w4EL0czQlFW2JJd/XGScU
c5l1YOlM/kUJQjNVK7JIQa9ve1yD1R+xtAvRYzA5xU3ZMNRbQvcs8JReSp/IIkHj
T91oKkkGToCNDzEoSQWBtyGoTLHz899dICG9QWTa6PxRWZdfS8N//frH/zh6OsMi
FZoiamcAnhS7+M5KR9tOc3qdm00NuV5fY6FMosXMRD/UbXEVA++VHfe5wN7X6O6Y
y4uJfoMPW2iN2tA311OxegvteYOfLg7i6CbD0I2zTk0xLb5/OTS8F6MiYfTRex+y
3RaLdZFosHB2Lu2eW3/9B/fIi6BHurdwSPbs6+VGJm7wk93fyrohYLzaIDjSjsFP
UrlXIe6GsZE2a58J9d98mQZGnZ9yOpcFJ7ckf52yzNJxsZAIINEuEhU4FBIMq+vV
eRtkauXBTtA8zUeOz5gOY8jfyonEl7PcIto0BO/GS5Py7MFe0aKDbiUtakcHeVd/
wOvFZb54teNk1ojxur0bbpDikdxZ7NgBcVe7VQCHDThwVz5Kyf9gML4JXkGN8uAL
RCWkhRXBR2qFz40tdvKF1u5AxCmeKr12owzOH0ukADoQuOPVbvz6ehQW98ECTnoT
yvzpX4tnYuAiSjC2qYjS3b22BWv8T6zJ2tazOzWE9rHnJmhM6asegnJ8fOBf8N8v
ZRTf3Fx0r0+ExSO8bRO3Jreh8Iy6lUPZ2FSC9nkJZadpCdvx/Hu2bAJFYQyZNdlZ
95sQWxocbPzzwz43r9HYsYXNIsqS3WIU4KGDnOZWS2uAHHfcZoPNWYJfpgsa14Yv
7dUkfZv9AxSvn2Kf9dAJO8ioBVGvhXGb7l6u/VeoYCh5z8bsc4dCHA15CKBNACI/
N7+PMx7O6dCJjP02MCsW4bc2680Ls4Y8OKX9KvMHLX+Tv9+WUipLa01nVD04sGEr
DlVUtiSCNpy6yU8YOfe6fXFIQwjZ9Cxo6pTOJPCBaGg1b7p+rak23Z4x2JPOwta3
j4tok1gD+P5+kftoAloWUYqSQUTJK0yIE1+nCecnLAdu0sSSvPhauh0lhswrS1MV
AcmKujGi+6FEwdGnC0E/Ous81EeCsTQl05pEMGj//9NtOTZ0Ncb+IGhp6lfy8Au5
XnP2I1H0YdMv08lPhnk1MdeA2UW1qb5OF5ZLs43tu4yGcZaERG9i8j/MN+OZV9rj
PPhmo+N7gAfSaAdvZ6prYueacHhIZeENOi8nq/YQSbIvXIq62/CfXnkMrBZV43X7
tv+KJVjtCC0PqcsWx5Uvbm4bnY/4cLTBqrnvE5RjOGFmGZA73W5EZAtWupwCiMh1
pmheTYqVCx8Bt1Kb1etHcpFu7mBK34QPHd/mUdOYZ0Z9OWPvkEHFyF8sXyRBvSgT
2CNYROj0DMqG02DVl7DdzU89VtPAIhXX6HyZxd1fR+ywUUa5P0V6aML4rmm543K4
4kWdlNhU1yOvUPnVAvhynXms3oFQxEmwri/8ZbIYJCLDDtilFItJEFhorvm2lDqG
45w8yCc+KNIneVPhJwaL3aci2e1k2vodHFjFOROzXaFzI8wdQS8NWxeVvD7dGJfB
LBTlpNMS5PhgO/Wc8d9OC1BaYpJdY71Q46fZf4ND24LpfbO4/ZAAQ1DfqTiBL1H2
6+T+NnMHEPfrlgB51XwMOiRpqHNEVN92JZiKmJSYxW+FYWPDsztnKzjnmITm39yI
BoGx9uJl1CmyLHXgNrHqKt5vtG+cmtOyaRvdX4CiuTjlIBZCbOjoCYglhZihnTsi
lRTtDJSqUA9k/RHG+aw3t5GL9b4HWPBn518DkYg6Le/5iu9opvzPyvDo0Y1D+zgb
1cSk5C0V0UVOXnPv96hEwygxkYJvIqAON0YPYH7Bv3rxsIyaye6WF7H9A1bSzK30
O9NZbzQAQoYi7qySXupUNpt+15zoyQBUsb0te8tTT8oEETDy4aceHDYCNP0JGVNd
PSKaFzfYG1nhOkm5xWstNJVQbmsxTEI7tm/2ozr0uPjXg9sc9xpZ9bTt3r30kYuf
8fcTSi0Y32++pcFRK4UfDhRkT/2+fUyDPHhXp26CDNTeUGdmNJ4oCuiw2qjqUF0C
YOqFbqBYwPJBnJBni27MFWRI6M4qWObWPZ+jb4o0flWNuRY0X5hWzFVLvYBtWorB
LJ4R5b+On1Xn6Y+VZWQyKtBqncmiS4pLaQV9rbG50d9DLzN0njjD11d7cJqi3v+v
dzhAhof15Zda7hPK4vs3azhFgRSsfg1/zm5pJ0+hB7R9gc9YBC7aazdHtjhSfo8G
8AezgtfDkWnQAX0q85mXqpzpLc0YS9DJYIH1nZN/TFFAFbjn6PvyFap3FZDWDYJE
gw+J8q6VpJ7XA5+6FAWK/jeFp3tJGUzTY2zuVwi6hLIAbDqyohYa1q88p+q/oI+/
7bzvEPT+dFT2MT0ubjXp7mHn6TpLKZq8TC8FZOkpInsYoTdYOhl8TXxNxEfcMeWg
ZKG6q+cCnZXCN6/JytGsT/9CAHgHnVge/SoBE496awHpdZ0dgD+bjws8rybf7pKd
5QyNaTKirAXS7oIhltuyOF2YKYc/St+06o4vtny6SnRfWDCIAtdjM9Em90+kOZKD
8+QQf5idMjvrecBRbeJ7kiZkip7e/xDxgS3RG7gsz8vbwWofDxH7wryp/6jfR0nP
0ZishctBoytJx5t9tJw8dFp62ATT6oNh6ZAVTCIQV4mvxenkAgu7lRJ8PfFBmlc8
KJnbwfoJ6Y3jG8kRZ+Ri8O30UODEkzm454gXK8oGSTIla6TVDM3jIz3iCAtfQs42
nXB5uCrqMisouUQM9hZGWMwfGw2sPlPQcOhjAZSaDSjAPUsfB4I9lfTTHTzFMU1C
LYz4gFh2SA3WyvZKwXNTxTU5sjWM+Sb84lTTlBsVMaO3zL+N+fH/rGGPEfjp/vh4
XxJ7QMqt7Zi0G9kKjSCTOwC1lvdWi646ANxYDUdUJClUvMkQcSCBlpqV4cFG+Tx4
9xDiOe6V0jGANAdKSXj6tXGNPbmNtIsF0SlVJRqJ7PqoxuRk+F32ZERPQ1CGIzE7
vpO98C0lAmTIxVd5S31h0YOAhU6gg6L42nS6DOlg+0s9rA5K7B2anwSVWs+l+sT/
d87u+6x2ydHFasRq6feb+/157lclQj9k5n88+W+q+QLOTvaOyOM3Kjd4VqkAFz+R
8S5z2vGS5xGz+bJsBx/QaqCzHZBGelFJgVEMEfdWdIkhYRDstzhWjRnVEhoF7ChO
en2SWQyR1w+1vLfy2ISru32LTSoL4L7p946PE02/Up74NfYt8CBsQ6VUNfFUCXom
W0wwfm9BxJnp021w8tTeKhobr3Ad1S8zkKuDroZzTB4LEQ8WndPgRYewkKHPDlVH
RPZV8yNVrfE4/yZ8Y7JTgeQsHwI2XIKgzfH9vCxi3YHpKf8Ov8JMmd4WY3Il7ke0
f2oxAVqawKKhPQd1xRfFS443rBd3uLmMpe/1COinSgMW4KtYEA+U6YFAoiSZUS7w
X+VEay8FWckE/7YTVrKVPZBRKVyctBbZ9/oGxbaa3+IulgQHFMNOVYtFtD8wlRAh
wRnwCfE2dLPYya9EjvRkJgju7W4jILjV5s0ElrGBhZI33yLbcRLujB1fYF3OrdKs
9Hx7rjQXfqtnT64yntWV/vI5wWZ94rkVJf5BoQzOL9WghL2/2dUBrkf91smwNUzt
vjRupJ4Xj3Nrs88IzL/w0UKS7EVr1vFreDjEQybyA6PDaSqbhKbI4gkA++17APOo
DbY7ZJJcp67lW2G2UBjQPMM+a8woA4uvF1haetv6ATooLtiND3ZF53nF0RsVoz7v
8PYg/wTEn5FmXtVh9ZvqIiKMxV+J7u99IOfyVp7u0jLPTDKDhXlGw+VXlMyi71AD
d3CZyhsKsO0iBcxX3pkgob9c2qTzgF0O/IbbWspc/wGr52KolZivvlkGy8SV1DjL
uShFxhY63Ojs0Nph0Z3uZAfKXWfJrhYJFdx5OTCIKhcajmPGOEoXBMCeCt0qGR74
P2e47BVYLQY+9S2I0kcSSnHAFsB/ROgJPx01akGzZO2vc4Kjq2LyILCuRzB7GHC/
QBBClauCxtyAnAruxR9sFiAgJoccwHotknEl1hrT/k9YbSv6mnKbQ2b/F8oMusOu
oC0sULwPrlRTzX4FP/BHO8Q66Ba4o6CqMTavtbzBa5T2vN1MdEVtvR/wc+Gozv8I
IjPvA6r7evtCIlDpr9mHcEuWXSTbqEXTTSRrY6wsGWmOXiPfBKTjZOWK5R/pn2d3
OAFb1z9NgYZeUyi9jbmNmItDcp6Ip3fBbh/cjyzB4i9ZX1PVoxPqpYajkwgmZ3k1
14Kpak1nsttYLQB9S4dbRwzveOP21GEgu5PuYLNbqoAiaNkCqB0S1EIJELJvkx9R
SV+q7pXjTB1FGFmAI19WXqB2aWScyxZ3P2DVnlOKLMuD2OeWbrKUtowDKYcycWh0
H4qLOFElpO3O2mw1Fg3zMeGG6Io8jTvsoxC4z24e9fY4XVVB23lVCKBwEQKAm0Dk
h3D3R1yau9x8qiSTvil0okQXcXtxT6BX60GG1+8fD79RBRjHcZMtAF6T/dKqurA+
FJ6P38NY0KpJRW41xMgMOExTl0s6vh4dFGgOg38fKhks7YOIyVAimMNVF2kGABvU
YGL0wBm0xlJKzijLvisiWx+iyMBCQMRu7QVBY91D4uei4KCf4b3ePeTvOtUsJA63
Xol18qM/BNY5r2lPPdK3OuvtIsVnjUGWuq80DzFwHRf7A0qHKfdLglCM9CqkcHyj
AWf8ILLyF9Ue2oGVLEC7HwUPy/kTPaTraMHUaawcmzJkeojDKw3LIumtcDNyGgCr
xNQDOQiEYaihg4wVfZ2zAKRzlDnXzBs5lY5ixU3MOEOZHVmBkZO8hOhwSoeVh60W
jFZYZ03Pk85bCSclpfVj4cOb60PNUVscyU6z2MyG4JxCC+keTz0YiCJAAOxeZLxQ
qnFySTBdzpXbqTrvW3tR/bXU3UDhje45WVre54A57Daso0UV6jLmi4c+7aKnKgdJ
+ovEOQ3mrhKhZ0qlYlp77CM3yC4/xb3b4xu3NnGZCmLUNJGOMQ6nv0hVSX5Y0va/
xMHh9mhwY8SASVL1zF6aFoNDHbSSnmeCizHlk9BRiJS/MHxy4w/nZz7pKPHjcqT7
bUKrfAi5Uea5kxYvrQm16Nwm2Z14JcPpOEuSMU2lylX34a/CkwZQ6qg0/JBvUPh/
1917r1oviEXH8d6U3jcmEljPtsN8hdunVGtAGPAQGHXUHdhEgvqQSIpvqG6A5OMV
ju9lLRxWpbuSwY5y7YMAR8HH4yUrzEgkmEOQnFbgERMB6XEwaCQlM8OpiY7yT76T
etBRLv7CtbYhDMLjeCS3Dgd0QNF1MQBl4Nq9Vju8CDp2MH11SlBR21HJyXw7H6ss
0Q1+fEr54f2FOnC/0kyoW05h4vGUlnqtOssFARYIVHmTy0zH3cwKOS2Bidy8qUm5
SgEwtEg8hqTy9B7j1fUrAM/lncBxPRGMe6O8eBXd3CjCbbngUFHJHqT4xXvn4Z7u
PpGWVw1ev9ObBs5umt81My31uMJKq9JlY9ZkjgykEOIB9VXRCnalUaCwERbvKMnK
0QF/+G5B8bAXCtC8PBQgTD3oUzqWpXwAWyer1bwySxN8E0k3eNaWcT3Y0JkaBoJP
ghzdwQjQ5wzbf6C+XDJ4Rt7KUHkyuocfQ7siDOMRspTmhV2UTmXrk7vdn+Jd171W
2KR227SiM54+8iaYrWvazQjzQBPFXAmcQ6wWyXU8EFYAJzsLF7bwhNuOL78VyKR0
+myWdN2jsO3RyeQAFCpJoQHRByJv0NJKxtFEH89ypMtaeFcU0IKQE6wefzElBh5u
v+5glsxtF7yf7ndO0mIM+IxXUZui3PsDDqh5Z2f0uiQGjdWvfW1JNzQtj7uymqpZ
IsDhEcdN+qyhhA3EHEzggfRbCLaD0bCtxnaxMLVCC7+cNT5lalNFNnMEduMsu7BY
ZGGsxsQDp63zNSlWCHQxAPiOMhxsqz43SYyxOiOfrqIyUsb+CaqZRcvMHt1pfYgq
zxiqjDZ+Twz3QeCvl4nz8bsmk2Nyk8XsBbR2QCqeAOkfncHQGuv3/1BKtg5lFveX
QbSs1yurQrJE5Gkcpg9mh2vbwwJzkg5GDgw2ERopdKYJtff8l3NcMDlna6R3J2TJ
47rvNJp/43nasEZgj/ZWaH2/PFWRdIgvCzypagGCjekJUTmIydglBKhGIIARb7Dd
dJIiomo/FVVbuYuI/d63ZGRLh1N+8FnTu0deMXde7zcxcmJNmaRsSPfd4F75rZym
ZC0nudwalEYa5ID8PlIATZmpbFQyJkHFh0xYZzUTIfRfvrR6Q1dBumV07FzPT+16
Yy7+4d4sPZseb3m+T74K65ccqjOk77VrRVfviMrV7pqCPotKpKR+3soga4JOuiEJ
kVc72CyRfLS8gpHeVucjtZXVcbCwXVHIVwpQEqAGyNGQYmAkzkfqNQcx85/ql77g
s/Sfg/39Ayc0fURp4Ic7QfZG3K04g4diCVnmTXKtiGVqIw19tZRFmyYb9QZdufiO
ofDhD8PUSwuR07pC/hXOQbN32EJk0+XhxhUx+/c2MWCzLumLBNx5ZDm7Xr45WT2c
NV/RLnYfIFzgsQcHKRoEsi0MMmX1wau1zkNGqtEAH4D8pUalBFzkrP7tt1wmkJcg
vyvepvqggLAxN4CvLBC3ihdx+rD3gfup6STqe/uBifBzr9B1Y8aB+sCXD0utQIOO
MEO61uACXdF/6xdEsAJfhY+NE47Rdb1lHVY/Yf7Pd6DmBASrYLxbSz1mNotV2dKS
7pupm2okjoOINWAEc1J2+/gKXVvpsLUeTbawGRPGFScH3OJfIJ7FS7BiqpOcWYL2
rpdGvPg1e0UknVNiKARb5CTL6+liyR1KdlGoGgvcMjGQ5Kq7tCNhOCq7dC2Smt1L
/nk0EcCsW+9TkHy2v9HRDWcwAhYzzevSDBiIE5plyC/6ckUBsMPb9YxUReR5QRqL
y3czNi8quolLw2VcYLalgNhdgRVezdKuqTgS6Fiu34tw9ghUCml6cJ0ZzEgZ5UEh
0Pz8CT0GASHHSZdHJ3tVxAuLgn0DoTBj/N8LZ+KDtAt/gMpokvBbjrwMQcTJqzMj
N62ocT1lva89tkCixaLTfUS1ZOmqesGGeifXy53EbGdkO/I9bvLMSOvlyXQhPql6
nk4SBi+vLxVWy2pp8nCZd+1XQfBW4q/QnZxOnr/FSsumTKyVIvOnUwP7YCUTtW2o
jUB6Fy5YIdHLiQXh5bT9uJ+Vemr7R39CE8+ZSQM6OMC3d58PHr1nHY5xmd/PRU21
xJxQpNbYxHdwuAXr1Dn96HqST/UC+7mWcUcVbWgAbN96ZP54E2fg8XMpk7lff0Gl
GpwxZfLiFYwHkaFv6mCLRVSu265t9YMFvJzFWNUEFIptar/k0tlhti/noy2C5R2C
x91VtCbRzVmjgYqse4Li/2f5aYuZIyVarHjmBD/ief+So/kRdDzQOUpoDhoGpQxS
O4sq6+7akkVaAi2Z/ldUgPL5XBr6uNGgjMD8KqvzdwD6WHzZkBKh88Q+jAnlIfsQ
sZS0slhZtBTR3tCK25aN5PBlFxBZ2pT/SBIjJddjQ8xw3LUExP8+UHRCGSVs7gsI
+Fnmhlu6MLBqU1c8cHDW6+oIRxu33uXmhR2cYaBeDS7fqRtu2Aj/GBy3CysWHbel
fs5XBDiUnk7xPLVpVtHDT6PDqu52LDkJ9pjw+O4yU4Uph+SIA4WWXAtNRMz0w/6y
9cNX4fyvHpTfbRNlmO2nW6ZyhcG5XGkaaTwhXBFCb3kSFYPnBK4ZKOShnmM+rE6N
x4emCG5MGTJZ/NiS3jzM0EFVHI4XvzcTIZXF1E0wuLagHpnC7sNK+oP13dHH432Y
6tQ6B0g46vyvIJnd/+LR5iANKpceCrKsjt9Fs0a7613llU8yof0P831sG3g7bXay
3l7E9sNH9jinrSFu/hh/HlFrZksRMOIlSNtK/iNFDGGMMkRcWZRTgqk3m09QSWNg
vHMsW/VlbUbUVfmKJa/L8KD8pYf3j9Y8j/Lex/vH7TPULuwtNi0irh48zSF98Wxg
6Nb1m2S1yw9Zvk8YuPClCU3gq/Bd08orONPb0JhS0JwkV0lcaeTUivsAzYdgn2s0
KZmeBXbY2W6vQ1gG2E76/FrVHYLT3qxwLztQj9Yyo94bP7OcPyy90UxdXWrE0AFL
tc+JVNOD2A9pZmIDyOaJEXGEr7xoA7+FRX04p5SNLEstWZZhwMmgSIUzN8bOol8O
AeAOqG/0FIy84PTr+5KHPVQ9dFdIqpMi3erhXGkjVA+h9VIPO2zxKKGIBkbcdyQA
OuUeGPWmEDnHJ4s4wZO8vsIEWu+U6r8ogT/3kLt/YjK/9UgCUfWL0y5zDqArryyr
EpI2BmJlcK4RPuAwVZ4GfUiip5UYpk4kH11m5J+nRuAOJf0ccvzm5g6ZOr9i/GfJ
s1PX8xyu7/RzMI6tSTbrtEQDdkoXN0etZE85g4A0I2JbVPTpd49kEleAOSVQX6GM
ZQKEjRd2akHFSCFzCBtJk/t0YTi7s0sLaQG3703JlAZvmH/eoUZdd+n2kZcZ1wfn
X+W/z+POvjvfglYRzlwF7pv9MAWUfRKwlPxVu/t7mNkj83WrBvARF0H/jSUTv583
ix/a9qblMuoxBwOCffc1HQhagDNv2zCbTyHkaeXAe9RMmxn4oXdzb9+WN4MHeqeb
bQHJXVNrIBFeBq6kNxvoGebFWLrv3siihl4pOR9P5ud1SdJB6yL72fe3XQtqOKfc
gjoBKJnzEwbKWqgvXrIKEB4jzlHHC+q4nTtenIRQJ7GKYCql4LJaYT42BF9hCwZh
D+FYx8BpD7Dh4DNF5Z9w11qIWKk7ugS6yqH1z05helj8VF8aHnjlwz2+LP9o6KWV
0H5NoTPsMSqM+zIPQwq9caWxxGRaTv04VOMR2giPiVb5OO3dhFiK358OGVzc8EPl
rElJlzo07n31Ef2ikLEJz/zo2SmqXy+BZvNjs6QlGOseWJMgfhEMAPrY2Y3TFLyP
UQ51lT0A2Kt0iyveAJkr1fkNtE6s/c9l2ty1wLeTbtcfTVivVmRLfBIL4NWM2cv7
NzTnYlQ6xah5LnXZS1AVu858Lq0cR2eejU3Td6A7M5Pt8CeJtjwbcWbhiRcU3Gs7
iQL5wsEXZ8OFqpU77ezDYH1S0+spe2J/+Qk7fU4h49f1qV9tb/qbkMW/ndPg7D+s
N4/3gJTrH8/Gpzcvvd/KSL+S7u2M0JZSGKKufgcfPMKmpYOYe7ZG4SlMDHdp9i3H
gWU87iNW9L2cuwJw09VfRI/s8pBM1+l1fbDgAn0YbsWWT9WmETnvB0CMjLNmoQ1z
BlKH0ZAusvyiJHggB3D/cg7kZt/jfiYfVrq36Izb6HQdHs9+x1Mtlq+e4GSI2L+n
MEGTFLnDlGi9uGau3gUur5InXznc/NhbAnh7ZWqlbdKIFJqedwi/wg2rr1QxoXK9
a81vkFsRk4wYph1YJvKXOCLw6jGADCgzUr/yD8uTEi278hfVQTl6uC5ocbBUHvFZ
4N0dNGLPijLdclfrgmGPBAXl3h0G53MEoACJKjQx+6ziq7s1UV2h3w6I/LxWSP4w
MiIl6W6Pp78TZ6CKnW95wS0+vjpbI9tyjf7dKMmdBrwezJDnxwNoNOBPa2onrO/3
oqNucY3sHX8hCSpULiuvfVMKv3+V6qcZMi0qmEJMnGC/H2avViPjSM0y9NclFZnE
zSlSjTC2nw601u2fXodRUIIjPKChlULuH8hdSeylar/T0Kp7hHn5SdbzuVoqDsH0
Ui7oatzLkF0fDr81sTh49DaGSqbiXQPuznWRLDjrPFMOPcGIhdJi3TY1Udq6yOoG
ty9TkOC8TSPa0Cge7aEtjf6wfiEU+awPu1dlSC4u1Lruqb2a286gLBNaUlh72J+v
6BwT+gVzv66CKIZ3F0fWsFPjBNACxkzbQNd+VUirogedTFt/IoY+Mjs6VBLR7XCU
xEYwWtmBbCTvyPc22I72jwZ0NyNKVIkGF9FAtxDS0rdlSemZ/ebNg8PV2SrTHA5t
2qMr65Y0vo8w6UG4+Ra4zAKQYHh3MkbEvKVjrLVe4UNJ4888oPZ1HT2alnwnDDbq
DCnbT7675xsRH5gs8eyTk29e7pAlCBIvPtiQZ7/v+88AzTHOwRRmPVpu4cFmEQjn
cst95jLqPguL73he+e0tVwom9r6PiAQDEgWu2Fr+9FAse5BTBM7/N8OWD6dnyb7a
Rss0DOccuYDPjM/m9IlLlro3k6iGnXgPd5CFPFfN3mBKlUoa3HbytZifqcZ8WJNC
iMhCvjuRz/zswierWAelzANRKkOnU3pZUeR5SfNZMQNOF/+ADrhaEWAXoafcYedZ
WZQUBrfTQ732pZkxyQYDjIt5AaQTtpyRxpqZHv6TIBxT3ayMX0KVbhX6+FgwYVjF
qm+pDdspw67aR2vc9Dku7K6QqG3eQ9zg7J5y+vYzCtgdOZ9ZxDRfWEYr6TAH+2/Q
bNeqvcOyboCAFLqPj+IUlCiBYcu45Ykh6wsHSbhOgaNZgROM7w23Z7JsZKYt3hvE
AVvudcgesi+xT9xZnWTqE0qN/8QABUuub2I9FSRWhmpRh+TIlaHkpl7eu01BDQPi
tnuqfF5u5Bz0msolm38C4kSFJxMkuXHUlIcbmnHuhimFdOA+lKWpKoumQBBy1kK2
UWxUpHJaYaRxhSrMRO/m9ulffkJunTJ2ZezqUMGohuVrC0gcoDiSCskB7NgtAiAW
Apw7Myfwn73U10TFX/eYbZ9PC/Ilfkqn46W8vE4mLWnQmSuU71VYnBYhRAc53eEs
8Pg9MviZ+s5iCo5CKRVhE5u32PeZBydDdYR5c5slUhrK3BdwpNZYB6acD23aRws+
pWLe4zR0hvLg/M+vQB1HzRBzPenblMxqhQmsWsglCaSmVUBBhtPljxXr800ckcva
aUW21a/eWVmbKyObpRdOx9NJmfEphgcwbZp8QaYaeTFs/TR2FMnuWuM356g9fQzw
+X57b2hacLJYg95cyOJYsmSejWRQ966+6ueTNho5v5NSHsXjvsfOftiw1MkMljMu
n1mEcdKogsV3uSahf964UsWbfgegXznZPd5YejCztWqphY15xcTaj58+FliJrzBC
b7IVL7r2LlSIReCSphy8qgN+f0MUWmcR2tHgNRacXMZTgMu6pkzPMPmYsEACjtm7
8u6AovjbXlMlL7lq9EfsT/gxMI/DYqkhMF69mDx/JSgRYmnJpWqanfJneBc3E7x8
ANaUlVdxccLf8Gq0ySbZrvsN1a8wCi9O8g0M5edh12AvQXK2GeabSbrZjyn0ipRA
JecwRQIyV7DdG0TxZJAqYft+gxAEF45p+JPJdJG5ebqolrKmbMDLELUbu7iqlGzo
aka/PpIHrZKnn1KAcT4xk08+fHe1r67kgL8KramzRpiUaI5Y++jb48av55VbIHhp
gKEE4XgqijD7afByVXjuivPh9uCvNQXl2ZHgeVvgVLd0QsEwkiQRWf3V2iM9uPVy
0RYujlfcPpjVO9dc/ALQYFZ9gy5hFU0a9ytJyDN6C7SbZv+udrnrNWFfxzUwNdug
4AJBXLSzCUxND3/CGgaJJ0rNPbIeXuTTvGUfqEeMg3F+dfoZUX+xcY18hiuTYDL+
KycTT2IJF6qFhgR1L0gPr4BP58pZrWPL91+NjKSfd5af1h2Zq7cuMDL/QW6APJzt
841rDKJR0P72PQVJABmerBzyHKgmLdlNcmwTXU6XBVBcYJW+OuXr5DPb9YiDxics
xwe8QDcP2vzmtWgvhu2o7SlZAhoYH0T26aKUjVa9egpHzGQbb4myU7Ute6GYzPjO
s1V6jhM34xKDzZnX3XECV6aagoztCN/fO+j7NLz6hmomk9LLNHz3pjPLQR7/RRSq
sqQeK2offnnfOCnrh1Q0MItCBN8JHLI+1X/EejRgftzJ8Mj9GF1l32TZ13enji8O
rvYqc29kN5Xqzo8RnhKnjx8l7dGx7ZbrYVsm5oVUW97tocGiEubX8i7OEOhe4rwO
YEALsfzejrqUYp1dBbyuz5ieYxKTgw2GS/wNQ/mtFKrz/jF59BZONJ+SYyMb0WCa
ckcA5WBKGujbYx8O5Ljq7wGefPW2XBYY5SFDj6vTVPOYx3FWc5vOTrrPeCGS8C3d
/8KN306GuyBfLzBo6dmH0NOqOJADWTisxtPDmVe9C9NoLsyx77vqGlu37hqBn7yC
Jc+PI5467PgMny5NyxdE/hH/oQccClPbYL4u929FM+YGk3kDg4f7aKWZtZ2F9eCX
2iFgz1Mf0GP+r4+aErBZAhRkFwXF9t4QLYU9EKKe5zfxhH6k6XNBQwdRwuupzbXP
ISLqVl5LHmY5SKclIBo8gLRE8YoQWiZnuU3T2kQ1NRKJlO7gvzG0xNrJURWEo4Zq
Nqcf2nWvj2ZekK20Sv0lvn5DHYpI0QA+L21739egt1O8//7Iq7hKomtpcjU9qO6K
wAZ+14Bvvo16+J6ul+ocrXftSd3m92TvyqHMtgCxwVDZVrnGqm0e5ovq9nhWkMrC
DWIBEoRtARqYRSmHPKNLLlqQbXRSrcQvigWPevuV0mWxDmuiH6FRyFSBEM9//Kqc
D1c6OsBoJ0IO1+zzUFtTM24PtF/yfnIGjYnbuDitO3WQHbOwS5ZKi7QBQUeTsXn9
WWpHSnj6v0+Gl8lNC84CElvsmVJTxz+kau4XEjKH9zo96wUzxRPYlhbxtXoBDYGZ
A8ZAT9tfFDK7cIMcptIKky0IWOmLDnFgEyNIWc8NEs3F+PONQCBXGgnOG1v2Uida
SMEnbH7HNukcST6QBIElXzyX6iM3/om5ZnC4152xMfzw3svZjEE7MlfX8L1RgnGO
5PqKyTo1IYWpBnd9mUJQL24lYQ7HLOOCsNoSIs8bvp//eSsxJej2g7I6ixUj8gVg
WxJaKR1vU/+FojcG8a7Ifz20qcpOvvMijsyL1Y8jtORkF6EXTQYruhR5Pi5W06nl
9RQteOEVi70QyQMb6+p5uNrm/6dKciVagyAcCN3TQxO4F95g6+PFnCQ+UcJoX9AG
78GmOIjDg8n+EBtADNmvEUYKHA0eC6sjydJAq3IfLzV32kKamS01kFFJ1M1L0Y2b
sVBRX+NlvC3VYRIwzfnbvmIeKan8ubXuVUjYygsNZX3KuQvuvdG1/SkHscj5xNUi
pISC7wC9IN1ZCTIu3ZjTyizvxuXg6Dk78fFCx8tQ1/Qsu4PpLSAB5yfYMxqlola7
EiKhaY+bshE+g7mnYE5MMC/Y0RVVmU+orLlZOekLCssV88z2+M5bNPhFqQPGgzlI
CVZ3Vsvpkae1BeISYq0FHlPPi+E3SAapRwsO2cKXaDbihGd9D/4saQ60Xz9SEsQt
rPstUqi6+eusfhTpoqgiyi8aLcsk84p+b9TVOOby/T6sptDX5lL9l5oxqnEjFsmp
0ZVAQLAuwk6G0cp1971TA97kg7sFVFK9ZQk/x4DGEVUBE7NsZdruxsKjIbamWcXb
JmzrafqSr5freyXwXkjmk9eMBnH3QRyihl17+WGv1ycaczXQxZxJLDDQ8ENk/a0g
UwbtT0PnA/+cTaAkVvjucCQlan5PXrompmcM+182igN6tSJUJ0hK9XA/a/ak2pyu
KSdS/xklRSeSn2OpRjnYozxGpDDJghr+lfaP373YHhNwIVC4EETQXsD5JIrZStpU
RiPjp3imLYzAdJoFOWyym1JhlmRWjh8M4fc4FXIPFtEd9/DfA4rlWEYI611QoR7Z
SbLqCg48tpoInXla/GQupw5PdFOf8CaLRKX6ek3nwqkA62uD1UldFTmfA+vpLYnd
AN08oNJ1oaZpx4W/WsFczA5JeT7aWQqDQUloQMosdLWi4XAApletcMAbw6yMndzr
WWjcESE5KPqv66mRJZ1Of4gAW5lihs10KA5ZUlW/H5knPX3ZlWOpr2N14xBH4IXJ
JCGLPnsHSs5UeZcDXc3/SuqQ0N8PASuAN6DzLwpcazrXyL3dq1nb2JPr5iKpW22Z
I+r/LA1oHEz7ZPI+wOKftOTGRk1BbtoAEmWwz/Ib4Jx5T1gVy/Eq65HY4eRxrnY1
hmnmXQFjNn5mz+QN5RFGiTUeYpjPLgZu/3cJ1owsdBwDHK1YfK3GYVAIm90sgt5v
tnRQGR5Gw5cZe6EoOTd7DlOJsBtClS/DUU7Am0tGMhXZUx1DYB3epXeas0zvCdUT
p9dfRSQax1HEqsmosG2fDearctS3mbeWc8FUK42B7YPNnZLOnYE6+JPNq5YmwvOS
ZJqc2HqNto/S8HiTyh1mlEPj8RmK3bQawgbJ+4NmSo55B/KNrLjbHgHv6WMlKgxX
XfQiDKyMuI0f3QYff5+eN+eObxInYO0Dy8wEyeCuf5N12ehEiiMFFkzxrnWfga2C
FyXNn9N+OGE8Wn0aMUw2kri8D3yoz+7Z+bvx2I1JjSp3nFRY3i96BovXWXJnsUYy
xBRvsOS65Hzy9sqbAbeN4GOrbMDesaafH7K2AOOKvl16WZS0seT1i6ARbTZN5EDf
KTiiSGytYlvGSGV+1xf1qe+hJME1a7SSX50L3JoN+u+3z+A4uzOv4lmcL60q3mDP
+pCo4dClm0IgguPYhW+egFYmafH4gp4HRFITY4Zcl/CrYMzntmznNlpZvxbpJAM8
amOMcYUHa9f++DF/qjt0yu8/blkGB2BuqHgRAOG0noF/5mdtLeoc30wbCMYTbnda
V/Oy/vz6+9owraOcPyjs/XlsjQ8wkykWtxLykqi2rMm6XBMTqharm+jYHM4kcB8m
Ua+Om7QMnmE1c39TSpkEZKkV0UuJ1FW3la4XcWRlZMB8Q+Qk7Yd5tHGhvypgo1J1
ROXlJlZwJP49ZCo7SUvEq8xNXLxpbXEPdmBD00axW/9yglJu4Rat0Vl4VIb+o607
SJrPxB6GBg8BKWP93a4WjWuEdsNEsrGfMA6GIFOYralnn2eq9/ox5ew+pXeNO7ej
5hFwOE0vffoq8yQKa6nuWHmQQFDl+vRAxudDaPVac7iTskK7S8+3f+CYgQSNv3t5
GqGWHaGeF6X0/sDOIj0Ovzm8BaH3IIIZAm6oPWi7Ta4NXN+kiA7U3HSp5+4G6cZ0
kS4GAHwsC7NxiKJT0b8lTBLeiaFbaPCVhw3jMC2TFeAic8VvrqENsX/PDwivnUsH
pRpxhMO4EsPq47K+TSjyMst697vKBECmPUE4HCcoSTU/cU+skoaP7QuDCPfWRUrD
vvIO6BNJJqjMB4b3Bo6Tre4eMFWwaLhWYp+DFoWmR9Lzb2c4CclbCzM98kDenYnh
KINalRKxu2FFje4nOZEC+uxLKOA1h32RPu4cRTS0Bz8lg5PakDLT2ZvdVE8tRPjA
WlqYKrnlEuz+593F0UGMhsgA+ASzTTTxyUXowiXA2fWIjyHbHat2PwZF8tvPPQ2M
nS5AkrH2SRZUBC6jD3eg5sdn0rJUInXeXc18FyC8BrtW+m9CQhf9mgqWzzSrlVzc
A5DZDXJtH7yzaulgr3sgmb5dBcgnRrpSGeZ5SdmJPPg8CS/afDyASfFeHMRLL8CK
t2/BU33mf36k5dxPUp3O1npP1Mq7D6QMAnjnGNi2vU6dXNn/IjJCXmbdEW1uP/sX
BK/u+YoipE+Go69cXlrTjB90cGz9I8JXjslAqM23AR47y8Xq0H1mX98t9Vtmo7Ul
RbAgsgaHSJh1kDrZbn9sTAWbZZtJddVQdBiZShcqQUGlt7a7fQrW8jxF0VdnSnh4
pnKxZdPrFG0xztN0ozG/usUkLTvIX/38tKTX9wI8x01tLIYJsdCDffxAhFHDUfyH
zbiX+5ebA6JpZ7X3SvAX2GgYlbgCWFrQyxrwgUEo07qmeQZY73ky4EGLJJ6j/0jO
3Wj71Wmmh5KomRUT8q8Agcx9XBTNdS5f/HwEz6flKKInwIHP1hyl3K1AGFpDe5H5
s+Mzg7Rc+H/58ME8UM+snHUTtUM2ilAsNxPAeLS9SGacDzWB/5mcYCH7cacb0TUl
0ADGbwzW8K2cLZyNjtMbu4H27UgwYdxLeNmhHzYaDg7ZAyYpIxbdShaWLg+KY+YH
qX4mx0+nY0JGktQpXCdixZyT+6YdtTznWJ6eoStUyMAExqxe9ADPGKwbG7aPM/vY
fIXDyYMG2ogYUpxHDvNClK6eBqJzqTN3i4vmV35xYIivcxM+nxkMTYyVRx48BQWE
VhOpiRE7MOG276SIVIpsAzP8fWlhknqGT/YdTGqC1WUToGcZsieLcoE33JHRfX8P
tOwbl6tV+jFenqCYsiGuJH+lUeloZC8Sju97IH9FKv5UkcO9VJEvEy2qXrtc/s/B
2in8jqRE/lz5ppmX+6lREzU97bymG7sIKDuFyq+/oXpd7i5dr2Tr9l85RVEoNfP4
v9BUumRQW1OarwZ6gaFTmDve4pgU7KSoj2kGOwsp6yoHKZlWrLLWl06QTzTTPDTO
tPdUT3WsK7v7GnI5ZpScDTybNAVp0ukFDrI7RS0SAxblVhrlk0p8g3tnWDBd4j78
dD24A6bcK+fvZv0VA1jHrvwwII3K/bP+Yt0eBv1RgZhcdN0uMmFlwkep9ywF5GB9
QLiPD/c62gH/fB6FJQmozNJ+nA/TAAG4pCcl45vfS1u08gxWqzCvCfuCjIPZEDqE
6pt2TVMB9ZiQSdYKjfxijQJLuRUYWnMBo2WaZqpR3XpAC/EyUWrGlp+POsahwPpn
apl0DV/OmNQlL8OC2xzHar/kH2UxF3RnLrw6A8iRYsFycHMDukr8yEtxF/hm3UFu
yeFENTP44JkdzRl+NCgc9XpPMdWVfF/qGOwEXzrlf0RwvlhpsTKTqaoOClSms9Q8
51ajizWIUXWzjU9WDNqp5dp8ptRwd9BOiZ6zY5PBjqigjVwEC+7cAxRw3f5+dsed
IUNVB7PP7q0n2p53kLEmBnNH0yfz+ZvOSpozaUHDTSNemAK+lhGB5hy3QQR8HwqX
+2xR5qjzjuPTagEkdcjZAfLEHSN2+rjpGuWTI95h4msLip1nPRuFA77O1qK5iNMH
fOD/6hHE255ttGpOWY3UDVCU5WWx6cDIEzGg1+bg9ehoUXBTOH9DY2xaIOSyx5wD
qzKOXwClAJ3MYjstYv/z3H2Ec8r05swocceVix5T53fnFeEXCeeGD3j0wL4ciVAt
ExVpxad+Cq6VINChJYgQrNPj5S1SZ67NciltDo+gOLNzYwbr4Gb6ismGy3C4oyLL
YBlLFjt/bJWZbQuCJJNzwiC6307Io7wLLpnHrqNGmzQzFOj3iaLNnCY3i4H+mym6
fxIkGjcrQhO2iFGyIanVw+v0sMFFX/TNi3sa/QWKIk76DvRRtwJ49YrjrBu81Yob
U9lBqI75qc1iF4t92siUX2sMi84hsUMgOuVco4R3a/wX/eeiZuIpgx4RrE/HdmEB
boxY2l6z4tlexlFN7qkMIe9wQcKZw4LktxR/7fLiBP8qQ7Jxv5kpZ88dZWIXSqN/
8zW44ofCqa/ZQ52RnRHycoM5Gubxm97GOElKVIsWknSfl3zlyBYVOil1hfzkJVvv
llMo+2mpyRFwgykoiutHHgG4fbsq9mYp8sWQqHcH/tXKDECHPwWp+lVe1vMtslil
+wBRv8J2WqJVNu5W3vWs0pricZwuxzhchtH7SXxlutNuEnYIMQc5kQRBTZY5WZ8e
BahJkz0DyYA0KNjpMKNG7vn8i5j/d9IP+zMk3CmOYAggvNfe2tHFhcSEPOhUpv+g
+w36R9DuJwMR9yq3i6ZqEr8Rw1J2VAHdt2ph7xBqnzHOlxnuapMtcNsPUsFWc2wY
cfOkP+CRY4UYx/5RtGywhnf4LQEbK7pRHkOjPCUfZsBUguEf09reVDIlQdPULioH
gkQX0wcq31vLHLBAy+lyBCzx86S1Y/qt9kULdG3+h8AdxAGSYTE2W2RZ9FbmF2sr
XN2TN87ek16EFVriT5qFFRZPU6wiCpoLkpw/b9K4QM7ZuGMuMcQe237rSbUcXDd/
lVfZ7+SaArDsiwxdB20EfQqW3G2JPL+MLBaL1tAVW7LRY0ihCjTdRRen/T3kWm0u
QycVpBwMANK5PYZu4wMaA9Ur+lyF2OPnRiWlQB3T0rsVZQOsDauaBqZGhakU9Byd
j3BpBtcVeUWZ8+Dg3uE0dPcwv5WwJeB6DpIi/8FufalfJaHarR3HFV80VAbKkf+I
1hig26Iaql28woHSoJ9YLmO0qi/vsZFIyRfFIYXiGVHkbvbEmD8ouwYw/gT6DIrJ
ozhu/098Dl4WtEXUflLovqGreO1TN/W4bv/5joAQqTuI51xI98W9SZFmppC8ZGIs
Y83k009c+PDudjTl/4jetk90BxoLMFFX/sCoFLl1JETZr83i611G2j3g5Jk1T8hU
HJYaatcjaRX+CaVxwhOyktZB/wqrG7k6+u3+X9WLS2/268h7oIa3logqWrhmntEZ
lkQknBbtXHhtZBRhmzWRePSW7ujGSX8NPpwfeUZkfbnq4CzMMY1ujbdN55o2/V0v
CVa1NA2iow0zuwYlbYCDayiANs5vyCqffgCWeixphd+xSsoEC/AItXHAK5X4wQZw
U7FCSPbCHP+OhhYnr+lSwGBbdQ0OrdVS5D45uL141BCTZEZoST8cikBwudIrAhfM
BlLSOgs2RhFG/ql+VajI7bMRb8uhJw6VjYTzx6dKE1xvg7G+yTp4P5cOrvXoAHDN
ynseEUvjrToSrsBZ4xby86MO95B9D3geqMjRzqp5sxpQMJGh2zcQacZwe+Xx1lU/
221KDiRRxNyzjyueZYegnb08VrAYD6ELE+MAEWJAQQhXE68gynA/16Zwd9dLPTVr
p0giRsKGic8RfNMFOhjRnp3+rFy6iZzzz834fAzMokNH+TrBZgwF/8zi+jksMXUl
Htf4twrFwXe9IIL3873r3SKoz/pJMZeGbvI+piemPHVd7YEezbwf4m1I9uANY89D
thIKWhxczhwKvQKxxUwlxH5SB/jDXLSzKwssJCCs+hZBaiWCVH9W9SHYmYyOd2XG
pEKYonPNWg+MJ6QASG++BnLQ6ktFnpVGbqUnVN7QXoIuLLaof3XVH7uXZK6eK0xx
/zTC+tFAY7W6/SNNIXUE5O1/DL51Ul9+0/7eTp6XLRK65i/2fvLofBT6B7zqgKTr
epWxBKSXcszMfwHSmvXwMDjhSUMh8jZsU192IgQuubineLrhR9Idb6ZP/ni5EErd
qMrqvBhQGpJ6UH4XSrzE2aJpjgzaUZs65ihtzf/mF5rWJr6YykMt7uomBdqNwojr
jqQjik3AvvblZdX8rtQHgmo7ScehfYzWROq4mZ2SRiORSRE7O5LtprRmmNl+2+jK
eC9Zv0EruNkLpG5ztm+Qe3riI3n+REh8RyjmcfqI97HEm8CVx8sf+Q3A1ZqH3FDK
sNEePPat5sPklAqv3V7uUi1LUm38LRa4wthgmKmMS8kVIU8Lkahmodz+JWUkdRMY
RCTnxu505kLaIKyAWzgZ8aoLnIvtX1Zjv5Gy2IeJiw86xYDeR+f/P7gua09Bx2HE
2AksQYxSXYZC1pO0jEmOw5BJjRWCDJu3y+fVSMP3iH+9380gq0PCljDTQOKiwodW
XHxRmn95yPkYFVVbWQT1zbf1PoLKJNJnsT1vFd3tlhE6/oZyt2cBSoN4ykXJiOj5
8BK/z4EO2h0xhUyb5rhxQhm+JPHqDJuV2OqC1MqOO76Lqr1VtpNJt4Knay+xqVZK
HxXmdtBRG/ZuqRsqDKeg47zSPa8+zOvb09azX+yWWx24xXe+2/H/rZ6L8ZuxN+qK
2Jd0FG+UgGmVgcMM6o4zux3Ch99aTK02A0sko4UQbMHLwPBcWSWoU2FGXjDQ7JKA
p6YeuNGr63zNYViymSQEEBV7hJW0PgVJEZd//072K7Ig9P0TBvVZSxLz5o7OGvZO
86P/GtTqSGlooEipHQz//U71+S1IX7o7+SjeWq1qPnJThFLtCyldCYXH4YFbK6Iv
D+XktRXzCqLFn/rA+IXVbPwnQRWYyh9XO8XNaxqg9a7jsRdNcubCIrxiyv6SnO8B
ocHgZ6u5mPgaFqar4431D9ibZh3RIkoDDstVorqGAK9705srggZjiRvCgOxU1S8B
ccmfUG5zb6PwPvYSCmLy2jP7Sue8Cr3iJhRQ9U2jnYCn2BNBjvG16SB+j5iB4rXv
5y/DbYwE25W+jQvKEPJt7XozCtD/sw5rz7Am4834QRyqNt/6Dnk1f4B1LJPEw/I+
1gfOgxl77YMpiC2Kv9eLrVPFBpyFj8E+c06hILyJDaZ1qKWJWvrgE91I/rEkep4q
QPc/JXcwAQ438QCOaSsqUlJUmjGH0gfiBeL2yqohKWl7XRMFMTOqrl5xZih+winD
0i5fQPzTP1wnO5c2vWkScW615CmqGbDBbCbgg/Ew8WiPg2ossnFvVnInipT3hBr/
mnjNBPMY3bz2d31ZyNvlUzWHMUV/DGRTHN0LRWOfoccY+NJVMvWWhBfS9gXCmh5U
XT0bdIWNU3q2Skxhn9sMbN98yNXbBKRoJfAPMYcqTpCRMYIgCQD8XS3c2rYK30DJ
SkmUe8TEqFN3k4jTCh/ZNjbVymh2fD1Ta7qRwANqHuCqglmIwKzu1p4Dz+m+yCAp
yM0457Mr17ow12h+O2aUtXJaS/o8wHxI418eSwcNE3zDjQFILSnQMesZyVed8tqy
MUBiTkB0AEP8pbYSZyqKIrJUG/WQ8fQuUXMmu7YoMn4FvBkfUVFwHQcQ8J4AfAVF
n4rBh4uER6QH1gabONMfKLeejiN+b6ZSxZUdVrIQRjJ02foW5GMavcSJJf99JJRS
I3Qsfx3gpEbJVS5NSWbjsPX4RBJIKuH0+rKzqanSD+WHSifxDiFILQ1chlkoxpeh
ZzWs2waoLgIrh9rR858Ms898L6QFJ/Y77DQzK6/9uCQabZIypT2srwn3hYr1fV0V
wmgz1RZwwpt/lEYkVOq0HYFdGfO2cD86qspOyNiqdp2GNHql3SdahMLvPyuIkN53
HYMsClas6jEOafvYUJP9nMjLB7PGibnddAfyI04kPkz2XnRcR9N6L4x3L31hOlkL
tL/rx6V04+lbXNVUXzeIt7UnyuPAlQDnwWGg+NjqjMKHkNqaCHiyffLhx1S+DmXE
n+OM6M1O190eMxI0I8iXc0Ocg+EL07pODgeoZGCTO3LK5AFoOpA4XjBMBtqxbkGg
lFOcijlgwQyLZpuyxUqNKRpmirZ79KMvesMt5pKHzTQBpXX8p3OpBzryYkdUMtpj
XvQQ33aRh3wwCG/ebR0wp7JN3OQuZqXcRciHXLqfStW/NkIM8kJQCLhE15+EEf1j
/erHtbbahVjYf86Vep5Zt4Pcb0PjJ2of+MzuSH9bWvFc/o4oHMCO0bU8Uprwte58
rXUv1IsmIB5T05kG2bPu94T2axXo/sQYQc1mOvG0jxPhvwUEAFksWENpXIKrI+t8
+6eTIQJWJjsnv35Zm3SI3T3vHB35yFL1XmMTIoSiq4XqPr7Dal/S32igobo5Vt9r
uUNVw4FK2SKqsH/tggOthf/qPNmIm5fi9UiksD308ESz9CXa5INTObOb9mBQ4vkJ
o/wwRTc+fYKgpJ0BVzjjPyq8+Tp9wPVVOMCXfxOoWhvzG8IPTKzxj18hl8jscxgV
2V17RnQRhU3KZlPk/M3Vyym2mu96T8zA261VpAsZcE74SByV9L7B+wNTb60MJgK/
5gqoJEeAu7HbYBLE6g9drS1clxkkAVpaaWdjUKY1hiLSCiItX/AmwGsdZhqZ+cIp
oQWl93YOQnxGLb8zWm4vlQxtX5SuHSmPML/qreW2EgEwbJYQy3muMPMpj1fdTQb6
Yp6TzpyR91h0foQqatdMCQ+iobba1rJKk57sX0hZUpfgZQ7K2BpJ8H1LwKlEPG96
GW3ha/qj2zFegC3ACW9KmgowdqS6pkBlw9hxhZ8wsow5EhCYr1o+qAIMoO9Hx0XW
PM+lMJbDdOLynn2nvyO2FFlvkBDNJyLEB4N/GeI4UeYAf+S1NfMYBR0T2QVVvRIp
H0qo12uhMUbdFGIQfnqW9NgXuJ3sho5AwP7fg7itr85IQT/PjjEilgD2jbUfU/S7
+q324PFBT20HSm7D/KZFEnmy8J3d7obyujHsoI9532ZoAEkHzLqBSP9cDrjMETn3
RPXRIITyYgxKQCn7TN16DlNtpvCRIwkQjNOFO3ZK63clMRD4weXnqNUY5dvvZe2M
PyXNMnj8KIydnRbAUvsNu+wL7IVNvkCR3SD6sDc2y/Lg91bY594UrkJRd2vWCns3
CN2CD/1xu7ucfvkCJmFGSdNTEYY1iU+x7dr9NpyYjJ+KiByQoZr+qFEQgqTOlFB9
pD/bKFd9fLAWcTpsFtMn7f5A6g0c2TOJHs3C1lCDD+q7Yun7lrH6S9jtiTIdkem4
c9KcozM7BzHnqNBUc2wxeL/nCWszWZie1y4kbTptZdttPOrohZr37Tlxm1HG2F4/
509pTPTTL2fWcBr7Iq/+0XL9T4+4byhv/ba2EIMNWDuXBEP2qxLYVfB2V3i9moFA
Bf/SoXj+An9dUWNqBpz4sEF31DBWkjshC9aAmWmzgR8qSGNGFSZfjSJa2ARb1hos
pLj1ZYj4VpXOXNf3ucZ6ZsZPWXdv6jwtEDbHZ2opw/N9aOJH0ZUf+bI2LOCDCWu1
PZXP6mTr0HyXJMWGX2skwBwr/dYz4r5nODopN2Rg3IG1JqkUu3j3KI3T2PSVG+32
Psbmgr3XaHaibd7BNHmf9Ys4YdNNgs0tssbL5hxSWyhmNcWxQVF7iivVFvKAFOgo
wUG7ByxlFUO1+Z0WJtwcwXee6nQXXCtFVuxG20BnYhGO7EG8EK08DjmM9TATWKFn
qRN/F86Ieoc0Y6CN7pH6WUe0+dRCOD1GdG8bje4507cFqxV5KzaeVusdZLZXLmZs
62DmhNuWATIuKfxAndCP7yDO36j6CSwuUMXu+mmOJc5fnnFfW6MFfk2ZbzJNNXUd
ZxkWkF3pM0tjIhzTokCNRDg8+N3EONGjCXez/+bohwj7b5ngSizUqCeOYcKXCAlJ
u2ObNQ8Mo66jM7vm6jG4APRsGSWZQjtSM2Qw8Z+yY2Kud8K+z2wC6GlS31xk5rt0
bKSoxfOAz8ALe2kxXXVf+wRt/YOIxSIOePkqaySvsZ/BLHU/Ban3TOa/CNv62ISJ
vIXfWTxBNt4VtnvzIUwgQB13lpGLJurJaBzk3w6FpnuIUoDepPnWmv85E6Oy+gPP
Dfj4UAorLAB8tc6wmLggf3ibgxG1mreCzPeXRz9YXqUm2R8egjJ+YngEIBddjh7S
C1pu2SXAZOwNRQlZfRm9unPa1gDhsssuAaZ2qG0bq4DkBfBH/RPXGzQLobhT+/XM
D63iw1vdepOpu3C6jTLfZHWsOvh4ChWMB3sZADrtsOvFIm00LMmcbeO8WUW8Tl3B
jFpIaW7QhlER6E2APMso42KGOETJZiH1s+LPL5EIJG0Z+qVG8Fjg9REgnwjA3jPP
Duoq4plbJyGBDfMSkHh9nB3BsO3ykL8HODpUeflHa6by+jW/qy4CUAXAo+0uorB3
Gb3zbp7894qwW5m2qher6dhmncLYccaCwP4o+z7obC82ua+M0RNeEoYY6pggzbCh
gLyqFhRvkRr0Gu5/hRjUMo/hDn46wzhsPgGArR89+tcuTLvnCawQKhzYTxwoZB9V
4iWmt5/XCDdSwSKnaZ0j8uWxjlN0upNB3dtL76xOdL2EGwbZP8Bzcpf/WbV2nl7B
HOKB62KUtikZ2JGN/3GpNYXJvM6ReuvXlf5Eth5853CxUmVJmpPl+kmvNmT8vaba
vxJF2mWctPsTj6KRSyxZiGcLin8QeX7knEav3OiUH9MSEUJZZoe27uzn5ml+8mKC
HsRaLTBk6qt1u9Ct4NgaNFqanUvh3aqM/9xR7F72VocPuh6UbOkHVWYoZKmj6/j+
u6YvcN+U0L3a22KuOJ03GDr3Q0qdTUEmaANhjixrKZDfnf1ftRTDAZEfSCkJwBfL
ReXVppOBgXXdVezWlvCDjdGkmETJxKMm7T+8O0a0RWf063bxNVh2LQ9RoJVr7P4n
RIu+R46kEcpvMPOIiyRyvgVdvSd687Q0c/lgWYmBOMn9/DgpUbKKuPkl+zaFIvB2
825wnTdYaFqScVF9CbmTTUoD99K0iQVxEZ+cap4kA2DTeHOhq6HiFn4QyCVEBY3u
D0GWKgoJgrap9PikSXV51hIueRlSn8UEI++a3ogYNaCeMWr0DfK7mXadRxbG3EOs
0cMHWPUtJ4rqkw5psWzcvtsLmd6MK+MKGIm5U0hqb591JZjFJjkxmn201k51NkKd
S/UZkH8/ml0e5jXfB7fZQk1SMh09RKoeACPGInqbyZF+h0eZE7y5YE5f5w79htRj
49aHAsuSL6CMLy17kEgXorfUABrySUCgG/2FnRJGll40RMw+hNMwpgqKajffYSRf
AEVDA+FCWJnr8IUg2HXvGtMmFtYXP0i3yEc6Va8JSUvZfL2Lp2Iiw+9GYy9D9WQm
dhOSD7klB/IugjOdqHmJWu29+MwPPfKSHoOJJupdJHXlQN2kZM8K9/sPDnONlEAx
+KRuolnGBDzhfKhc8sMhWhTmcH624Zo+ssN41f7N2LifNAcNIlygSridxmSqluns
f3klONKJ3Tm8yfxX05IO8vK1Rx24S9LxtzKe+Hwl/UW6P0H3sZIr2+GyzKjgeqew
tXPbJC2VnXBgkcym3NyVaFzMDRcL2mYH3RYV6P5ZgdViLwHwWyTnf+0ZQInl6aOn
9VhgyBJzDTOsIPUOSWtS7RgXvjWLrzOxbk0fmMQMycUmIIFlmy1ecHXBIFKEyQuz
Dz6okZnQ0wra9/SzCTz0dik6fO1fOptk3XO/waP+rVC1ic9HHaScOLFpi75tG7F5
78TzPkPFYtVhz6XP0JJNsOOk0l1/64qP7q6X11nOQY0zyzXIPuP9y4WhQa0s9B40
rOsPooO0Eai2HfVXNjgsfkD7+37RvIqIkG+UbUtYL1gZyTKZYsAMNPtEjoYjsQ/D
MbSlSmJaMkqGMsm7rXkH5OGiS3RfCONegc4o+IZezmR18xq71e+GKc9HEmxiS89+
H6EJKVRgq7EIIjVRoP/zUQFEib3KrT8qu4N/da/9jZk+3tXV3jQRLkw7PMUafGfd
pOo9t32m8COsRf6VSfMrXUrEp8br3sfyaqos1fzVC+w4kaNNeTatFrxPSGuVoxFt
AYrZe+IH2ivmK3RDdBRMDDGdFdIXSALPQynJVjGMGZ4kgzv+41Q7hIkQ1BMVPRe4
r8Xw4it8VgqKEsXo0EVEG12sWAw7Yw0Y+yplbmPZTXo+f3CZLC1wuu+PvqyKKr2q
CGy1IHMKBjXDTLC1xa/FR8Hl3HNAXNCv62zbUsxP6sE+Eq9/HI210RMmGilC9uba
KurvqwV5BMUZReE7O7rgJwKaYQ2q37blQP60y8HRqLQngJyJ/7w3F0vAh28TB1x3
Coy1g8ZglcLBDU/4za7Zd4t/vPmMzyRK4YqAqh9KbyFyIDIX/lC4mXhLwoMX3nbU
3ZOkbjgLldlUkIwoN8a+fV7ndtl4qA+OCMRW1EiOT8dczZvsG0QzCeHFAQgTIZYx
MiFzC/LQH6yKqPbOGifUDVi6ja3pihynjqwJlz7sFw3z3g0ljqzXvlQvb8pYL0EJ
Przg/G39WsPtpODmgKnvhPuGbeqewAnT8KAYlI3KTGCoDYUJR0kQ0JgaguqayuDF
xankkGFrLVXQblSl86q89/WMgH1HE4XxYm3hH3ceW7Bd4RkomZeRS+6TDlmRZVzG
z2TE1jg1gQqbr3urLQkhacOxrQNCLVxNAuAN8UEyQgom9IaY03Ea3xK3LY7l1TM4
Ziq+uA0DwS3Kf1n68wXLF8HSOdP1rxDOBeyOeRiKZpVRiWEZ6HDWKrcnSuFV4Zq5
QYPqpbdvCYlLiRm4zMfKvSPCBDFeliCWfX96YOOFiXbC4OE6246IUOWH3gLIsiQl
G+N00vX2LaViRu4Hj4BV3pkjqLpXEvitP+fKEXNUcGUvOKB2kQPzfQLTdtDRTwSL
AZDEOczqw8DetLmnwp71SNFrxj9a0Rv9Es/xQgZgYCn47fShhmt57evNBg3ujXS/
dfylkdCHwCszOXRLm/Y98nm5sab4seJfD58sw20AJLc0eZ7D3L8Q3pPx1pwNNp2p
NPnVQ6ER8KDIjpaG3ZGfwFcMqz4f6/7f35H3JQBtGh4AzPwne/QFXnt1egdNEBmA
0bKenfEe/EFOMiaBlXks2a6BrxeuM2mxiU5C77aAs9jFt0LCwVZIDLsBnEilfMtA
PWBtqbF8a9FhCdq6r5KFAAQubgWTCtviZtzS9Z8TzPeA3rSY9KH4ezNeGtJwyIsL
06auHErIZcSD+Wyk8V+mgVfroC0vy37pvUm/CxEjUoKL9P0eI6V2dfB1W/BWXZjC
8c+oCUTXQOEBC00aNiquHSncrKrA5qRnopn7xn3pnWjICSselQBx4r1eYFkjBwId
IiNk4x4KOdwknZ6DiAGAu7W51OZrRPVliDnUUCe7gCDrt9RcRepOivSC201T9TEs
VbgeU24uSeicaAY2Th6FZqN21Hw7Tw4atZzKsV6ALAVgdgVhL+MYxnUy94+e7/hH
3wC5S5ps4SBdNhRj9YCjMhg7CB4iQC2KxD1uVtvw0863NrR2sh0YW52xMBRz1Wfl
aQdednnTNDipNx3XQF0b/FwHIcjNFl+v29WLpxDXol9Ou2J0YmX3tzUuowWyhkO5
t2830N2e/6wf0mELSfZ6OU+jiQOeJCP2ffwuPrtpG5maRID13/um7L/jdgcgOPNp
9P5gWkJ2WbHbv1ynBFlyIUoQsrAtJNq8cilmGICyThInBHyjKo3CUWQMbVMRJJ8+
+qINwgKzUWux2JNdG2sbZm+A7VBSkXb21NUZnqyxwPov0NxdG3AzEyor+QvhM5q+
Zc5GHNAdJ4G+PjDDwT6Z+HgZmoTK25OT/9JSmFIXwV/b5z+t42oBkCpa12QmqBBp
CcltFAuTWAdHvDf/tcDoRekywcaLLqVnnGS2KlpbdHtGRPjeX4sRHdpe5ag5hJ+X
R4x8YSVV2jGpHcBDRyhfIZtq+2aC2/fzxf9+bPpXvsF7jCGIvf6Rks6S9EshaGxj
e90/31EYwLKK+1htYVe/NjpGESHau191ofFo3jeIBxdqrUXQDypHVDKoOt+pHse2
P3+aY0AlGnQeT534CLbQXbCWBx9oElO7wXccnOe01M+4Ove8jb5AhE5fPCik98HC
xLWwScgNlmCfX9CiHVadSdT96n/U+h1KFnLziPzS7/qopTU22x+7UlOW5AoyCNo7
taV1XrMrUk+ZtLJetmxdenaHTNPRb7Nro8Z/ceLXS/krZw4hhp9/9p8x87S7hAP0
eyN4knzuH89qu8M1eqqZQA+a24mTiY3xDKSY22tgOJ1gVVKd3xOvXgS+5LzAq021
mRHG90OVNy6r0As/PCRE8cLNsCUr7GYenS7rGop/VZTNLFf7I6clKQ+brRBQN0LU
CXV49DyJ7eIME8TZKrlYflKN7N4Q5/pDH4qZCPbn69tbzvQ4tQo7idS+LarJQlQ6
y07bKMLVibmfsbKQCbdZ0XDnhBOub33/3s6TfwJJgBgfBbIR1zLJkxDbBytdJ7Jp
GBklhvfAY+/8+9TvfmN4IheLje8/YxuH5mLMrQAGTSqM5Y8tsNIyXH4sUyriVzK7
dD3s1EdawTOwNb69IG/x7GDcZHKKchtPn/D8YA3fC6dJRXvrobttJU8Qti+zAJ5c
ffUgDa7Hebv8U34Kgkza9wSRKW0lOtUUqW5JqcK9s/90HFYUKTWkWa08aAx7KRV2
5vAz4yOW5d7lGd0c8SY4e4kZrC+7FK4wY5Pj6P8eBgIEe0WmykgjondCh8e7pzKf
lgEZJzUPcbJ6EZ2gsYxjICox2qUEXXk7yWcgFusa6oZRtDhUcWC/fR+u8DlP5C8i
AW2vXkO+PdnyG1T5AKraJPbJ29ChDpptAFGCfbOIb2mpzMzboaXEC7tAXHv0wC4u
r2ft449B3duDU5yknFrdyN6sQ1P5ryb1a1qQAZDzG/tT0k8oGlRxAzwSlExwDi9N
MAXAQW7nWcq36lJdUGdCk9jgeE0UrtKvxKXb1yx51fCYiU3mSdCuun8m+uM709Xz
qvORUYyiD2PiwBCfSHSlIVEvf26f0nSpsYJLHlo9v9stE7fMOm2cWuMZyyZCXYbi
FWXPy+njr/soTHK8mVY1uo/Rije5I+AqP+uiBOekexLZbs3TW1hfuWbGBuHQcIKs
Lk4olwT4OHgi7iB73lfitIqLxddnRsySNi2UTzyTux09Bb89YP7h0SeCOMgopF9l
YXb6g2UYtOS0y39JFpznFpJttlU8/orw37YkJFHvXsQnDP3m2CNQjyF5HQiMjmWd
9Ghz9IDwmYDiQV/9esMiVC7iNxrom9MWoZ6iJEUMq8h/XioKzhSbkZ8Yi9RyF8Fx
FgoqclSj9xTge/Bgr8vxIPR/46XbgEH4E2XB8u26Pb3bXngXRnTxLu+KD0IqLajj
lpGksEH3NExLqSwMRwxtVEX434Ims/WUU2NdvwttnkZD/vfBdn/oKm7QoihClUgh
oX9AH0KJ/sfAqR/9kaSMSIckJN2hDrzLTZw8fEU/LuCeuiG/hDrz6NuuiVda+/yI
/LfGA/6DRcmXBsUYeGjEd+yz7IOUUDuIpJMJbTINOVKHErJ+h39VQJ97UdqEfzk5
jztVGgSsrkRCRbYNWghjBTCBb3uPeWFugUKiPhp5bAMpmrAeDT8IcQazNRua06vo
OzVk+5h8zOsZRI3WfdG3gzDdsq5ZMYn6xwigDbwws2B8jRa+OOx18NufJnkQ0w51
ZYXwEiBcJnQeVPn43o5yL/rUEBdkYcf/Dw32Lfs2g4HwhFtKM0ow6tgQeBTMuH+l
relGU8czXtD/Ts3PtJb6YEVF4jP8TgBqyji0E4NAU+yKEkcMxZKb0WZ3b+XNQ+YT
qxalRskHAEvngXVfwaw1W7yy5hv2M1790k1ZuS9SUhStQgJHgPhUvQcuQP8Xr+Es
vCi8QFWSNq343WFKol31CTskqne7e0DfMAo69swJAShHyOaWtFiVv/mdvEwLFOuo
wdEK6xF1Ukt+p3nfUrRCJMXsYo872HQxSvf3gYt6AgxxQ6FbVST3R7LtkBOtL9+w
2q67AkCEMTrTFlBiFK6hMwgPYBz5btxElEhq2I0cRNJKXSbiaZcoSGllVhtyCRRt
+jq0HxAv1DepDupBPFJAa5jVMfxcVyi/EOzBHkBAvWKkppEhBWpAw4z/b6GbDTHE
EoXsDHd8j+8PJfpqSOwH7fN3NKsvEVKo6rBb9K573r56xHcP9IuSY8VzGRiyNuZi
oVc8KG3pUy5X8yO7zTKI4RoIG61EUN//QH4vG5XQFAiyCg+P63XXh+uLpn0QF+MN
CNUSOw/X3r0xmBvySz3hBe6FReYJx3VqjGZzIvEirWfi1KwYcW9+2TxexHTBp7st
VCrYSUc3aMBoejLcxdzoUx61hsnTdINP12aJ2O7ci6XfLYPXf6iZf2OI1REZ0bXJ
cHVEL30TKbwW0AlpWpoiUGp0HUCpr3VeJbeH5IfDjNLroc229L22HgqUoJ8Jobz4
yMmjmb7JeaAougDWpwiufZFQIDpGqQrtDwVClNAWPwgdTukcYJXjova064yqBNty
6EmezcstHDOUOAW0jwbV2OuJZDKLwcCwYKpCwtM15Z8pp+1aEp4aF0th5f9aNrjY
WBtG5E36FM93tt8PKd9SWFoJ+d9V8oHlQqjhzM+fKbnx6WsrMDsMMk4Kxftjr+MQ
Sk1CA5yzOZ4q5zdvLu9/7rQcZswavxrVxNOexDLFKFJgfFt++Rp2n5zoha7tM+px
j+S9kJyiebCyWsCDpI2u4HQYR9foUe0ZA04M6y/cXnazs+arKp8CnW4nA8JR6n+O
7nIcTHrS7UB5iHrDHb/Pbg/0JcWAxpC8heJRMwC0WN1BCCWJa59Z/MQiZ/ED+yxF
CynyWkJKzVrPRWvvtbCMfYQSCplJ7bB5uvNffVYm1PDaxwGH9ZfI4hgXyq0R+DIb
V00cqkQpFZi/hXRtkTATVM5A2rSHmgDuXIGhvj+bEzw1EI72wUSxChf6V5NTFLV3
W8HthJL8NjTaa5MtRT35ya8UjPYRG/gUPY8YsQPA2andOeffcpPrTztvaNF2GM0x
o5tHihW6FBN2cEH4+konMfwAsvfWPSyD+exF2KryTSCMo2GPefSuzdeYYPIKs9yh
paJrpNPiD5h7eamoigwya8q9hGzlMkadz/Mk5DUcx4vMF8x9vFzAGIZlxKz6WJyX
4uLiPZH9qaRXdaRHtvEXvGVpFjbjKYKy+PZ38ujMrA0JhYuz+9fM8vA5oe4z00Ae
Z8V0x+SITrppfIm6Me7x815I6VQ011PmJs08D+eNbcUELiSbErsZviRu+gU5bALH
xEl+KINzBsnWLqqm4WNr6XC8clBQ5LprdtSs2NE79BcTf2UuNWm0PfxhcqQgHug+
/A+Mwrh+KqTONpiPMxCncIjx5jWl4sfPaUHQBUYkWpmZTJgCxPDwzuG/PQXHb329
AKK70vqS6VTEbDjqYfTp7eNk+enjuN+QWRKQTSjottrjqG3yQdcEMHHxhGM2wRbj
VsSrrGDVhrRGkcjVzQGZvc+OQn7ZQMLaJnnfTornl7cIk9D0mO1bVkqJVHSV1CQi
aVANhajBa0+sY2i/P2F/0M7wQy3cGUAOIJVr849xGsYAHHsOKJX09Gh3fUasEb0A
h2QCR+AL6fc+fuM+euJH29yIf44Rz3r3ZrtZqcVc4y80b15gp4z7oOYsz3m9+KVF
s+GOdXDeXnU7Xv+EeFlmLuSCc9g1Hq80EbkH0OZo6xtfJH2/EkhSA881GjCbvscc
lSnYP3hlBk63elZsjTUR69qBZaL6LM2+E31C8kHEfUPiL8t11gL7Miee+OMMIRg9
hgZm3tw/dxGl/3k6eWwBMEk55nE0+Nk/bEKGFJo74bo+kNOuUQzDiJdLmgFFpNGo
tVW0LjMk89VxzPyFAoIESOee9t4kvww4W09ZhtyFFwZyF+eeEvDkaMqgmIFvGq/7
WayMHWvJd65HRBYsB1iFrq4BrkXfHt6wx6Lpu0kp0coiKOqQkG7A0IzxMuyB1RTI
8QmE8zTXgiZf5JOa0QOF1qVClJuvGq03K1rb1Ue5ogTDV7V1ME2z5L6+lMUP0vqh
JwRkwgyBsKwE/zSu8Idk9Ht02kGjn/bVbH0WAJLUnKy2aypF5Rai/y47j5v/OrCh
OWk8ynN6ZhJXEncjrhRAgFhECF7zPcCxD+Mca0IaeFswwqEG6ljPwJ40Zv/9MZoN
8kpXQShsv3ujWbr6QQwBoZtXiCVKQob8mkp0DHsOpKfYjyg4LlT8laP4OysPL/qR
A9Dt4ylJqKL4sq89XmbPvhP6FyqGqHnOaKniIbKtKwIgS+DrWBMN4ewODp34lX8X
0IAif6a4azrq0OI8gk3fqOW8+GupaFQ5RtpGgf1+l/FQst9QDsFHEX+b7L0KJ+WK
UK118YB+8ELhr9QvM7FzahPgfjgw3Dq8jy6EQvcc5OfVU060m4vy0BpI0IKrTHXP
f4mhtpLz8b9JFG2GOzAERM5MZWWCUmZ80owFRA9yRgrUUVKzD9vyzqeCxbrkxSxc
mjmTPsO15pWMrZosi/vbSBk/BNoIbn6di3sH4gogOigK29SPyRGfnrXBu94RpUoE
FmUB+jb8+bUMeVKWwy7yNEXHecUHLUS1v7NIyARA85Xh01dDNV6KNqKOdqnr29LE
fJyRuxqd1cHBcW2LZLgod3uRwjlP62vDrCf+mVHPewXfMG59E3b8tPO/+tzgwFlW
8qZ7IMVrKAeShuJlB+bFLy5W9UUF/TjXfiOkCGxLIVUN6xF+Y3h3R1VmN3qJSRNd
YRkyN6yQBFnC7deNUU9qaMDPbMhMXcD+e7R0qSvbJnr3W1km1sIyh9h7VKkDPdzx
BVWAEizoo0/NJNxBHT7VM/gIfWlHcNMZZSODs4TKgyPT2t0sYl/c5rXBMn81UV/R
Fb1JKlI+nXGYQ5ZS2a9gW+eu5fH71zr2hSXvP+BiGD9kGB1d3mUEX8qYukwzhE5B
M0gebsRa2tNXyF3Ic0vynbwj8noQCpLQY3fSEV/fO74LGZ/IU0iHHZKJD9KVgeuW
sOImKVAkQRognqNISLT3JTSC7E3Q3yUlyJmZDnA5bAojfY3MtJPvBsGBJMZo5zds
9kdGUHHy2hJtame/U0xxDyRbF1m5cR4fxf4S7MITLkH4ETkesLqhM+3xSubQuwUQ
3LDDsN3UCmJxU8Me5k0YRVSwFx4IXC/kZyl76otbr/zosFWl8vYaKH4NAmfJUDm6
05CvaS8SDtTqVO5LXGSZ/M0NLfWiGv2zdg/sjENuulPg3tzf+ycg/pha/juDOv9e
KES8iYWEBY6t32rCvi9c3rOi0zBwFBox/a7EoapxLqvYWXwVXSrsBwk5++qYwkp9
d5k88q8Hd3/UZUDbfgB8hiESCJAGomiq9zo3yEGZiLNM8MCTGq+/UMdqTv+K5V7P
9uvaUsrf3Ypo7NtA5rbeGANsxkIVYUyy0pac7TsJ2WPTzjyawvg1yXtnYMQNVFir
GFT959oaHKwQhSH2il7qlkbwsdtzCy09HYXvc6rs0qELhDRMV3piMcRvmXt5lIjb
Ni3M9uGdjGNWsLJbLLNhQiMKaQz221g9iElXqxefPahX6ThpeGq0gCezwYwn/I1b
W+ExnfUPiTwuphPr9pcTdGDFmQ8cl5d+3q09dwIAn6JReugN/e7F8GkBvGLHEmjW
VTMlLqfVd4/NiOEAUPk+xyhNSM01c5Pb4IZpcFmbfKnpP0MYOYcB7B0tV50JaJp8
7ovYNZ1yV6UtDFfnxGWKJLImwhSuJB51uWolwqypYlJCYP9H482X4t3SWR/NmqE4
1xW5V7ae3STyEf3LPSoFZIMedQwQdnoX2NcUsJH5DK2Kykiu9R45tE2t6Kzm0ukx
9NY9p4yTNSOg15oaIW+lkBZia8efMKzHgZQYElM6B4nSmVq15ENHl5GGsxax7Ceq
v+lsEKJ52XbNc2ogx1Qh37rRPGPDo9ba/4C9pB77aWtRa1Z0pNqZTV92Xu7y+szk
IkS3TTfQMCGJnA5LE4oL/B2J2RiLSn5XmWoR2FWHnj4HxyJrLVAtlNovx2woke/m
OM1KVpK8PPWZF1USyVYW/psO1qNsGuwrzNqe7UlhSIwNmXcNBN4McCTdcGiRd9d7
MRM17+AiQIZvo4Wdgu2SmL4goKXETZ3KcmiE9hWCy/8yabxw07Wb7GXaNu5jB4rh
iVh+gBT8wLCg8nPtw+xhE8CUTM1Brj06m71lM8+y5zMqeJtOtPseuHZF1R8L/wjI
TPC2sPZCE/Z4ncJGsbo0rEzrITD/3lAgGd6l0O93vtqJg8kIe6on+BwSrOTvtlEU
uFva+2V7xLun6AbsBT7wGwiI5toTQrDl0q0CRWXGkidlRf8GKjP00Co9oPDdakCC
2u/+ZmOiSq+ZduVldyjpmKz2OOSII9k91B+M1+E7plXQlb0NWQViELeUsOi/hqln
+vF9icOTvu+jtc+W8NobU0IhWuAjP1GrB7hdojZY8xuF9Ynk57w8oM6PBLCtZgva
WjMGNRjPrs8jCKQj6fPYGa7NpbPrNtMWYZaVfGKzmBYGtg+j7b3DIpo91Hjforoz
aQRCNNTwqBAWZDv/6Z4zLV4yODh8hMM8fc8RWl8wz5Wm4vRT04bwOkZU8VHM7qDL
TYn3hYolp7VyJEpDibtO6TDs4BGweMb3ZDzNgr8GAOpxrh9WkkANXojNcEAZieTb
xxGFMUy0u9Xd2iF3zcbULM4ZNeakWyDe543p4glknK9j4ikQSLTg9cqqVxa4+lOK
9ygG+wo8lTrVkkgbM1OQvqhj7uAbcFU0+Q+LNZJ6UCdU9w8lnIn41SVzzN6Doudx
JOf0K0C/mFhYsnjFRQTPP/MC9oEiOrCCE76UOrim7o3flrWhawYgzN0qe/Tz1Fhs
JH1DC8fl6Z5biV8Y1zS8Ra3EbAYcQuXppnAGdC7yAWf1okibrYKxCPQsQ9UWNsE5
BONAKxCyZdf5xMQH64kYSoWVMAdOoOWzgQrlXvwWy1eo66w+/c3YjZg0YeBFhM7o
RBs+SYm8SGTu9VEj9qMKcFQdAt082hoRPq34Qf+PZFdplSizeZrPGng8UFvqzgIS
NOjQWdUFKDnVZwqE6CuKlZBdTLHiHVkiPfw/SjF61ffTFsYrZ1xGLtVRQ6nsgeJk
+RwBwaBprhmkvB7K7ggb9xC5c4g4uxA/pIlvsKSFxilfkmNkiSYrMdQ33xC93Dnz
uCtoEAk8etTao1hxXXRnqvql0DF3R6E0A08ubiXcdlKdlzm2TZjt2KN97aJvtika
+GsKacsimSubgVvjVTT6qCRvwJgAij8ON9BRQgWDIiVlhMuovapreSZIKUsVE8MJ
9/DqkMhtBYNseqXrO7bJKkXFhEja7lZysBSnzTNXPT9lU1MBDObN9KzuhpAhJYBs
0KCfSKp/gLZYxci0ufwHjqdveXnbWbi5zeqEnEcns38SoSSwebudhcmzdGGmFddC
D9Z3sWduFXqt1iKi+5qZdGOfsqTeW+lymMIl+mbGcuz2fGWTT7JP8oeo5AvVbRrQ
dBt1KGF+yUblT19AzpF2V5SG1gDQsCX5Ypxggj/Y/YfjtBTG6VCTTpfM7yxgxrc/
jhLld5SaY8IzCuD/xj9raBgRN1bcJCF3z5KYDUQzN+AS+OHOeN0oGN5TJIyaSWp2
ZQA9/NyDBKTqVUPKAxIoixO4Z02wJggBOR1sq0FAVQGSeNvkN/V3ZhTuunYRvKjV
E8xkSqhEsS8tOPfAIJ6Uu+Xnj1yszN2YOcWceKOwooXoGpxphJ3nPwXNTbkDZDfU
ARzlKuM1tPw4+njODOhwXDnae/v3bfzBrEAWNTBvYO8RpKYwo1XthZQMi6+jqx/y
PeSvEoRYbNVWTem64cgcosVSayot9vs04pBQk8LgvsSffERQ9BjUlIl0TlxVjDOd
pKQHcI7GeN43coJS9/nBefeDGPUz4ABfIa7LH7v4RKAsHZ9S/ew5qzmyY4xiGLSs
JQakPOyox+dLkyl4Deepp5IzOvoyRRKZJM1ej4Qe8Ju8Jm6hTlRVN40zIU0XcaQy
cLfeB7/SnsdijJ0/tCzr3AuHIYSayPVz2CnShSBOM3cP9GS4W6YMk4C07gICA1Uc
K7ZbixZ6FiZheY7QYxT77CT9tFkw9L4sISMj0narqGUrUR3tLAatgsUD5Abxpl3r
r97UK6ab71ioaDugDdKgrIITq1J3RX/w6DeZuOaBmAwUWxtkNBOO0uxHgMd/mXaz
d6sidN7wLnRLx/ySikE7vbRQWzFlp/D7w22VGx+OjodQM02bo9alTbD4oIiii/JN
B6vv+weH2RO/mdOIF3MCSTKhLyH+eEb/rPkMnyM0SqzIewpRhExnSNHiYptL+6TF
MsImOay6hcOAJCJvbYxuwal1ghNbaQ2w6ezzU5cjlvBR7rCVXR4CL4I67PyuLZK4
UJmaHqDVb7DA2N+WeFR8yQJ33H8MHSpvLcN01J90H9NK4+mcpIqYSCnAp9b2zKOg
2BmRemiqGG/Jlso8wkH2wxe/6TMGd9HEC3NQjUnZU4A8QZn4BSSAeAdw5VwmkUgq
VTd0Yzhvs4nM88om6ezTw2Ws46QorRZGN4XGiMS6WWbVyoktwp2i/6CsNcmLTiyC
MDj1ziRPJtQJYDPmu6Js2uQxFsuGSgIu01xhN/P9W3bjTmfg/mPtBi1+ot8kEewr
Iu8W0+EQhjBfWLhpqNhfAH5TjzsClLpl83WS+9MCMxzHP9F7aJ0X6Zv6QUIKT7BC
mtBqyUFI+RFmLc6oBAWrTbCFX+fxqSvWJNHSrgbOik5tcmGtJKix6Q7Cb7tYd4gr
zd/oXfpvFPKhOfaMJIy5mJ3fGPubcPMBXmDFUgqmv60VWUHrZ/WuXRPI0r4gGoLn
/I5nZJHRgAdpyuwIc/l3TlWKY/H9iL8Wf2NWx4ZoXx+GS6A9rVmIG9rddrbwVxKL
qKYQtY7WCIkjEBQpOM4jlIvPugSrSR/oculyRbsul3IsRG7UjfHdNIlrMWmKwD0r
CCp+woo7e8TaljWEBPyNpIfl34ztlhGeKSFaUYY3w/wfubU/vCDiJU3B+X8SE/tN
Y2y5ifoE0Q5Hj0JEfI2un7XiLlYk17J5BqenniOOptwsIKcAlo3TFkz3HjtWUB+a
8j4pM2pver1fut0xkZPWa1NH+GW8beD2KIPnJo/ntmGMvcK1S4dKzAByVQHlHTLE
ZEyPwIybRReGPmWfgLH0pZ8IEnEypS03/YzA/y7E0QqB7TUDAWSgFs/t8WGjM6g1
r4OqQ+Fx/7/c+eK0J86/nexlif+SeNj0EVJA8c43NAjphFxtHhkYiwEYwyTChQCy
kyo4DXEB3a2ljRIpNXZaBYfwgKc+Ys8KAe1cHd0VsWNZBTL86ul16f3AdvFG/Zky
dTJMnC4H5GXN4Imq44ZnbfWOA00PaYkY7YjMw7wFFdpfz9Eeg9xAcExFYppUPHrX
R/pg6jL+V6Jo8Fk6p3gqJItLZeFaeU8GLN3CP0tBPgijQ6MU0+mEgs3ML6kDyTRt
tNmiUmHYIWurO0lCFDMlZNoHaDBGwH++MZd3gf+vrVJg8HAzF09E3Bc4eoRvKRbO
EhiHHygchS+PLMj+ObLvWrmvNgWAjypuR74LkRW4uMvzriTL6w8aUc5IMp4ngTXi
w2wr7yAKor50CxQ0cCzkJPpLeTioeDCzb7qm8iPg4kJOSvW4OhowHNCGeV8xCY04
tb3v+GQzi9zUUDrzhX9TKG4IRoCgpYziGzx1Jw/ah+Gx/6/j4aeCd/dHICVDLY7D
JQrE18ca6PToFNR1dQQvTrW4OkayeruLStCheZy1VSYgYtBM5TSjcBHV4vHeWp2t
25vAh+WSfl9FqF8S/2VDauLqw1LrJamZGT6SaQsFAC+iu5RWlF+E1PCgv63nMmUd
9vBLQfZ3Be7ZTPM+QBXuiHz3zBVzEEcRdIDqjw57PnHvyTAOJIjMJ2CornFJqJQB
2UJ8xVLAMh7BvK9NqWzQEhqs/CdyRUo90hibIXFHXnZIXOLSJv5oeD3XgG3nVUZ2
qGHLUxEib50HDoScq/X3AgTQuumpn1jzVXivY2GXy0WAM794NjeHfai5hLsu+rw1
g/oc+OcKf2Mv4u63i1ZjAL+IJkL6M2hZwVuk95lsrMc+aAt2vLeNV0S9XJ9N+p9j
w5IPIxazoHeX7e/5ZCrcucSfZfLYsVn/W67qgZhieLKfGrN9n/9716fjDyZ1VMb3
VVrIbV9xiBpOLI76thJKn3zien7ejYUz80272OzBZPg1mWuH5fTcM/Y36aE4Gwqd
cl9grRnotalayvjKl85CRrdQXuhwMFwNKCv6nvDhd5MGXHWNn0J88LC1wVXmKGsj
NBe0H8XkvXW5tuLb4kTcpHuab06aE0Oc18EnFfWdUWXfx4b/P8LPG8sCOjGQ7qf3
buULxOYy55SlJuuOeQCaHD70c8m2DY5PP2Y9EPV45X3X1ceYQfdY8VnXplb2RvZM
tvs+aXo/MYULH8xdd8EQ/TXJhsn5RIAibhyY8+oSpvO5zagddxQrPmkJyRJusSr6
cYeMQsyxPWUAICGhcU/9RItVQ+QwOTHwf+AS4iiElz3V5urWrHFXXNiRujvc/Da6
DxPu714/fLxU61bjC5GnYcuuErA832YG9xg+NKAVkTnRWOX9/iJVyRWLymc60HYR
bamBXYd8mxogr+Jqv1XG+7fpZYz7pkOwV8Yk6uR/mLuqBrEdrZJYOSdMZyZT7cNW
K149WezoucfZaUgEEfL2L2OPUt9z6yBIYw0c4OePXeE9C5LybrW7a3zqM4Ev/6LB
buoyGcYt2XsrmXItBNZ09e+evpelyxhoEJxFwIorVh8X+0EVumAmT8fsNg0kP9zm
UXVbzX5SUmYwvEGw85PrvKlpXxxqc2xyKbB+uv9ikJwkrqkntv917fUgHezB8Iht
ORCgCLDOtNtjKznWi/0fAN2eHFU9jOS4w4lz/Pr7ir9kar5Lp4YH7ovlDoTAhuyK
okBsfpdJUtxs26EBd7DPkfuE1A53KlrQEQEm9yUSqn2sNYEEdIQ++xFu0Cu/Bn8z
DLvnaCMY/AnKiJBDCmIAKm5abU+1oekKPkxOzNfRcodXYVQETYWHZz0ikRR0L9uS
sIyNCQW5ZTlhdwgReI8/sZdLJCMXi9XmwvZhSuX92HGBynnR3/BJ4nwSPLWcDpWO
WPYob+ybkuI0rEVQvMHfjGTCPrAJH7O0CTtnMu2zfcpPyrKEZdPMEjhAWMIyUDlV
1SVJ8CDM+csybAXE3egD6iZIBUFoKL3+FvtfRhEfj3l8xiOw2uRGrgayOXXzmUiN
s/dLoTCPBunUtjWySwtt9PrT3vl/k9g761F2tKJXANi7e1cDC6KYEmupZSwbXPqA
hgs2nQRL7/NDAPAgYrTCmxHQsmzQo4cZFJivngZQbpyloUEP/3WrSCbTnVzJKq7m
ZOC4KOJssmkwKSSRXfnGwbVNtGNL7LYyDTCrFuuuQSMQthvgLH+JD3w6MHgjW43A
BQN4QXoBxA5P2lCJ7kIKPRPEPvrmdQYbOyPP5joQbjo5ClEvfumPN0cMYG42NoGl
Dc50f8hTJxPTnUVjAKa3soeufja67rlJFw8H1eeLFMCpdPIMA6SSCIAeRxgrKHFs
6VUIryIJCpT8Y2fqQXJCQy05tgx6rPviTGzq+Nnhd+p3Dl3ANPv4nMpuQ9PuZmIA
tSYY1lOYe9I+hWxdR9GhcQuPYGhuwbz1+RXRbiaTwPElXNUbVYxrpBtMeUKsFh4N
Fo9dayv3uVJS9KFn0xnwnt9mv0YgYDfnNWDxE/wCU1QjJmZlVzV8iNrWUuIgDwwW
hbTt17JdTZy7jL/kFWFeVIIqzwlYZJgu+cJfAGF60nOPKJs7ljcgfClXP5EmAYW+
fTMpHFw4GWyQ0cIqU0hWzWCv/qPFdzdxvPkvzZuhjrk6bPF3f5bo9U3Wff7HpJ0t
ezyR7huajLVvjxnhUOeFuJqqJ2BSmn8X28MAHRtXswgEeDhrQ7hNTDjuxC6tsXzr
gRxZMA2Y4wl/QieQ8Li4EuTULmFKDM3T1I0+kaZUUFNCjrGmEAZbypK522GnRa8W
8GsSo4Ddz4/YTAKfMBGGgZibUPVg0BEwjbR5SgFLW4+chxXr00nzhZ2Il8o6YdUc
sTYWRjge/fxMhyNSF0zet7TaklkJJzLosJoqcWa65+UK0wif8Xm7fgUUm3tzeiHf
EYUYrBdtMMyg2kH7jplI+GXat6e5mZYqz4BZEsNNSlilnFSfQFfpiHDOGNNX9X8C
ublCnESL8qpvoe3D34GiDGqoaXQOYLC+C3gJft0jAkpuxUP76nW4DzY27x+/l8Ws
mZllyUa60KoRput1EH7rg3tJxa9Eu+mPdRZUl9NoAhcH2yymKAdCZQuQ2ccST0rG
EsQp8UZFqfgvm2xqV6UomXLBsP2cD4uUXmyyIbInuDvuf1Ljc4dlOqP10k0/4eG9
NMUXuQx1sZDidJXqNmAmQKmVzOrsbtC0LV98Y0aAPe7TMy2XcGAjpvIOgm4SE+az
2rJjY1WSQt9AL6inlIGpesbtdwsCU+BkQ1sbxHUXATt11Gi80zCc1o30LKe6UHOD
u6fhIFrmG2yMopsxmt1QMGicvcghzlTE4gXCVspMZiUpip0PFt3N2W1ecY1nPjtB
mlWb3pYAXpszz1D6qzfhe9WaCktGu0seVNf3HBBx9wEDb83ckjdoOSd3xMzwTr7P
GNotY6Z/Dz8MQy1ORYeubmbudZ5EIz2CQPIG45dChHvpyjdPQRUrJhJ5iQLcZmhn
4joTzJQ8WNmssINXa0Ic4igG9cTQx7ltbK35vxiGanmhKSVB8DMLtrlnSIh8T6eF
//WZIaL69XCG+6QeTYSKz2pZ9FDj37eYc+2HdDiA7avbHhjzrRqbvMqq55aLWgN+
wHBMt3NflxGr5hhA/JgtF8e2TIyWAJu69AJUMZ8UJ2N+Or78CKiwb3KVAYcd3MbD
6fk38Of8XRh9GAEx8hVKlduGdJzn9DU7XWqDnq+fc0cBBVDFb+T5nSIkfvn0zaIO
0ZKYpaNW9N6X7bnjwABqpFOoMv7Wb60JG+8TBTdmjyS/Q0BJ5BJ5kdheyXqmS4RP
1mZ54Zy1vpBxTZ/B42ndag7LgMbvS5ydeLAdwvKXe90sZXzA3IdfpVf6pu5wXmT7
TuEsw6WSg/QUBYk8BxcUqzgjOeKBU1DLVgdgDsr6cRtvAzU5NnUf4lRdq1V7oEHW
oqpB/caKkuXjVTMJp86H/XvV6+QW4VujJBhu0a6vzThopVWWhsxAwQoSYhl+j8Mu
QEhCWdcJdLFm7ZWLZvkhNJbzFyslXHmIECbFd3ztdvOkrdmkZg+fKN/3Kny+aJWt
SA4HpDBL07w6+qOJjb7VYBRLmbpAMKEzL6tEHuyIHaPYo+4DnaEVyB18KN2nU8G7
CZh2ruSXZxXole+VWQ+onmkB0/XCidy6mztw6GczTPQba4zgzn8XPGND6E1fWSlb
2j0wutQ+WYzu0rAkkr8G7sXuNEpKRkVukc98entZHVSuW4LsyYrX7kg4IAwXEhmw
3tx3ut7JdE+7UFxobXk+Vx/V9esWvZNYBivH8YZivQ/OPFcpiXdIdYd58cQS1rB3
Wwc//LjqblK7/FSTyMu1Rmn8DPA5O16cqLEtO70En4G3AS3/3d2DGOwI9pvccxLy
q8RV4bYjoPFoinkmPUmALli94rT/mtnGzDNseFbwBE+OBCb6ZvLjEX+QsHZkQ9Ei
GfQHAbWn7VWtZKSjGjELpA5h0geRC6finJZXctAybn9ZlORoN6FxLuXuy6yrAPcR
kxQ+JcWcQrY7aNJ/vx8ybrKpL+Xhov/xNHTXcBChXRhJVIs0eEzabF0grXFOYjwV
IoGuFq9p6ncNq0cRmxmmsxSlSun9umUgBH6Mwy9MoENxooLRJk1yzCZlrJj+Ga5w
g4Jn9rh9Q1Lh4OzZSaT+vrKt9NE6MBMCo2zBxcYkcOAsdM2hdGRk7owLl6aYLv+h
Dz2RTdZyt4GWz1Tf6d7QzmGnlMJRBOAAmC3rP7sZOWqwtTXHlV4giHdaZTvr26Qu
JX4EldsU5hVzhUb2J6540Md0PCDA30Pn8qqa6U4MMjALnPHtjZLIRDBNE1bOkvOh
8BLeWIWTmL0FGzb5OqN59SXnHlZVGo1Z2rudMgNVlLDOqG8bHLD5SfF2lbh+Lg9a
gyYqVt1qr/eGXuR2RFr3GR5SorXETP/2jhe+VJqCXon9Kmb6KZFNGOib+S1oZ2dS
17V7qad/MmA1A3KR+guA/LJOd28mlIJ2P0WLTIajV0fZFkNZVrEbj5Iy/5vVFFBM
EwUxftL1xiwiY3iAUvckqQIRg6zyROKEikJPjAjLijGCzIZgtsNgxwEWbVRccBsd
xDSb1GenY4FkZXK2+X/9jCls9xcyguS6AplRnJ8+P/buuO1T8WpcSEolRaWK4uyp
HFsZGQ+ccA60srndZRWllEA5E5Nu/gWcaE0C4fpn16RlsEi6wVVnvRriBgUl/apb
HU4FxdtFDMRJ+PWqzrBxKtaXHsKq1sXOTjTAteSJvhhewQNVjbBDPIPTZYzMjF4t
STyuSvvZMCE3BMuHUF333moNMEqPDfUebsR4yyXCdun9jVZ4bvMhwd55kzyFP9Nv
m4nJGLD7THfx7va7YXWeJHzDa8COSK6APiFbTkKjsjGQwr1wgaUSPtAKveqXiVNf
jZWffuAz/3jGtqovUQX3rers+dJ2E5xzrngXy6xoaO3JaLGV+Xtn8JFtL3IYyWVQ
BM5tltEA88jsZj1/Fp8ZNkUkwrsHMrqrUkATcQLzXL0L9AIU8yvC/4RiPNMDOSQW
suBMXsRL0Lt7/V2J3oaF3I2lLpKU2v9sUiIR3Zwpd+ncaQ5eVudQtxyTJ23wUvgh
+e2N+MChe1XvcO1vemHF0i2ZGG3DOwo8CVVQeUoSjSv2imG5MQLxZ2mkrQyFY5t7
lXwTELKQ/zi2jaljl8PYxItmTKU7g55VElsldec3Ydad7UJnI1uaxiZPb8mjtpdQ
qKs3X699bXTNTSZY0avEo1jZqvMouIFH8VyDEw+MJ2XRY3rmmblT9Q358YWXAPdH
37YUVBX6kkOPJzkIYkNiLgH49no1qS9ym1Vtu3RnlycU/Hwt5aj8YQvAqJCHDbwA
14EZDvfLrxOe5asVA4w+MT3ri+tTxzuU0SwgD+/5XCSMx/RcqWOJxcuHzlhPD3ci
PXBQKft7jC6P4TthYv5vWThLVuqhR8crL6vSE37XA+2g8uKwBjEn8haMEtzHh7Ub
URZ4e1DXnnijEV+jmmS/Pwy3P4XGHuIOyr58gi8rD+NnrKkQMvoduulM27KyD85P
e8VTc0rgWg3OhkKnZ+rfd4vvQnIxhq5xm9PPhgJMwZjQsxIAp1kt8XDujWm8yN71
2s0BdyA6lOON8l8pUuaYritmjj2I2AVwbRdz4tNOPWN15RlR9fImY122uwt83Qom
QPodcWR85C0FfH/LliLN8k4r33jWpHpvSKvCD2hRsvAa/nIxznvnk7RIY8RXPhZi
x0B0FxPZclb/6Y2pNOXaeU4ywEnB2KkuyYcxgIoVYXzSYFMTN6uaT9VnAVzadGwX
4ZtzC5FM90F8BolgF/VcNW6oTE11pJEReiJxk60BxJWr/9dgsdsWxdk7GB9KLjJR
EqTv83AYw2r0rhpGGEt65GpNWxQ+xHnY65n7iQG+AYFvagN9YkxI7p6zFe1oKWGV
+dI628thDsIr+A/I59whK8nEQm9zLIh8QsdOT3LDzEZOwzxJHi8he4I1X/iHayAV
pwNrft4x9gsk4lKx+E3u6Fa1mZgNbgDtJNff6laVu+r56fGzsqR/BXykkzt3A/+a
Cv7EwJSVZKFQM17Z61PIkWaJDQxChwHvxQAUaG2Os0kdLfszM//gaXCCvW+Y6VAV
5HrXEJ/z02bdtWypyAGiIA8zElJVacW3yxtKksk8+04wrBiXhRrE2deaFgsGNcNk
wfSYiOoc/UyntH/Xa59c8rxNqQCX7LV+AeicqBOfcKYV492T7Mzdi725ehpXcRlB
+ymw0uMGk9ZxZArYqjv13J6tejajNZVFZZxNwKYoI7CIGJYxzJXHadWQJwMr9DLt
Enyngg7JwuE6xXMHAgMgDNyDwzV1ZE2pDJjC1HXXpCsbpdOtX6e+u6vsVUR4kXCy
9rwXFSrnm5kdz+16KEW9kAVa6nBKtS+qXeLjqR3NSKuCrG3AHfDFTHByKFSORdMU
0L5eR8jyBUj5CxxaT1Lo5H510jg2C8E5fFdv9eh4HuUOCwgAnvZjqNk1vG0uTyHt
hUBRbI1itmHl7Q6QAP5Td6FMfOItFxhNPlttUXfDoQzloO3nJ+uC5pRcy245YiRa
FE73L6LC8YDhrEL+54xXH59HwQyNfyrnEK0VOgHfZGTTGKcutFSm5IdPk+LfFUlq
zwbbDwGF/gcdfDiRpMJcAHeO85NNTAZ5H+731ZbRWi+aqXaRX6lOIwdt7YFXcjNY
zc5Exp5Nc8rbP1OC0TF+Pzl1KyL9/IQg8noTbisXyUVt0xFHLBWP/F4qp+zeGHaH
jh5seVphbFIP0MspFxW8/H0+aZZwTg3K9O/A313AXl9uRx8A7YhSKd7mR8eSvzhX
95wZlBZ4+1GNutsehu6ONVF79E4+au02ehYrlVBu+ADu1CaMklpD636HRXCbd5qh
QYmNxNQTj24giMM2mu93hDT8Rkbc6B0SZu5jIJ3XXkF60eSrXV09KCw1DXcbk6+y
h4qiFVNvAOOmlxcjWzrOCUybzaVFAhtInbbkMnLh60XKQvrB84Jp3ojyanW0O2+Q
f59os1pqXWLT1+L0yxpbzXi8DSb1HXJwGTePohXEX7XNVfKY1ijDsDDc/jxanHGC
5JALMxN4CdZVDIYdqThEz1mr14AiOj7vCohTouzyZNDIzN1NfO7FUuyzUbcLJsa0
0jZMF3bT4cbFC9slCOP9dFE/55rKdiu4xPYhDfLuy76hLQqjTa+N+uv+elbVYG2g
EoiyBAOCzy7Gf5kwPedfhrv1x1R5+AU7mlpx5vFIB8qOqmN7/JlcWJkjd18nCN27
6rGfBDfqqPiunV+tXxVzy/tUbNjwC5CVpnWpigdMpE0E5mQaB0PSRXacjf+NrkkD
FqUG2kx85A3M8ddl2bMR1avg+aZgSSK1Q08EO3CTdhLxLh3XSPNBXWD+hyjK6EPy
0R1U3bs2nxVVGO+GootOoPHK78PRoKgabhPyfaSqnnA/fWuikZtdgjRJv3ePOb3t
wVJ4W1eYm7qE1ZeRIBD2EF1duixw0kCA9ILfdJrlXDlKP6KNLjEf29kvLau5Tbgv
YX6/XxtCTb8DYKAIVNp/DoSEL3jCfLZXYVwcAc1o2X25rpZtefUZ7SOKhPoGNHt9
xMTP8Sbp6AyQI3mM23h05GgxLsT/wsm4Y7sXrIztSvsnW2PGzrGJUZ2Jdp9dhAk/
CqInKq9ebkflpDc37/pLK/hhP3WvdhHT92gLR1GMty2Yn2g8Kn0mlk4VoTnWJ60s
md/pgCnRj68YyEv5o9evnmXOM2T9BA2ZuhAhkHb75Qo7FJS5raxZ8ZL0TknQEE/T
QQJPxggUe41/RMnQJDeEAQlSAZYLLqy6oA6seDYEsE4Tx3ue9zQk7KT9ETtP6cfg
zICNo0V2Velln4WY6o51GQrODWEhz11NfLh73sa1yqeMSPaIqWFwHxBwPaFbWKxn
wSAKrHzgV1TZmVpnTJFhCqSUQ7FfXQys+euslqJoVLvGnwZ9A7pzqZQeu0JaJsB7
JMF1e2/Vjh/5yk3MiKB1E4mgjRV7dlSVp6GtD5YaiIBPY8WONNhhzUz7V0pYDjM0
SmWrjfYkKa3/cVlh8yuJu6VfHjWf7hWV8H13T+bjWB/4TG5kP3wcrNj0PZzGBdaB
BZGROK0scW2qgWGBzbaGGzOf1ylRw2ERem+LIcH2zkJWGaVVY2TWdcsLn5wIdNym
As++2XULjfLUlD2frJXtll7Preugnc2q1Llr6DYk0KkTg3FFx9Yl+HWoF0cSCy6h
+aswNyjhY3s39vgcZLOXgHTQFoLI+cAkOejyc0wKQ11oyuS2I/9qwlaLYxT3L9GL
Q6bloO5KaaHjkTxF6zA/T0TF9IEjJU6x1J+jUU4AvPZHqExxgDPJXF/FJhdq9CFb
FSZ/wP7dWNAIxsYwIw7br2usJ7w2JDvGvw30A1qqzgDQuytpu8ox3u6bl80v9ye6
PIKPdNsPGTLi3taJh+lNDdg1feg0Ybvraj6rMktf7wwbhlUmQhBH60i7/yAuMfs2
p6wxS7Dz16Qe28wrBbCvubEGgsxmLrO4Bk78iqIqzB4iE3XGokflfLbFRURtZCRr
7Hx0r9hkMG3NCZLR0wpYzSDdiR0dvT8ExJvVxiAgeU7u2WsoNyQwM/vCr7jwdXPu
iokvBrM2Thqyzz5V0stUH1L618aDAQyb1HOK/XpuuvR6XbIuDbTmFE9n4g10UIqp
fUehL5ktFbLtvgZ8RgWyYjvRn+CUWdxmLWWBa/hXHcWN7swK0JiOohG8FXeV5u83
hyEE7i49LWNvUVaEeWheqmWZ1xoU61smiPOIFOKkEXv+FXGvcFcDvz31cpZ6g1F1
IRJRFZuyR7vFfyFIv0CckaFRbai0ZH5BQGOVdqkAxwzF2aSzMUfYL39GPk4sIi6u
W4I4Mg6JwGhVR3doZo3Se5rfK5h9ik1nMdnQhVL1gzpxMRp+vs/ZZB1JGXYUhfNq
wuwSp7B8j5JVgM+vjqtEZ82i40dNZPlYHcmGHqwSr2vzn0IDDU8E5x3LKtVY6B1I
TugJNmwIxV1aliMJrghJ6QnMR9l9ofVTdgeHe3dS6ERn1fO8ck5m05OGJPYfwNa8
6HVNjSSwP3vp99odh2ZGgl4z6SafjKjvRM58bq1w7azN5rXUSXtD2Up669jowmnw
4No0o63dFJpOXnAbepZ4rtta4TLe/dPkA8/hbhVTWAnhflZdXtO7LSKjqXA+2DwE
vi+PqWzSqLW5g0IxaqVV18P4eexce1nxaVkb8+iZPpT12QTC0lTdDEsK44Ht4avw
WTGS60IuaxJaIXo2A7pEzhaca82M6RQdGAriohfGzSPaaZp++QwCJxl2KAg9w1tO
x6fNvOM0WhuHq9R5G+ObKtaML5NjF8UfmEZKoCfK68TaI9RQ1QSqhu+m0F/kqjza
WmV+NRh1IK/gW3J5Z9dKBU1mvku0/TArcwgOsGqUS8BIVV6X2n+nI+XBtm62WN0/
nwN2mJvyxVxc6Xb1Sb7zXAIW2kkrSC7s55RnwOyGis4VSVrq6HshtZ0qJJW7W3OY
n2N7QJREI3QbX9TRFey8vWRvGTuNnz74Iz1n7WKljGY6/G2bafUZiSgSr20Bf3Pw
iOXS6gkhqgDbJNjBxg8gfocYmhu9e7W79kf3oADtS/1O0Itb1CH1P5p4nL1/jHO7
dWXjU1Zue+Xz2073VU6dYDneA8t0OK0/8BCqIGXe6LIHXfnvL2lpflFcXikmIo5+
0boeFc2/0EPh5qVaknyR2JnqQ7ONf/v6TNl6+sBndW/yJdP3Ijstn4QFAROGi2n6
CpHYgzZMTnYBFrXOkGOrB5IP/ggPntxCXx+yY5vOk0ykd3yjKfbLeOEDfgPbjDN7
NqC82zmtVeBuOxCI01OjoJ4GHEOJ10TOaL7Kp0NLgUfH72jMqC2/soCro+YV5D7p
bXzdfQoS8UQdxMJcE7XFj6DVQqP7nMI5cY4Au9qjRZWFFusbW2RuvdfrJ3FWsaD1
awp4DyYTnSESgJ+VjE/yatpyEFQk/cldZrh1c+88xiceaYuoe4s7PgBwWqAHRTqB
1TP35IAHSZKEOB6iwhQ8H6Xwgh2gFJfEDPFksKnyCdZFGLZmH0VMKtBtkMhLuFYC
OzPHEkRfghtbY/E7axXHQVJfgSzAx64P4yVBjudNCi+DQKHSLVaGghinS6+8e4M2
nfGbQwrvGt7qc+WjLxU+Kb4Mezh5xYKpTWSN4WvOEkbl6LG3tU8f/OaLJxd8fMZk
221bk+rshitbTADD25pNyptznbXa976XPsi1GyFrP6CDsmhuJBTJoQ2Zpg88ohQ7
k+oXUZVG/BDfT2hZfP5N72oK4AS0ZPU4ntbYkIujL/JorQWV3z+bPBGdHLfPcvOa
zN+SvzU0qdODM11bvimOXdUlEleBl5gnwrx7UT+N88X4uXDuEAntYoAbdNVGcSok
+UQN7UKn595T5KYBnSZagyCDI/7EoGFDmGYQRIDAEWtCltFgozcmED0FcWw/CTTU
foUudfgyJy+PHGTXY9W4SQsY9ZjRc1RQ5ittJa1yq1ZC9OKNGa7O0+bHdxqilRRy
EVxFE68AkpaJSK4t4Y8M0kZzpFbt78LTAlVdVk5/fu5i+TEWjdHb51emRHHKZ25C
jrAFpkk4y+uE8V1ImTs4ZyQZTIUK7AWWgEbSaYIgvzOc/G9F/HrFBrCNdVkCOf8+
67E1w0qFSlnZZ05IH8t8nChnK0nrpUpI93O3FW6w716MBW0SnPQZJqGzqwJbNZKD
3U6F8vjTv5TTpS1u9N2w9tZJug8vilaX3I74TMSHSeR4rbF4elK7Nj1/SGaMPAQA
IYonQ8/HIT0P2kveTMUpOj/SF91EgpCDLEld6kpiAWorHoJy5sbtrfwFtHdVUr8D
uwz7Y18vPaoIXXbIgyFy5ROtKF2/E0rsSPQSManlIVOpNB1OuxrmGwGbR9GUiWTs
ssfdJGYPtjnMyVeFwGfaINDXG8OPC2ZyLp0IrJA+3lyJl6qH91cFiOsiXGQyBPfk
+ZlHkaXCOsw8ER5gkOmoVFrE4U7ZiSf3z/khZBC2DiYFXDRG8ruP8ZlXeKo/kj0A
55apw2rOMI2rAwg6YpRdq3qc+kNUqv3crlcotrAMsOjv6+g8IolH0CP4WLtXGzEo
9X8aHKoWeow85X7OnPGjcw==
`pragma protect end_protected
