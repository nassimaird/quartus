`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OY6oraMkOWZYo0ciuPHFU2XJpxJ9Nm3ERfkX0pRsKMmE0uLsdSK7QmWh/R65yKgy
E9rdmxIILnfOkAOmZs8nE+tIrR1ZB2LpesA8SblXGp60awZT0fI1BZXYSOUcC2dQ
tmsr+qIz1PY7P/bzWvFI0Y1YBzEGFrEtXb2kVRy50qU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7680)
Jm5MxNAanNVMYhkEnpWHMZXzIAzMUtKwhjceH4fgDMKV48/mvjIZjwhh74qD30Ph
Qw+FMHK1aw0mCXIFqQ15e0ODiMQp5FRF7LFO+eV7SRGNOqa6oD9159zzRWXQLs/y
fKroJIOAHecA/G2DOCAFQj/z/fiTweKeTgO5NS1eae0rc0qTqcby9wf7GtRE48sn
GqSSf6k2xSc1N6qO9KP4r8RHi+flOod2h+04tQnb2967Xm/e+cWmTG87QxZOgmI2
2UA/tD/LNuZUJx3UC/wMiUnWOQKZdIa7bf5PC7SW7ZT5JGCxB/w1OcVjGa7feeCw
74+bB+cMOZtDmpF/VHsd5EhPhJ3WpHmmNbEOHTf+F7r43z9DAxaVd3ozSySA79Yw
1UhM8M5qboe66YSSjlQlbk0s9o6W5ItblwJWGQFhTYH4bMOk9Qo6u1C3KRyFNzLe
R3v85mQkH/ijjhUuOp3SLDJ/ShorqAsTFGR12z9MZ3DJCY2zmdkDnEDLiRc/tVIw
Zg/sS3VL7kUS1ZVeuWZpwtxHUi5nxUdS1KfA34OX7DusLcyI8lyA931quBynRpde
0QdVScMf7OJq1RuGWi5BU7kw+zE+SFGwH6YIwitpjsw54s6Wt1al0nlJE0THluMh
9XG1dSigjsvvxo7WaEyvXdb4x78wuz+QaADhWASk4hvKwG5vLoWdpdVH1PezYWMQ
a7RzmWSnr0G/U1v6v6nsSP8i6jc/ArsUVqoRj/YQMYNS+/DBozUhcrUkjH6US/xC
b269SfMc1B95p5sWu2RCEZU8rZLdcnTAir705k3bjyRcnzTvkns3ZEP/Xs8+JNow
WcNqY3Y0h3kkg2wykfBB7tzzSoUc7dr/EPAqRKIEjuskKy5oWW//Lzv1kapUb0AP
e8Mf7XWf5U8X7M5KFnw/w2PZaiKdd5kcJ9SyteWybjamLH2KOaJ0koLgVwz5dNMs
JwYXL6ok5arNL9CpznGYXeDJyGmLhplmEhm2OZZLN1H4P42r0210gp541CH5ohQo
PT+Kol6lmotLCy12nAMC+ZP7PLBZ9cdjeufGbV2k84TcDMtO1CpHi5R616ZggHC7
7FChcAb+ArzfxhV1TX67h+DHOjUDDs5b2YX4JrI8NHoaRxR2LNqYE2wb7SDE16vP
V8kwODQ4IllDXGnfJoZrxPOZmo5i8pIMd9X3JmsQceOUZPNwgJ3D/RxrQYjWBn27
9aeM+M+rWlNiCbAvXHy05UOBJj8tFB+rTPydazj2pEbwKkG8bsDm3n98ApFwu/Nw
7lOIJtOhOzmEQZgnOU60uQENsmFwV15BMMM7Wfjz4qSWK/KKZZ7UMg77DylVDr23
bYh0fmR9rn4OhaAA7jdb8DPBBjDvlo7OicgDX4sAslga7YVxByQPY43tIEDUf1ja
jqkU8+MMeBCOzD/P6+G4jAwZqXYnm7+KqgB4gOne+GUSSW8vNdE+STqCZaFTTc6U
s0D3/m38mFtLfdqUwoi8PfuwgljIf9+5R5NOsjDphC6XzZNBE6lRVGT0oW7zIKDB
kjL/KLsPNFG0W7PsnLs0dp3eamGeEGssiwO28Wb4OO3UZIU57K6l9Dk2o/5HmZEA
yZhgn+/1fVD7JtaGeD5Ew4HpTRi6qYxAANPIeuq7ANb28Qr7S+mGc076yEBziwiD
Em0HOTTec+GkmuJU9jGgQSkQ05MrZGwG5tCvDTNo06njwuRNNAn0IS+8+9OREc3E
S3x2b02BSVd0b6t4/HUoLexFzVbHN9sUU5RKpPgRcDE33uW5KeNfaIXwxuAQWxlL
of+6kIFESdOooiT5GfBB9Ujtpo2U7Ooh/7q2Cd0tiwYc9wyknLz9G6MnYoiXAuC9
yplbvyk7c38RAaqRV9xg/RXCvyFbrHtEsZp+I1SFwuyWVkReyR7o9ESqLyBFkf/j
yoVQAVWCHidceDnuF9X7txpJ7hhQajfzUDbSWbeQ5ih8AS440kCYm0bS2xx1VCXd
UrXRAEZvW9kmUN4DhgDG0SAlTw4sd1PbhDPvIUu46Uc/XvVyEHe6Z37NUkgqDZbA
fHWJVSTUaDLFX+W5h6VrnEPWGTWMlJxHlaoX4cNVVc4sg96L0X++EthwgQMBn0vi
Ohg09qPOVfbGS0kL8cQq3ScmWKIONt55Nll09eompUMAih4hkIho6VQEDM/KmiTy
okNe4BFjNqUTNB9a+115gTbR2q5ViQShwdrycj6CYOpHO4JY+Lw1ScWN3PeYi6ux
7Y0hAZWan9lRiLVQgGdjGt7djPKPg+ps830rlyKiHOaF7yHd7ip8I+AoMlkrPFcS
jso0iXmb4MQoFPXqWU/7MuOiLdtBnuYplkRyezuECARCQvCCt+Yp97VI5IdkM6sO
5hvmobghir2CbEbfz0cxV4FDp5kHv8Vo6HSnZtjgJGjuIUB36ER8ef69I0VzgCqz
7g0k1LYjj3BPhfajzeBoHbPcfXxsDLW+zq1yruzn6smtoURSaEwlb7zXC8JxZCbp
QKuSmGR7sQ+7/A5dDAzDvX46YL8mcb3c7r6XhmzpiQQL0wTgfUhsUFrw9sjw8k5U
dxWoT2QdH2SMc9hGuio5Piknwb23+hszngOCa0xhB8V3q7UwYsTcC5CZyI9wRw2+
u7mAedXz6/8K9ZEncSH7YOr+DTaLaFrdUrXvrKqleVsiAYR0G8q5EF9L4tQE0X9O
csMPM60AWOJm2kxh3jltxbpXuort2D6YTp82asGS0KR/ynKNYRWfez+obgnE5DH9
0LgZY2GHAZPro4kjhGXPIUju4ENQldLkM0QWQhcAhgWEQ2oAihXOl18KjiuWDp2f
IOETt1UdchxAD99VIjkGGd5m4L9ZXx8AtAsK0P3MOOFzf5ukw/aEMMYAE1BS4tDP
aemv4BaE9Z/QYg5gHEM2+JzNVh/1VQ/Uk8vLt0361Ojf4XtYWQI9r2hwKFQvlHVu
frV63ZJ4GvesgnL+bgR/JpAA0meXZAie5ZkFFiM2pI/IhNBBe5wRaKXe1uEOkMEV
jtnvtLYM2JBJ9EzU4gvw1JqQFGIQcUaidUuF/GkZ0prVDEdthEfZM/HG+k9WKvsU
0uZ26hhoQce0NBtCA4eLNpKm3QgX5OCb7C4J5e0RrLDgtlwgFZIHfChltBQkT8bZ
6388qAaMXw1rMWgP57FxEA18odVYRa9zTUe+FMxeMDHk55ZnfE2hylU/CKmPYRrj
7J24Ddu1JXbWxiTGkcwANGEbBVGPVdmxkpGcshBknSqCdmzaEVeX4IzTZEPyae3p
lFbLduRjV6Ye1q4CpbzOd35uADauOPqOoxN6QolWceO+vp8Yi17qimPdaTTB0XIE
SjR6SYJ/pdPd9aiBS31sQAtPBxplJjl8ALUMBF3tWoqDqigSkY3oF9OZia+N9xd4
KTlduMF5XBKPaPY2Yz7C19u9vsI8jfrbw2Cx5FpCHYlCjRIIxFsVec5Y5xOZ7jR2
AtNnJ0QDsEm7fkiqwsTY33QqjREsKjMiJfpRWvnJvcBxV+A8Bf7i26gY6vbjycNc
Yk8AONZdJrvf8dRJMmwXGT/khz757HhgBWgkx7vYaaLYl6q6+WG3rK6/AeiGpZyi
DJ/UlDIX5LHpNtsNlNPHLshXNkmHqQlW5O8aUtcn4fgEmZWZhlWHvz4SfL1+5nvj
A64f5/5S7+VoHdl09QEDWYWhjlIrLCaLPawV3brdJ5Xa5jwmnp29hnDiDl6+nK79
7vG2bj48ZCLgCjYvNg1wMagK7VDuM0GcB3HDRzRSfrWQpL9165COhXsnhW/w3NK8
tSKHff8BovI2ojdYA9ZtwrVpzaoMYiKm1l60dLM18BlKOxlT940E0CREYf71dZ5S
tT4ph6P9ks068DvGhDlmLtc6jdcp1S3rCoFHtwzVLH0ErG0qTz8/UAyBZgj8x7+w
X1mGRfXshV/ov+K71S5XaFajoH6Dh6DcNlbNXWPccl0rAEBG49muKCRA64SO5Aak
BvBd9F/zJ273MkqxySLvuZd7Nyq7G9tos9nJfu8XNbyNmMbLHFdSieTekTWZ8XKI
ivAbmwx4r2A7U2RUjo6PAgZj5VOAWQEAjJnFb2P8yt3B7Zj1m/n7d0gMrcLgIfRI
QH8Ec78DEj6vtD7l7NKw/aMZVSm+BDEfW0TEWdLLxoJ9YQqTvZ3L9KVXr/rVZJA+
zR1oWfAqFpbFG3m/rBFL/eJzCVY0SWk10TywZiaNNFpQETtTJfGGCJku1C+K3Hse
Mpuy6O0MOPts49P/hgVv/eWxUr3KMeljkbZtDBla083F3z8mWLDQUSNB0MksBoNc
sJB1DJ93ZO+d4ApmiUCFTE1olhpko9zS1FeSfxqpMhhcz4klrvOut/6hVH+hV1fq
n0zNL9CYzktm3oUxe8wfFD5KZ998AyT8CCVv/5+/UAZTjHMEySCJynZtiOwyTnR8
MYvt+1X4Yji8zrAQWDVMkckCHId/qL5yNvWMc44Jd3xl42yemam5L7Cw1EGlTdcW
29+vu590dY0NPRM0e2qmnYxELky5fQvTWliH6FiTZrboZueOVzSlmSqInyxdtl7R
3+jiCZdafLBu9bJSjDop4tBN+8/QKAfaLTWVW557xZYrmfOnrwQMxyv1ueCocRXa
zHmMf9lwf4YmDLnstkuZcOTIoYCxI2415bvUcsLCyqYNX5wCPN6+r0H/pai0Yjdx
P3L6ryFkMVaBnkSFxqJ3HPBg/Re4WxwzJUa3W/3Dlu/yzSCPO0m5C9d+ysrZ1m81
1AamibKFApj7mSvunFL1hsKM32gDpMRmImXuKtoX5bEfwj1iWoGGE1DXHeABdZ30
YeGAiTjCqiExi/12AZxi+gy8UJYh/NJmoBB5IGlfVTJd055G2eVGPM/OxCjzCZR1
UzsVAAQJUWK8Z3/4cztmE/tD+8q+EK4DOd5kxSfxC/kUL54pJS9zTy2qoeUNH6Vw
aQy6Fs3slZZg7YzzzVoJrXLrSJ/xbu/ppmqZJPMfdUhP0bGEN5PO2BE9NTwXS7UD
JwGSImgMarS7zp9xMZL57M6GOxzLOZxexUiiLh4CuJCumjLay4sjPlUWYWKnIpMP
FwiR8zHfchV94dpe+xyQVeW48rd5ayq1B1L1V0PxpWUSkhQsH0yLa2gCuoYXIFq7
/3LDsEDBSbNLB2joqZv5c9F5bnUwQl5WaqmAnMyPiRm7Bc6nylPlSQiKRpe7ev8F
QmDcGvBIWfq31ilXJps+5pAHH8hNpGFOhMeYQuj64/IvfFc4WZ/wdEX6R1BZ+HOk
iQLLz3+iizAjJY/bRxk5ArtCKwM4a2v1cZ+z/ZBT2f1isF1FUC7Akz+kdgwDQYZN
ahrh2W/9zweBLz/N4PDDam9jdNgByGm4616XZK6xK6PpXHXKTbW3NKGUo93C82T7
o19n/Sd90YDaPwXBT8Fct2Wyc0mueoEYwr5zvNRVcSAU/s29fLmysYKADrzK5cmQ
wHgg9uzNB4UgsXl+OuPYUzZq4QMH05x9B2iUi0QG8gh8S7OX0U73jFtlCcx+wI1Z
99k9Zrdwx9Mpm8H7QGKiq5XpXYEpWbWcfdUohkQgu1xuTcMLMHxUOzPA2OsPf5U7
xjzD1AkpG21BQiSvKVbyfIAVzJ16i5KVrZxc5tGBNQCKzj2B/bbUQqI8zM4a+XLd
44KEwxxeQQAcvhClE+FMr8ogfaD2Zo7cTaFMvJ3wEewAS0Mjrhenr0H97BW2K02Z
vZCD4tWgNDyZocTvPk6dB8PSNXdcdM80+z8ZyxRNm/MF/Z9n6HR+dOLkbpZThhbV
p9ljebrJ2u7tKcVnDQKDJeplwqlAO73El7OyLF0S2TSM3B3DtyWImq/KMxxTzoB7
J4gHPanh58UxGgG53fnZygWwXkG/ETJB8VA3zIVDFFpbku+kx/QO391b7DFq9UL4
ZzftAthc8iIo7FIgCOUDzSk+RiEofyBcT7N/0tt+RYUblPhaCIi12bWcB61KBWcb
NELJ+lU7k3loAkV1nD6TpzXr2P5CsYZ7dVrG+t9+DjGmD8JT0ym96tBXM48K0bbL
Hfpp8CL4wqHIjSpEcwZGoFlK+mdRvGwBWmLwA62oD1o7sgo1DO8YroG2fIbQUfx5
c9Dpjdzd0Byi0A727Nwt86EZbRgOyK/bdbhznTmQ+ojzTUD2AHWy8/ONShZkgTKE
fPXFEYOfCY7qI94bsj8Adat54HYNHobAQ6betKsxa9Wm3lFhE470RIQfIr79+ad6
oRq52uKIaSbTgZQJHvEmW8Eyefi519fh3z+xvaqmgMdQ2+psEkaZRkTwuWN463TP
Hf9XtmEVYv7thuhXrBC2IeHrhH6N7W8xOiLQ+GDP9Gq9MFV+Folxmw03SVTJRzZa
psBVyg2P+woYeAUgaGDyZH0eGYJ1TWW0q6UN0qeKq1kI6iYJRAH+gpUcQlcGYP1W
gzvY4sMH6lTEWCA/gVTVLhRCagEFsIS+aLzKe0H8ppcovv5wikOtnSKAs5nSmaCz
mxkbYBSrhZbfut11AMnk1iUYy4TIk4Yd97ZQ+k4NDqDsshbj5+YexHHG7Jf7+vxJ
0ol3Lm6xMnHy4YR9tfb83+V2fe/rCcJGxoauK4CDdEgrABFmtW0gl8lJhIaxkhIz
orlO7bJh1hiHzCO9Hk3Jkbd+Nxo0/fdjbZV7L11Bb/M873Sis04wbLBJYA6y86d1
msNLAoih/0X8W5enxoVZaqg6p8Youq0dgRWTjUjRXgKEsi64nFSAPH+RAdcxubvb
i6frn5Tp9ShQpdT3YnQHH9DErviwROf2RCm9gMZ4MHaMUwKIJVkHEEQzYAya8xi4
oiTVioYeGMPxX5Hv0loC2rhq1gpdWg323+Z9SgMncXoyzj03wzVj9yUqmZC5+HQl
IPxOvThkopHHMOlse/DfpJ+E3+TTVX/92NV7cLe3mPb2F8nkEXUgMWF0zAlDSLHR
+RI+VZxuiO+ccGzHZwNezQyssVJ10g/D9dHo+KrcsHN09jggy6LTogrxjMFN5mV0
2lJE2t6nT5+nGJbhY0IevA6qA0N5PcRv56MclF5xfXQ2N01OIDi6ZSdzcAM+PQ5z
9Ck5Gc6EitJt9ZIkGSg58QbMYFMdk33e1NpiCRtzdRCWYBaw5bkukuviqXR1XFsJ
EhGqwnCnidYPRhVXEuDfqhPzyNuY1n7zq56IE63Jd/T/x4jfVaBXdRSdCLzFTHye
rxZntjH+y2Mz6lC9x7n+Lw1B4JKYh89ZzPyWA0K7R+zhsuFpgGEzF2ciqofWgln6
2OOPbzy0e+O5hwKhyypCNyH+H6a3cbCYkMKiaQWuB2VRg+qM+SK3Md7hSwzZbU/o
Q83kS1XgwBJxbCrzQ7e5ZLC6afko/8UX+3lW8sOQ3PobQM6j3mokIv4mZO373Hzi
soL48wjodFYKMPcPxkAIDYAY3EVXIoYIfkF8tbSpkV0ut28PqYqxXkC7w9vwE+b1
3NuhX9XvlKiXxgg/xLBthB3dMdhagoAGm6cG/tcqAVL642bK3hptMO7huZXXc/kN
DBPML3FuzIaQalrLSkhnvssMzJV1gC4T0NJDcTtHJjiwswjyteVtf2DrV4jDU6MH
jFWf1QlG0UzVhTgfrsHb4SBbef+a+caPm78UKHVt6UVU6K/yfAR1C9S/i+LUSeV3
UmOEbcxyvcey/PkNbHMb4ZL50d8CajyrPOTHmdel2ljTAHpdlzG7Zlr4uzpZTPEp
cMD8lh4Jbwz/nNgu2KU/pRCC669bkH/gqat52j/4bKO2SwBalDsBUrgTcpS81T/b
xHV8H8WL43QsVlduCpF7EN8AasSL90TNx9Xyw6rj/9Dc1NrA4a3Um6fZCZ4KRipZ
Od068uZxvwRQ2oKmKwuLDO7NNM5LCSO5N1gP0YfOIRKxVXJFE347s9TEAcvRmG9c
sJ6/4g6j2yDyZAtwM2IMoZ9xdmNwxNg01SttEBGlX9PILtLCrFwgnsfO81N+vVX6
kAx1H/AiTXhEuoUmZF2NuXkOklcGZXjyM27c2xtEZxR4ajLb0dny8i7/tRfsqraC
rIqsavZu+ML0IvG+eZ5e1hhOfQVpepuThL7giCX63ZgRCxJ8YkmEoVYO8Gf6N9L9
/G1G3fYULYCGwu4dDNW6QHOOxKg2HOJvA+Cgnv0XBdXYjynYi1GS/JWH3EvSCqZ9
rlxrdeX+S9K/rg23KbcF+WLwvT3TP0hL5FFbO0BuiUL9Kt4wIxtGWcR0f/tRUYPP
vLkk6Td47TnNjtK+1TAvn6xHdumPzE+w9XhpT6T69N+FoEuVZxj/Pr7Kl2h2rgp2
Xs352mbIlaoLxtyLFGh/LcHMBMrIiMCVifsZNXnjOPckJNipusx5/YU7/XosCtLG
7bokurbtWwKpuBHnvJjBVAmKc49Cmv6n9z6J84tTcsq+MrPl7asOF9A7nhldFhI4
KEIK0Jk3fQpCLALdQlZ/BbyV681tMhSBcbc+lpNit3kgzfiDa3RSttDvCSXPEzqi
U6qtvUn2TyuyyY2s9JCDz9F+laB2jyNV8cXDalZL4U9O7BNccz/0AOX5c6W2Lj4w
q+6TYBeZGIhNcIVj2RnvWqo78KXsialCTWsi7xNLh7BzZpAQBLi9fyGiFmpAJuvp
2WOtguM+AqWQ96AVEQH2gT/zcGPky+Wm89TkjLP8y3Hm5Zdp5dHOT7phzFSX4osI
gRSUq5lyg0B8UCt4FpG4uLLgRQNI6M9orn81ZmtPFhoTpX9gzQ4GrLnljvad0jVn
+4OyFtouW3/BnRCOIR8ClJdXDRWDpKzkTDx8ks5DO5fWU5FzXyNcS91NNsVX/Vqq
21QCAqyhssVloNF8HQnv+cY7tEG/EkwVitzYh5Zh4/0MaP11sDQMPRM0VTZIK+XY
8Ce7a1wrLiyLLXNNAK0qO0ttuwfHgjy+JNrIhRYskbPdO0p73fQtpvYsEXvBETqX
2zvKroDRQoxb8bHtOlftFGLahMvQ+a2eV+IlISpYQhBQqmxqOSGMwb9M3kLKYZ1r
TVwlp2VLKkgM+DSU87rm4rWM4EJSzSf0D6Q51vqSiLDcyp9GZjNDP268i7Mo86mn
LhY6J1R+mJ6xs+FV3Dorr8iuYcgXLiNwOLGR2KY02us+VgQ+O1yBpVUAxpYRKeb5
83V+w7G2JXJXaM05UPZCLt7cBAGTpP/uunSC7vsNxNybp7tRof54pYhtl91hNYY4
0iFSFhXxsWDgYeEy02s5+Kb1UM5u2JszApzs5T5prXpaBO3D+cy7fG96KJLIHlbc
R73LS89aDipztJcHaD0HuAa6KjMOU3GUhjl7vcyjs/Gy1qxxT3i+F4CSnw8226No
hVpRVMXPVeQEIJq1JsS69UFCLZdtORq82cJHH+8OpqOQLfwTfGTQ7AtGgpVekAxg
vaAJUCnXfsnTsdRIt73FzjPlLGY8mKL5t3UdgJiymIvlvahNZu8x3lWZBcffm1hJ
H5amVuXZ9uxRMXy3VE2inJ4udGUCaT+rhq56SE63vJLS0eijuBpY6728oiDLirqk
JMO7Oratf0ZHfelDmCTWm3JWx6XBua++9rn1Is8d+x/wgTjg6x5HzfXm2Ef/pD5y
G1WvCYOXnrQFQJdvLvl5fZFnd8hk+gMjdujAQNSrf33AUCxGCXlkAVtNHxJgUlB4
RrrlaLv4SHmrYjDsD4rJW1o7F5CHvM7rfKGSx18R+oJKJ29garhrdbF7umpa+r9Y
OxhOf8X5Xvvz4tAj80jXBW0E/cB+5Zt2QeVIMi9Xa2XTNk7j2SxDGgA/Tm8WwCDC
xP4tmU6l8LLuQ4GK3YwiL4JrNuHDRshWDvKkd9HrFwpSmoNRGOiQAVCjB1BUhJnl
qW0eMoPCAFY5qmLwV4wSANGC+Tj9UsYq0Ndp1TV1zIMEw1Lthow2pJsu5sSWxDFo
OOLVUAb9E78UMbJ5ppXBG4BuTI0rggweH7hHsbogxxuo0ZSyF11dXmyAlBsBaewW
LXh/HbP69MmIOa6n7nXvZFMIDnZunvvj31Xm1ayLOgU0DutuN3b02CH98EwJlE45
l6vy+xxi3Ino1AyvbuokftcdZOiYeQAfiRM3VZzFEF7n72zyaIOiQOFJ04TdBnJ1
omlRcyJCGxBHhkNIqN0PQe8cx5WDMIubux8YclTqVc+BbF4rSlfD0Cxt5Q6x4m+g
Zs23PjI2TnaAT5zdj3i4GoPztrQtzKUemQiBOzd2v4yLeCjK2hqYoQGgcYVJt+Qc
AncGjcDVFVFWmfuDAVVLgdaJdIuFPWhyS4Fp1Z4ujGFdvl3UcPCy2JVwWWhkZJBl
`pragma protect end_protected
