// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZqvSfOj9Ukmklw1Z7o38+oD9U1r3KXNGZ1eoLjfM/r2cq3puJwF8NMzuKKesL2auMhCKPkV6YPWN
s3p+sFuYrKhTGej065tAqFnR2/lNFft72yw89yDg4AGv9IV/MKMT9Q5ruSOFr81sq5NCaRpIziy6
Fjx6SIxEfp+B9/qa2nwbhjQ3oiO+cPpFJ7BGa3WDdifx+nDEEjTgS4eCnCrMapBI1QaIErOThKuC
VwKastW3cg6bfxU4XOWdHCgCyo1+DbAI9RBNy1WR6aDxYPVjcRWkmxwNg0ny/6Hft5/0E7CG8uYi
q3/wvj4zH9B3p5UEXR8RSpxJhscqg7XZxqGBPw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15504)
SLDheabrI7QzniZglyzfkF6ZSKVzFTwisUWfKbf74IDWx/7sN19jQQBeqTXSWF5zsT9+7nCIser5
emqqaPcJ7dm6lbzHFVRrtxUvXFVjyqrDGqjI4gC9SFMZEy/wAdhhy1UjSd0Wd8rLqOxAx8ep0BwJ
SUGxpK1LzbsC0piyHjHhPJXOe7lrQSiQ9IvC7HQcd6rH0NMQI5PeSYk1T3gQb1vm+sFnpq1rZhyG
ym0twNfsZVx0OK/YariK0HLnOz6un9hsFCPQgq+Zm1pjBj87TZ0/njsR2tVMkNXSrg8x88R8Wixe
QZtiju60qZfgxljl4yDfWbNNMANFOaAM36OoERYaVctcXEM0brBpQl1XB+EJo1evA6+nJoYwT3lm
LGKCAWSkPZvbHYt0yi3htMX7IsQ2wpSzazaN7BE9Nz3pvTC3G1CnyYLiBQI7ThQ/EuiUvK4mQ4VI
QA+9qDdk7QwvnApNgnbjhEPo6UINz7jRe7TKojbEZLwwvJcY0maBPOIGIJ0oTT3n6Ivy0+Nf5bsZ
sXvA4UEXt8rX2l3g0ioI/2Ke86LVtNiG7wnAf9rvi4y6U38GDWzFP/js1uPXTxvYMRSsj59dAPFm
QTDVKbUI6KGb9v1UzFGG8nPJtc2yAMyH3zChBsqchceSwfceWcUISpSaQVH5Vf5Ajx8DdTXinrGt
BSeqpJhSgkYj/3VkIh+pqCmWsIH5Bc8L0K7+Joc3pWvwy2547xhwqKpV82Fv3kkm3ajLmy+JfPFo
iY1P0RhVYycyEPjHr3egZMHnpffog0B/T0tx6e1q5V3LfUJdjpw/ZsNUeHmJ9QHVFWxPwG9iTsmL
RHbB1XYlzvR4eyZLUEOqwjn12Px9wyLm8ETtSoplV58XmcaGC6nl/xkJyHhUoQMZszGtD155/3wz
qeP+eZhptwKP9OSctDZP/n6rfboE1k6bUewnzidw76urmbEsrLYHIdly1bCiLve3TOaJtuNiR4H2
0tVTeBprDr8QA5mwNBKQTdbSF6GiysXqCm3yAZBe2izsvDGEJ7b2F6v11j/CIGTG31NLVMBpnMaP
o1q2Jn12ejVAEedrVLGfu1UvvgGft4QQye641nqSnAM/tppfFojmQIpFNZ2o60p9HTnuT1gM24E1
OAkK4dMNdAA+QQ5+F9t6qF6L9OGzcQoScE2tYtWp9m7e9XH3TfvkVUIo3G//D75j73tvqQqjuEVC
ecVpo2h1Ebt9VgStgqfyUfEJNfRgrMOv7T/fWtFM5Sx5gMabaGmn8rKcUEWPL+szm2RFY47kHl2K
n2yLEuJFAVEcVzRLMQkH3UkcWhDIfG8OTAF7o6z9QrSxeiDMuBDbRmmQfRjeUEBGWhn7ZWDZT4Eq
eg+tBUDU3cAIBH+F65d6LErn6jJiFVALbWPQWzTg0K5nFyZwncQN5q2gqDDpMz2HR2dScpe8wSwb
SB6GM2Y0i5atYrg7Z3frLuyuMpEQV8lO+83/PKBPOS+56y3B0aMaGNhaLFL0qOU/Kqt4VweoqeYO
o8CqeebyfV25GdhHRfGf39vosDma2qHB2ZlL/Qu3ybOxxrSvgwJXzJP+jmEibwIh/2kdCmDUgHik
TFeSRkp1YJ3yDB0R6EakIKt+kmb9t0LVMkz9oUCd8VJ+LhkQJcxGxJjM1YuAbi1fd9O7eFzIM3Se
EwfBgZHnij3LGjYKHC7V5eG66Uac6OSHtHC44W24U69wjN9203/HJy6rtCom/LSisJHVvCw5oZnU
NVnYwkGXeAuk+GWBYjeHyMSgDg0F8z95zPYsXfnZvIHjNlRvZhE7Jq9HpcjBQeZ78kK7fqL93yWB
/FEj5A8hXXZNYiItw37iTwcb+mgu5jbgXBgGyUneV7u6k5nU8gS9NoqqTJ4iByTQehppavx9sGiV
JugJRq8tHrD9mzB4SEWiNC/FuPWejaFh4gHj4xwziipPLLpZhkThGelgFnQrXe/ol426kzJ93yEc
u/92H6XjxZlSsk4ZLeBB4JiaIylxQY/lCmAthhI2IJkxgcRwQudy+ZU/TaU71PgcQU+r1aGgLlWV
snzRJcnLNyTO12wRTQ35ty2CaUSSWJjY55BLNtlKayVpu6y4bUcllZ7kSJb3HmhxYdN/+n1Ap+RX
5xkMVx0RFbsysT/OPwO5KX8E1VSE/CZitZ+8zJdZg/dPC6KcoKvX0p8LZKGMhLRBqEpPcekY8s9C
Ts4UEN+ccQbFXLlTgMQczTL8pJ1mIgW1A6rz5pJ3nSj3RUQJcDY7gbWFnI3uzhprkFuhe5owJ0hm
C5IvF9k5iI9Fn6TDOxXbquF/jb7Xgq+M0toYnzUZHuUwVJg9k8HdgpOe78uAj0bsTfoj7zHllT9f
dyQK9bQovBxn5CR5HVFMlICScZh8RJJ5659c35Q4yjkbzpdstk7iRdnVmpvz6du1zird9KqFUL8C
Nq7EHZkExrfhZlrpUWk7dS7Kx8YrKwfwwGedj2efNGrfnh0MLW1B6dCnGWZ0S2aLgjpjz+KGunR0
zpdyqpdGXCm9vAc3cIFUB/er/CASo7V8C/9fs4soBAxTaK1IhX3tMuX8uw6TZGglqI5YrXSuQoAL
eg0+hqGKeqgjRxFehkN7wxHVXiy4XsRjQgM5Q2G1vvnHDfIjVwJqMSbFqUlecQsDrPIWv+rVtfxx
ke0bd2sLl6rBtho37mvMKplush3Y3gWNCG+1Vn2UDFDyRcLyJoTpbw4RMVqPUYLFHFQ4kUlf+eSC
lQv5wNLUepwOvm/HeUBGk+cbkYoDDAFdQG8iylFmrAmQKj4lPaSlUMUpOOIFHw2TG5nARik0iyo5
k6Jo1gGT7rWLA/z/f8hiyoKBRUHqIFYtXD1Jb96A0aMgQayNxxww0iPeIIT77D7HQtV5ecN2cIh1
l7UYGpxZpTDud0bPgZgSWvTlyBDmdg7aDfNHUwPWL2+Pjs+moll/5/ghivHWw9zljCWAX5tq6tv2
8pMz2qFachWLRp1pu+3d4P5gvDKleiX52FhPTuQwytwn/ESS4YxsBSS14NL+Gw29s2mfamdgGt2C
SR33NE0OYKuzj+1X3Sikd6NOkR9YRrzSXZsEhosJZ2c4u33VycELuragLzMkAs+nQ0HvtjO0ms/i
jJFHWBYEyRAfJ7z4EwIGaxTYuKtPR/LEabXCMBrAfV2Mn7/VzZ6CQSuaNM0Zz7MTkzP5TbDF4OiX
SryPRpwpDWOLWix70RctpN5CZXtNGd9TZTbvi/aBNNsdRwYXkSZU2LEECn5nALVx7M053G35sio1
y1V9ZL+pP9eThmd6bDSgdRXxIHad5Ye0/6zrpZTQdy4+x3YMTiV18V1LIsfvkoaWp0LuFI79r0EJ
NAIOKssvqlVJIzHFW6cjXLdS4UTJ2aJbY4087mwGlZ4iszmm54NwqezeWkfI1Wb7ojntbRZ4qLs/
qu5yehxIFmxbtbJgxmKO1Kl+1Z4NvGS+SGH9NBhXzjxLWcDPqVA/waoPam7PPOSAN26fYQalBitj
mNJwUqmzEZrQHsj70Z9xP5fcG5XtpFY/HKsEFFNzE1yWT+efA9maSZObWzxeqnnXWGC+z5Fg9IlR
0th43/6hJWqz9+1t890gjBRQAR666Simv9ggSYadShBYHKX5R35cv/eqHl2gFHOjHGZGLrk20CqZ
L6y/IkBxgQp8IUIAnVKza4WBTnsBq8amJelTDfZHBvtVQnihpKOkpRvi/CyOdLbZYumnv6M2Zd5k
SS6Mg0Vio9wSz1dNItxEgxZPs5mQw8ZWpD9y49zmaCGl6leRqaUs1Jp0dc5PD1nlsnsvuoCLHu6D
NkBIHADcvmvcS5dWCSmb7f8By46sWwF8DE7VTW9y6oI2lhmlMJQ2/1v4kvNMM9shP+ms99Dd8VMy
4qDFEc6Bfcue7OMsEPo7RLxDoDhAvc/DdRhieuNVMOIt9BAwh1LYzHns18QuZavPqR4XTuDhKB3k
WpSIESpOriDBWWzXKXY6NP05tag9GWXkIjateOld6kqanC/A+fXG4sx6Cm/xC3p4QbqdOsERGzFU
WMo6ral1CQCalZimBP6lqoUGkjydQoqlh+/5kHcOUm5f+Te5b3smKSci7pcba60j3A5Tkb4ZkhK+
UnsoLbSJA4PPFkrUj2ws3RtZGg5OHmGsJtdBd3r4cNQP8V+dlbN9EQc2vubi3Mk0OygCdjir1vYS
gmusx05OUUljeMvuj+SoFLGJxiSYSpRuhZ+qSLva2yL24vm5DFz5G2qGMWNk+qJ02aZopyGB7VHR
Kapkewz2I0ivwYNTY1ObGhrfOwYGzJfrkrLLBBLaXIKWof5bbU35aW0oq8Bux6trVgliNntkhu5C
7HdCPLjZPJ+ymthWLnbxJ3ch0iXIzR6Y7x8wUwkqT4BzEMeoiSY6oPob3Qj45RPnAG8g0InyOUau
TarZleD1FeaTEMjQ06cfK/+Dp49BUU9xv8xxw50ZNUm3/Y0f/WQILuPpHCobhh/oF8r7v+sOCsnH
nnhMYoEhgHMk4YYQCXOmDOKeaCxQLECY8Prubp0RX8l72167n+htkePihsEfSpC3NXJ2n0Zg9pdi
MToQXN03q1XIfAiv0WV1Izv8NiV2zqHZvcOGbBIJEGE3yxmStVMbSHKbwTWjZLu3sH7k2w0pkG3v
uJVpaNXPyZhPGYucNrlprpRoA8inHYuShAR7O6FyTT+Pwfx/DLNaPmlK27cJWflgMJG/ZpLNGFUa
bHDz7mUl1tm0U+SFz4s5yyULnYEDBj27mdMruZW5gpMUq8vKu6wczaz9p5tIXAQZhKt7exZgu4/v
JbuHo+j2JQVLu3YrRAH5QO/a0UEevjlq+TigltvXS9y6rKpQi7mPoEJrKglU64BrG9zSiZvMP0+P
/rh6Ari6kIDoU+x+mp7HeoD1fg3XMpJinbadyaJ58OL4seLrDGoyneZ96mBCNlqE3plPKGqM7BRq
Odl6uveKdMtyfFqOyIS46h3MSL2R5eAFEz9Y2MwdeCRu8QdEqXc/59gv5T8VAhKG7/0PW3Ipx58I
cuHtV6NU92IBr+daLHiF3nEstum0xA3Qyk1QYuB2Zr7u231JCIGDUjUYacLZKREJApeQeS9K2igx
P3Lo5MIkgY/qNWRgbktl5p081WWN5UCE63aD7bXtFZmgRMqHpBAcyVVt691HZhIJCGiHUigXUQAv
N+gY1BJIRF2np8FTZ1EmaaCosS5f3jPiDzyKzDc7S52z4bxyVKF+KmTel/kBv6hkQ7hRYnRl3bNg
R5A46jc7sldWlCxui5lziq59o73KHr4zCGtbcGcW3jIqBLzozr6FkDvIfhlEBuN520Ch+Ei0gpU1
VwZ8LNxWuobHbvwGjsl9tWdFL7HbXHQw2L3ubTYlnM2LCbqrdacaGJKLU1yDBE4mXaAjbHNQCHsY
Vt7k1iSTevwqKSY6qm507HqWNcxuaMG9+33I94vGaaigSSdt6kWxMRE2L0NH5QlsyeKLdr8Ql9LL
maEDzU80SshpV21FVDhvDMtHvK6Mr67SWYcMM6PI2J7t2eCOGatDCUo4cHnMndiyVVvC+rZbp6bp
wKm/JvRdxmhSMkAlFv9I7fCVT3XHbuHwswMqEFfLQwlUw7QnFowYbcx9PaZHXI/co25fhLR8fu/Y
6ZEtEAHovJ6lMvSxBPnIV5RGM13PUCi6cobZfGnwUCVIiG2U4g3dZMvXw4WRYvkWw06wXbI05Bw+
bygRkncrp8MBkQQ+iu5R9m1jClvD0cJIuyxiCmCmWOjeT9f0WauYkKs5J1/juoJhwkWr3HEcezaZ
JjBlvqC6S+w0cv1F1YA/DWLc+tMUx/Jbfnano+fr2wuICSFkpluvlt2AYn9OFTi1TcNaEQcmKfLI
djKIL5hMvV06o8OSmYiFjGgxcKWARXxVN6wFYCxy1jYnACxOEg7XcvW8n8SJJeUCJZfonjt2pmpU
0Eu6PRbfs9xywO5fXNTkWDhuZLPHdkZYVPrFoT4i7ZjdOW6gHOfnYH3N8CQ9vpxM0Yqs7DgbaPHn
P9JBkus/IeQ+yef0Mk5uGyApyKRIFmxlAuiPmFlbtdy4F8xJSyMZrH7EUF7hkFloBHAlVzJprq64
6I+6RpQbuWjZZRqruXXOoGEg2hYSD7EdZ/i76fAzsNIdGHBu63rcjp+acE/cn9pd5oGNyzDUQkVK
DBpBJExONTlXJYt3vNzDt37B6LX8bFJJlk56I6mV9MgHMzT7uBdSdt4IUsFpsKNM70TxCGVAHio0
omOJrVwFGEWYMLkxaZcNYPb98RgDxsTYajTQLVVaK+2YCr/KHuBNA7J9LAFlXibIf24EzdWPTtv5
6nx/wyIZsfjS0/W0IBCqsKH5201ictSpu0RT72d8fyhrFsJAuz3ItAsRcSHM/7v18tKck8NLzw77
+1SYDCM2fXc0cKGQhDn2uu/geu/O/0PZJ6tMeUgX6ZYmxIB7V/fWvxWcBd4HzOUbmVCJp7up6Nq5
+NqTpyXg19jeM9c5R1Zjk47BFNRVH+RcGS/3LDGw1SsjY+Cg3f8gB//ge6H39LiWpLsDTWtXkjMf
SXoZwxKGlZs0p+HE5xw+8/0j8qQWzFmLLgQsUBsAeqvxZ1iVoXY/XvN8epLKtJPPicpiY5/6Q5k3
NxgdpMQFZKeGZ73tVfyLDIRkiFrPGbmGq0lcaoY18yIqEqdStRZP4ipKMEAo8KMI+euGvaMau5Mg
5eybC3ooA7f1QUkajwnjfXpz7jZLwACpapHUGGz+9giKbNZsVuYP160XCBR+x1iXyju2eIdcZVcn
zr2tBIkj7Exs6u9NyZHBndn8o51LnVdI4U4m+So3HRjXT79+TRJtLfc6jbMq65wK0qu8zcnQkamx
siLkSxOZY2PmJd/lI1v7UlAUSwgqC1+wzvuJhspbYCHAu3iLRWZPURokX2zSAyR3ERhJ+vdKDCoL
ofsxFjUuIG3JxWqBeeMInSdt2x0QtAwlNBdFxVSGmgagijhHwPKQFejldEytjGOMvfVDhQ7fL6kt
scRexFuhO2uzV6lpN93rVDLdCgOL8iCX407B/UenQRqxNpA93ryVZMAr3ZKiiSxLigLBTteBtbxd
8GqfmaOcS7+mMND6zD8VksDjHi2NbIlkdnbLqkvI+iFYMqNN+j5k2L+PUB354aFKRaHnJ4HeTdEF
qBPSAp2F/zfYCGqQkpcFG5Q4kn6qa4qCjJlE4JZjTz/vdHnfP0VaqPQgITL9qCD0B/iN5TiO3QBf
LNTBZnRhZQNqfJOS7K9CHfIVVPyb5oMH4yKF78sy0d0QOoY3uD6yY7zdze8Mo+ufjBEJCv/ASsqT
hAaLw4pR8nz9j3sYl8NpRaV60sUktc6NxLjsHtXdNNxCMk1Z4rjp4x62YHM5poItT2lg2wDqvjpc
n/laico7Sj77a3Y8Cs030KgoOU31uDjD/u+A6DgcITgZa+cuMpnJ/iWd7fpAA6mM3kRT4fuuoxb6
e58HV3vfghBBB3ECyK2vDh2do2ep89SiiSZs+q7eWcK7a9hTnbyifreoICSg+1U/Ynzc8ezxfO3p
oA5O9yeuO2AWBKCCWRJI1jVNE5iI7OZIQyN2ZyQhq4H79+L9cUN3Q8iMS8v1LLLAyrU374RPBM3o
Bjeon/8oHYHGdQUsRD/hCc1KnjP+lykNaqRPuRpR5CkZMNYTB/sZpVqc1vIsN4O0oLQYtgp9KsSN
3iiMhKx0vT8NEIywyU4TV6G2CqCL8q8PQVgRotauAB9RiVQ34EOEOPORBXrluYU9K2T0Kfl/nA4Z
/9QOq67sBeWzGlzD9s18zla+fHUjLbx9k1PDeLnFfwlyZH37sA5tuca6DhWv+UILgT9Kvi1jpaG8
2H4RGxkFnNGzaZ7HT4pltzvgi8LOBSqk9rR37Zwv61rdKekhx9Ov7VT3ApjPXg2DvH45nbBezCsU
AknrIs9gDSyS706do4RRcLbTVbTzb0Livigprc8GmfH+8bthaAvXq0sl1i/pl8UtQPpZelTEt1z7
r6oJRY1g8t5zYfg9kuDpecVf+72lL6GTjVa7fyNDW0qzS2RT4tx4vqDw18LGErw8GO+pTf4Z8no6
3v+OSRXA6KxhI1XspjbbcRxYjTyZ6Rf34dLMbuO3DmtNMSzgsk6y9Q7X1jjUkT8iZgibFpBEzZIk
nWyAj0CsNKpqwizMQjThm2yFfrVApUg3bkHGJdTExVBTgzurObM5btK4Oh/DsQtD1yY+KX8J3Ka3
jzadqvxKGYeZnC9ZDQGeQkJbOHEre9PLGwO6JPWNYENIrXx1cb4May9fQpDdRHhuGsuKxqgR80H3
BK/bGbKy3RIxrU3wUKnPV7sAGK6bBQTVJB0MX5dNI4GMEXnHNFv3fd0luYdxNEaCeGo3nPVsb850
hhqXO3HPhMuqYIGCVKivc6EGjKn78yccDSdp4QLzke2W4x2JTJvlqsqvTeyqkQrbEX/kK0Uc0kpA
37KVs6VymDdvq81CnCeAHpShDKAllZ3qCWB2bBhDe9Mvs2ClFXTGdXzsYhPhONxqHP3EKxtRwODt
Ojc7txCj7KwPfkdi/v7DXH2hw0BhymcFxW5ur2RdWdbGI52V5rEi4ctLyb/nkn+afFgeX6FpWqOk
jzdt1/W+AgaUQyPHMbtJVIA1QDPc+7sQ2MiCdh78PvYAa2D+FD67rGJQKdKbMmCM0ComP74A04DK
VgsRxqB5ZBXCsPwlI883/Rv/rq7qMIlq85dmSYXQsheFc7RzUVd6dBBJ9Q6y3JhUcMBWBMllp1iG
6ftcpMHWj7WFx3XNvDSE/HwZbfBREILB4iRI9LVAlPvlB0U2frJGfC4Df+Tp5TEzEyBtFtoZWn5u
0Ttp80pf19PL43C+3l8BJHUVCEpdfeU2E1b2QSS8NI+kLKwgHzpK1uC3XVUXV0g5HS0swJq6UJ9e
c2WN0pMxOVXR1S+1lW/+h0uly1dSG5+IXy/TU0k2F38gM/7mlRhBR4BhLnMnARV/RV1jzVm9YDPX
zeEhBnp7zbsRQeVgdf+DLP7N6mC3p8Nk9eh2wDmEmB9bjDQ+BhEq9XsgPE3zf94y6a9SD3ToxRfF
UszTR3z8nJCpBjbFkzh0tnLxA5W+YfJrRgwFDOAEGOdNJzcJ7z/EUSGvOUxQ7tlMCc4+BcdWGLjj
U+QxQ7PKMXFsJ488338I9mk0aw4IFGTK01NN9j8mqddCd8qw9vEUZEVLPy1N93eji/DC0mCQiSvX
uZ4vBZ3PMdkImvzS6jwpFcg1l37JTb/dAdT3AhUm+I10uOniDIh8A+8QWyRUBmd5e9kYHVJNhbk5
oMwkZDC0hWyOyJU8VYxojzqscOAkM39ki41bogki0hbhxSRXULw7Ol9K068hxGnGgpQufKcKp6Yy
IvltORCCG8wNg+/n8+VTEsVEDSb85+i9v3+/cSQf71OFP/wNRS58DHC2Qtp8BpW5r5UqsKPRa4EV
q02GkkYdpV8WzigGeNq9x1M81dNJI70LFCqB1PVunQTvo2J59yDh1xsj/7iB2Acga/pGTgJF35nH
i3WZCkL0pgZEOmsDYxm5Y9h5AI9aYuqLvKdmx55jeZsX3b55YYe5R889DgmsOHqnjEY2CxzFmh6O
NWi/rgjtnzCEk+zVkJJ59dviz0BHhoW8fdZ3dSoswfNCH77gFwcPTGC5sZxpQRvMShEEmhRFEtdD
N1UlNO3rnnU/iNuRfdgjeaiyknjbDUjAILoZ9NN5pRgR/u9V8CTVvVL3ydZ6Rc9QQekA4wZy5F9V
1PfcOpSZIyi/6Ff4nkNuspcMvBKr4EjbMwUbnrs2swVqYfRrNGNQN243C42Q4LhHhLH7jLosGsOu
0LwKW1uaWO+v0yf0ePpkYJ5ilU1Xox1DsQV+5OUWk70ZjqWOaMpge6PUDOzEnyg8YzJEKjiH9FYS
pTT8gP/XMrljpjXk5WVUDxGVJo34Y0GFtzIGWoNLDlYtAuIOov3/Lo9kn0PyXTTfxjRpBy6WNZ+Z
R3mJEFcm7YnIK5FSKB7II6nnKBuyZkUZDgrw7G1laX+q6sWiZLAh+bIpk5KLmwtdIllyhk2SvyWX
QtYanxFEfnTO5Ni0+PSjEE0qMPyM4nm3zmV5Is4VbE6mu7W9AxKd4KX0LxDhlr35R+4Jm2V0BcID
9nrFek6rwurhqrL6F+zj+NTXQ5JtkLFUpsPyXlbPa1R3bfjkB58+FxXqxSBMSM5Ff3wqgWIVDcwn
eqhYIkC9vChZZasJ797Maj+GrV0dhf8NAXQ7cplTmXGVa9LP149vdTiCHnH0F/78u9Z63NnUi9qC
6YxU34Z9jULN4ZAdFoWVi8zFYOR0L3a+UVbhEzmasGe8bWwcnUPE7lypQqSFEcotKfO87+NQ9IE9
P74z04tK+6CinIWOW+SfAxU0j2+0Q44DjoVwGXkyyLP3Eqchko53Z2Vk8kRk/cZV4V4xBnnqEkFM
klmocuB993LsFIFZPVxQIy/U8r/rq/Ak3Dt5o9v01u+wKhTuHXCFITUjOoReMOwNEgDTM2ThMKKw
s300tn2CKrtA3ui9b8e41Kg+fHjbagCVOntVd0ye5J7kdOnysEzrQoLWYvSZ9NFjIpNfYGHuJoNc
UkTDsJXJX96XmwtyhMpCIRrPdusVkaw1Xig8oG7U2ygIzQ+bBVwnTnKmsaPjpk6qfOezfd98j+2r
6TxuVpK89BrmsEPX2/pLKFJp8a9zTFcU71Flt3sFYXqIVzVxWr0vywl7E5PRknTLD7wNqrjzOnCs
dXTWr9guISICesF0diETbrPAGxfjBmarJSUKJ/dnU6xTYGJHu/eS3sgGzb5vc/UdIIGzNa8qde12
izmhidOgcvWe2kBUw3KYYBsCOKOXcJJfqVcJpz8QRXx+7ylN8cQT9/RNA/z5v+QBPeJ5dvpzfy6P
mNNUZiEh1bipYNIYAFsUnw/tdS9GX5ETviR2sPl/9gO0E6wi2gWZm9xBFoe2sSCJGfX/yqvLYB1l
CnRqarvhNsGaHYBAE0qBiIzsm3/46nN3glhmqGsCZCthRsruhgZJiz2MHGCUgsQ8/RoETC4Wp+9U
4hTs/b6UucnE5yoYKFJwof2kr689wh8llUVkfWOzsrQEYMepPZqIVKQXa0qhb0ZmXnSm5Q55BUao
0iOJ74hJANxaXrZ3JsWzSNsb0wue7ljuxSD1oHnqCb3VY17Rj5rCAZRVatZU/1rtxMSWh4nhPnLq
2KUclRusThImONpHBPStTvDa4mZD9LBvLa4BekyHNHFA6oozPsaSo2ZPi5vqA4/jE4UjLAwduTgg
OAd9m6B+1eIqBPwlcqs0ccd4vn1QBaAR1ix5nmB5oo448cRZIl4kF9u+k8lPX0TQ84hOCpgIkrTO
TAhlTZE2+kbew4UH4+dE3P5u8iZkqzowoKFZfaaHaqyD47lD9xTH2WdDhGroi3GF0kBq33+03QU5
fVasidyli+ilhQfdDL1DoXEYotPnW7JgojKFmBls8ILzN6kq+SuM6fVlQ8ApwY8PhpmVjQGZJ8wN
fhNll1DT7J+NNr4w/AMgyTmwHyCTFGHfc3Xb2K+LMmPZvyqDnWfR43R7l5htg9bxC16+aNKclJuI
eWKBkQWA3LyqCgC4K07GLhoI/iB5cJthMRue9D2RqkvB+zFIwHPytEWrlnx3OAdMeI4lxkVyLu63
Ggl1+mbdyFi+AfSKrRjQAnBFQcWzETIl2CL0UDdlkThucey7JDLNtI4k4r7I0inGjzaQAn7qVeyD
k9ujP0EcElFgoMOPj6k3w8HZupoBTTp8rFRz+41LGGeGGplRCcwlAvUvLz6M9pZurd4tIKAbNH1D
P5mq0+meM6OuwHPtAi9FPnvcFOhpiK8hpxa295l3COFSQyeoEaGMTbCCUA0nL1AzzXHfnpp8G6o5
mvs9itwZlGBTZpHKPpoel2YUvlR8FD5apEfe5Iipniki+eUektzQROUJFi0n0ORtPh+f/OY8d+zv
l7r/lnBrqisJlAAp5qFu8P2/osnpArdsH8tItrsATpVgAB1UeBCwRjpfRuMlHAxKr71tTDIzxhAL
gqjmp3lC1CoalEhHGq5pLl5X/DyvaH5JdOkuCnHcLik3Rq57SzLdzzUNkqb1bWOf02HQVP+WOwMh
ye2mA3DbOqTbOUX0jMOoxl9qR5HHQklgTTfYfvJ+trptciJ16E+jO3EwcY7JnNuC18oB9f2BdvaZ
+mwV7agybak8p/oO860IkZX1QeK9onoCfBKoHGg+kd1leDfs9pD0pP/7wrpDtKsoPCv3jzjJ4OhK
3FbSBAk5ZNWFFlG37r5lQqMlY7ULCYrju18Qu1uQHKex2gJMp0loMwoWMQtKvhy2aC2lEEdht7NN
6FfvrIKRsUNSGhoKNazd9eLP6Jhrsw73Paop+mKazeLs4XL8glg+J2Nf2g1IDrDVTn0rkvMfN8Op
rn919le+Weiaedh/efhIbxF0sSQHvzOf3GS6PQezuLO3/94IAoMN2WKHRUAJGCDoeE+BUdfrN7DB
EmZ6z/XRWkSYQR1Wnd6daU/e3ESx5XF2uTjxy53EolQYazV3/bFg2SFkxflkdHHucQawS82U+YZq
jclB3Nz1XYsItEjVY2QygLzNaA/R3k+mk+ESc7WudrigMFDUKf+62CnEjjRVpPIJ3lsco6dG/pCq
l+eBCEXRsUcvzeVLTrkYARuTs8XxZGrCH4Q2Y1qLeawcE6JJizIfqlq25Cw5xryz4volTRPHH9gW
hS7jlHcZWoQHgKZKf15ucZNNWRaCjQ3cdZ0UbxCMYVY/7mZFZq0F1mb/XbnvcPunRsTgJu6bJTaS
miR97s7+PlxNwyqiVrHTLdPZO238dSfDEdc9CGl/MLqo/CwvCmbMcCBKLcQFAjwqO+dq2G65z54L
iB1xACeDw3L93UgMin90XPs4afd9Xzopb/HjGVKL1tWsY8vWTDB1tkqWC+3sUOqT+TMYvmo/I1wq
duGOU7Mf/ysAEo5n4TimrsiWtdbz14IKmaW8EDgLpmFbH/QFOYpjpuWsvFQlOa5lKwuQw/vFiSK6
4/6Cl9DkEox38/PLH5v8g5MAjOVSwv1m8Qng5PnHXqMhCR512rcF7+epTrDMGurH9X068Uyv2FQi
g9O/IR8zqwjd9On0id7X7HCVQnNuAkcOuNgLe9OjJYUaOhMlnyd4bRZEfO3ZoDlzS52xrFBtNJhw
sqs7OSQaTTzVBtbsDIy4vmhyeXhaNLZ0jlbXqURmQekafeBdDjn+7iX/pJvJUtbKBL0gY3ETwxje
/yCEBHYpnZlw04r3dF8QIcbM5XPLVAg8BeXmkUaUN+7W6OgouTnCx7VajXAK6yY9EUwmjcSf1HXu
ScxhEQ/K+F8SCb/GkscmElii3lKUrfxKND5JOHn5QrdaY7W0aHsnIy7i12YJmNzfZliqtZ/oIux4
GUIwW737LPlxpDuz0pg/mdHW89WWESe4OvdOZ+94sgoJ3/P5wISyuRtV4bJnZJdN1ZWjgv1UZD1B
p8PEXcPr8nNps8GWkKXQ5dUDo06dI6zAVGgF0z0/u7oE7uECEoSao0xp6INagWOlcxnCHwGZ+yjp
OzST6Rq+L1J4mU9uwB90MkEHeOYE09dsds11PTVf1hrTOd6dJMDsTv7FjXXtVbIcN5HmEscJGaNz
1Ws4GjAO31gl1yYrhGHCArPpql4HoV8JD471THUkYMylO9vQ2He4fOv7iUYf5HqP3FlgU8nG+rQp
xKZWxkLTw+nY3JOXN+dbJJ55CT0u1vZQebYiFUaKLhZXdCcy5RwI4G3jyS5zbZEXXY4xpd0Y7IsO
qAJZJm689JgYGcGShyzIfXcADSAIPFMrxbVItUWGfXJQv+AHIVrgBcgieoWS1Von7dKPFsD6tIWE
quF3NcQa19P3TrjLIX2vFn4kf/EzfdMEIFTQ4A/6l4Kkoh2wuiVuEhcycGAnXpDheA2qsX1pWFtF
0BuKtcYsUWXoZ9pWwX/RYZjDz81O5t6VdJ3KTXvhVTTgcsQhdGiMgHB7RcS6Gi8/n8VXcddxVfQg
UK7bv6oU/w1GzA9i0UHqc41d6UBeemJC6XQ/fZgGKdfdFGbNqXwMx+oTRm7ciY13TfBhN1epi5wu
lHafC3pRXjc2BTpz8maFjgeON0AgAPJ//2ec+SvA+mGqfoO7b2xxHKpgdWry52ehdklq0herw46E
/3d+uldpQH+4dzowwkG02vGqpoB2J1b6XXzJ36DOBbfIBviofBLWgnb6pARc523G9KJ0dRM+t9Oj
DfywBwbfLLgKgCQmQNHlviIl4rHJChxNNXTkwGjrr0tf+KiI/5zRNQPCDsQTx+HgiR1046zazq5D
ZR92qIVG/Wxh/vxc6DM87INYlJ/JbU2DzQewVBBApUOQZxuQjRJmbZWw2/UCCGyVjc+9suYR6IWO
rad+KRjSmRi5/H/fdFylNEYCZR+uU/T+SGIqtFKKhf3CMjcGgQnUs46+p7b+f7wIfFpEOEE2F+wV
+Q79GWYTMLwZui2MEyRmtbRNHoxTSJ5oGVEJYEJIYENcxal3EKM7R61g4svV1f3hdGgStl+79gKy
JUBf6uvorDEK7SCKejJSC0gqbshF/aY15fFG4tJyz8C6uzOPMVaErX0uapHSqDVvtxp/2iEPSQjQ
IVg7dAkFxDgtPDDeUj9qQAUTfdg74CaGwPuEoidc7OhhyfFKn2pwC8yOFGvAXOxtuvyUOTytyEZ4
AMlwQX/jEUPyP3AoKZJ8bgWCk5ZaAXsA8dIF0pd9EKg5VBbZDFJoMMmYuVwxAxcZDpkNiRU/j8XS
YRmKMtw1FI2D68zgxQkcLYXBZ+G8bRD6kXGiwrGHrYmwEXGusywKxZ0+LznkDN6epRNgWBu2EKHk
r9uzoShWZjZnRtnTuRhznVQd+9zsSZB+0jjSDKNb2zhI5bEyiVxKbjy9hkMSnAZwUiAoGHzKhRCx
26DWrJG+PE6U4RUqsKGuoh0hsCUlsnfs3zEicPW0UMNdr1w1B+zv+2/T5dc9pp6d+zt8RlABYIOu
GLQKXqx95lgyCG2RVJyIgoXSpHlEmZ/ZwLFjS/AwpIctSoocD5wEx3sMZ1IZR/okseTGqB6frv3G
6nh4HNQnddsxd3cLKGPrdkGdMgcnsxkoSrECwkF/2wezTAfe3Tk6MXdYI1EoxQWpNM3tYYYFVKPG
dzrMbhtg5S4zF9xxlK6VKWo/3uL0exA8I+Cre8h+5HS++U1wdkiJaZr5FF3RjD9IemYub3azX9Sx
uUMMLVM+axQjxv4ItO+4ZTWilPdjVFrrPjwl4YIfxghFv8J/aZKTUsrRpotasxjeLqkLzhauAG68
brs3kTHMogjetRtO563Ku1giYxgXcskTy8hax1WPhqlKP5moHjEfXlByjXPngmPGbGw07a38FhXw
ZOh8AMFZGBOTVHaMmWQJPZ7vFOQzkamSIuD1Q0zUmR67kXnSHGe40Q1BE1/qTtvJ633AqmDcs7D0
9w6ZF0Oo85Wo9Ro7FVZQvFSiGAU/vNfv9YwKnuGf8NxyakZypq4Z1GqYtsQW3Jeo6WPsSSUVFc3L
EclTkor8jcuuuDs5EGOeERIiun30Ki5VzorngAEgTUQZT5NlzVRPzzBjI6PKGlKcIVFBBTTWnw+G
po89BpvxJO3C3k3uiJ8qhG3Y/v3qJtA/xeXGH4Y0fwlD4jXeJDW/6zbtP/zP8D/3j0cdGsl+nORL
Bmok945HJtVWisPoyDqQAtWNp7pNobizzQ5yHCXHdSJQS8M40y+xfqKEjnv26S4a6RJXfPttX4ya
j2aBuhoFb2F91p7Nw981BHjrSPQN7hD86UEtxmpmQjFiO3+qIYca1r/Emd6kzT1IFBnP5Ee16qK0
WVWjJO1rjuhGq08nMgHj9c07xgxOM4fMuS1CkqcZQ+D2Y1uLH29PybF5bQV/RXJq8ApgaoJ1tult
fahmqX5nhyWOxOCkQdlcSQDZbOuT4iKN7UWrM9QLwYxT3D9WZyG9y7kHJ2JKHYeypEC6+Vp3eO0W
BmSZYK1QBmVauBc2kjEPOjT/rZ5BiA6cEjpI6Q3PhSV9UCbLFC14fJScVwk0moG9SNf6df9smWY6
2FVtbEHHmGmEDAaY8UBhs2DhB2rRA6KV1n5arsAzf9LWcDvBuk0k8KcOSs5gSaADQnTeW18/ji1H
R6EyxTVUbhy38TBJo60HTUQh76AF4dDEK1GdrIt9K3hMsz1GptZp6uTUE9Z++u5wjqInI+j4mc3C
tX2h88v6QhxgDYBTzAn0dE/DT1/nKvHd9G6gGf48HepSy2yiYQH6C8xP3ykDVIgA/PdIS4ZkS9FZ
U/7kjUOULimWeRM14YRTExy72NDZefWPTSEcy0mLSawH7RETLdo0O1UrMqpDpXczdVdGEUtKM4Nl
Nqx/LUSwIUU54OC59MSiFL5kgRQTu11Y4aTRT378ZPukIs1N1HyPR46IyV1ugLC29rfD5TFNo9ay
AsH8izJeRfkyx+yXkCGSmswoA4Y+7VqeasjJ3YXuOZPNBU3TK0DF0IV9k+kx9023KgDruabYrqlt
KL/RTE80n2WhuHgw1g9SjkgtX2CU85gajWXwuF5GJH2jxL+NSJB/EVImlgsjWVozXLFbD5JIn9zE
C7yGX3wNQA1KeVM1QRoGwZH2b9GsyCLXCcKfmymLyx7OTpfbpYGQmSQPE5tT1ZI0qp9ZihMSfkUs
rAxN8wKrutAge/w62drS1UA1ARu7B7SNd3xTROGJ4nmHtTyRhLOmYHnF087OGJYgc8AAAM11tOPw
URsCX3BRjPMndZNjL9/P6E6tZWkS+C9UMPOOtNNPF96Xw2AZCFB+BMzVNigHIPPGNZXD4V9KtLQ2
mpQ65AOAlGwhy8k9ZgKoGdZkRKnV0ai0y1+6GbYKs4Zmm//UjmgOv0SsWx9lj3mJhyb0bi8ew4Yg
qOwm2ZdoTzrv/C3VmC5rQNCW/ERwbUXPCShQdwPILx6c26ohm61R5sUgESmnEt5PMtNBLoXuN4W2
eTH0CqU18JN3kaMs2n1ROIrQNTYOEQWqH59391wQtYEsYZObhV+OYUeMr+lR1Sd8ykv8rbxMIvyT
bPpx4639pW9to7WU/FLBGIkPMhW1eT5Kf9mnj4GWHmq1BM+SQpEyVyjXJb29klvKZA8SnBpuTfS1
VnxjEAFPs5QxlKKg898GAo5T6PQwRTj883y4A7l9nZS2taPrwvGOKCP2wpgqDptVLeVVXxom1k9q
9A17lqEEcngY4+7U+7NfwUmVHE7/8ipowUGug8gG9nO2hpdb+lqnAuevMLZ82LJP/WhXt4EXidQU
A/GpESYBfV6jGDtbzDjgU7LiFrNLcUt0ye+CeXmnjkRwL2ZDzGZF7C3FBLrZUM9xaM9FzHWfz5WJ
t7UVpVBs1L4EWZ1PJPlR01mzenKCHzydjJzPZyMCp82ng0Lghz5FzyHddJgIb1r6o56raU7v4G7A
/VfTT1+KiKFT4g8MFquaYtAPfGycclxD+15DLwye5MqIIngHpenrfhuUlj/PWpDdd8miVWk8Ehxg
qsL6RKnQp0AxEig4HLclNxRWi/2TwWIENvvozdNONKBAQYQKIIOMmv/abQwdpm3E3wKa7j7wDssq
8pCdiA8d9yxR0BoOJ7STlcasYzCWZEJuh408m9EJZhy0ujxBL1Kgeq7WE3vzjPM2YamtGvpNrD6s
JK50NOK5MGyJAxoTotzIUxudb3GJuCYjK3or9bVzMzaCnjeSUJMtL3BilnFrHf9SqxXY35l5W5dZ
v3X4fgyFKbxcwaipY4xCxZrh5Jpf0P6/zoLM80trOmpLhirAGkesBYcg0kp8AC7XkWHoUv+4u72f
QSE6FYcb4Hhugkx7S5cnUkOH6+t12eRbhIbEBBahgItX7OQsEznkWtXWVcU+3jSypeUkawIDjaQS
Tnuk2c6snAiykopeOblXLYA3HIGCuOQWSnFn2PuQAPvkWNek3G7y8vlPGC2saUv82pTwHsbtayvu
28dM/w0he2Lyk84onLQ3DYmmTbTxdDLURL4x2CvKTqaveR5fuE5FwDjI7goMfoEmmjd3hsYzYJK8
gAYPza/zmdqYLaisz40Rbby5HE/TNARnzFfA0+Z1XQzgjMpVSqbVBkONmit7YNm0vXt+l3kzWfu7
fNlcgXqlxKxnniC2HEW4MLkAOoOW+fRzuSpXchzZEJyVwjQXJLpFqUj0YX3LTdBaaKTh8H7wIjT4
olMeTwAJSIInOlNH94EF2uVM1ABs52bcJch94VJ94afCvnbD6tAtKHR8B46LR95o4ll56Hftzjr9
Q7+ojO6xCZBWRoI2bQMzgzW1lrvAT9JIwNsCiSBNlIlaVv09/X40SCHEzlEqPEoMt+MjP1U39yDW
fkY7xBv7WY6NTtR72mTsBoAX8j8UyKjOwURrggL1ujVigu3Tq6FJAtSq+fFwLv3svhXAwbNBLCRd
y97H/x+j1rw5xhrhAUDv7El5TlvaCju8J5eeuo0cfjE8b4m+UeU6XhToqBbx4iD0ftqS7kZVGNGZ
O1mTm6qrsY6hnE8sIMR5nEUvzKfpaZ3BSfAhtXTJjykM5/8Cj9uAgNBYV+2/z0AIdf2tWSODQkbL
hhrbn7EY9v5R37eUQFvKUDZ1lx7fCVogMHC7VODwwiY5bnGIoAhevrfzqtAt8KJanzDWCZB8vVow
IS/Mw7bQHdJMNxwifp0zPCt5lymBo3H4u+u4daieUBga5nWKLo+KnaQIlBiomPzxWBkuhtneg4WW
NQtIzwF9a46ln8Z8Og2ggDA284Y7HcjhjPHozdwsHswUjwtEB5bzpeiCNqD16bz0qPcgFFuNBP30
WoKG7iXsRwXtWAeSlcy8iiwYemszCwMnKhX7afW7fRc18doF0kHJZ9WZD0bEyHg24oY5WvZreJpH
YnbaEcYWOiDS4XqE5rlg0lM3o9WX3UJD9UxAPhtQiBL+7P7CiyM4+5RpdAP6VrHI9bEqp6wRP1hu
20dYfgBh2mi5xI7JMt7E4PzLrC9V3A+gGBPflqrtitB4QzrA0sn1z+TxxKeloAyNoZUiPDsV8jjd
R3GCrFkskrmUU2SkuXcQK7iwC5V2XJSFcPb7b421KVMDCsqbh+TvzrRyK7N12kp2by5JoUUS76Xh
0mNHKRO+BJ0g/trkGwsTjPAzZNK2RUWAhscZSYqjFp8dCqRuRpN5x2MYadFqXMhEHscQNTQKQEit
R3g/C3hmPk5ffC08eFFEa2YhuFease6c52GtBzKWgnlhhDZfh8HmiVAMG/cUKPcTgacPqJWYXXbA
Motlwy22IFBd1YZPwG7/jVCzEM6dm8GQPusZk66CQYCBozrNDlT95+4q14y2bhKi2y3zWN2o75Vw
tPcvZ6yep+v8KPLAD3GSfjKZUea1oNWATgyYZq8PwOHa3ehA9rMzY6z+JRyp/gYjC18db604fGLn
7Fmc1IYqT2MuSNmrVwgKg+zK8g34zfCwzKGczBN2ShCutbYxUP+XtM2uKY+0o9TIBiXk1RoqqLrr
9RUQNNoNuckdeZFTKrE90bWy8eYgvqjub4uyDQtGBkeSrNpfUf5dHDpDvf46aq9wIMJyTWKeGlHs
/fkyBtZTwoF5HSwXsiWLhkYqWpGJTS0P+XEPVJw/yUQFxNbYVBUbTj55oK3iCaBn6LfVE9lJNe53
1vB3fOWZcuNMGuxLTr9UGwyNqBPm9ebpeYtQjFIPmF9aCR5PNH8aD07tXEJ7QrR1Jy1ZGDL9CAyK
Qsk9YimdfIeBzXt8NlFdwsnD/fgDRGsBj32vN2rb0NUavslfc2nQyNtse0VL9BoWBQwftYSfdJHb
WNOpFFXfNJfkXlvliOMDOigMbP+UbdxOlREHg/w4kjU+Qo5P9CVrg54lB6dX9E0Slum3lJrYk9vS
16Y2WXd8uG1AtOWuD1c+oLq0LuJjACj2G0J5PN2fUs6EdPCOtYiDOMZ9bfrGVAyJoI4h8hwN5Yb8
T/wo6M/wZc0Bh3chSJtQllBGVgGFIP+T2DqIDQD6Bxg19EovXGi7/KP9orBCjzmdqERRtpwIkVU0
Z4rc8Qjio+mvqKkiRPRR+JHh7IE5uc8VaHgxfQJuNqvcdzzuzMFIN5oBOzYOrGpPXVY0CKSvpWIs
4uut+dLewTNVzd97OvQjiGSpNqRG1LtqjeSKxc0GA8yFzKvpvM+/N1qsSbIpmHEKL2w3+6aEQtgt
P7FDDpcXhWut9M+lCAYtlibbgvcAae62Et3ZgjicGN5sU/vHN/S+ABD6YxVEb2stfP4yAG30XUEj
AfIPbEzhgF6x1T2FMDSv+aeAbpK0vfkH7pARgZyVwVEU8aPOgSN0o3BWZzHiRoSgTvWW4VVyz6iu
ljlyV9+ML+4HqSZCUh86S0bcjmeQ6BjGuLY90ClOEnuCzgqNKTYWr5zZ4LkRdzIAW0G0FEN8HBJR
aee7VR0LKUYdD1nLtjgac5O6g5i2KCOY41f9xutMFs0ZFlow8d95cA+jcjzePx2/+mh4seaxH4Pr
Gp7OMePrWeItmYrCnKbk35RRSilKUb7Y+iSzGf+ANzUhB7I1lBib0k65GrjSrFqQtzITi+Ffz50f
TXB7Bvv7bPMPrgOH27byFK08oGdtRwjgkVMl46bYNjEzmWMi24fB9XWLHHGSMb6rwPE+nokYn2j8
DiIah83Dt3UYlQmu1EvkVWz4zCs1n0pKqo9P+RNa2iichIJL+5IDthkU7NQ9SGsDr5VuOZutx1LG
`pragma protect end_protected
