`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PjjfnTeIYMNtHIC+P8/tn+OhdLcEDzyt9Fw6O4nTGiTgR2VaP6A1+7qFHXyiXo4Z
f1Iefa/CfWgpUjp/j+hLJT5DteyOu8/VcBReEKOUlHAo15LZlG7XHPLOYbt+xRwA
MRddZLcaU9pk/xzC7QIQI/IT7GjT0z8zedMVgzNEdy4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3920)
rW8Y7X5ow56XlRD7fp439OdLgaKyWWlC4wzR1Jwceh2QUJ4X4QykonGylKYp5UR2
K7iQCY+KKaZwqy6DZmbZ9L1G/2Uk2uXgUJWQjD/XYQ0x4mXfSenb6NkzyduOXjzh
h3tSjNKuVBg7hIdDSAMHZkZYoewaAfOs34VIbYHfawA2N1ZaQDXpwRGLOU/8aZga
FXdiZMEvgpJ4iJa1OOabhC+oQYNg4amLimGBLX9ertgqK/7Rxplta2FVluCugUhB
EerlGSDHpsXI3tPOBmnL5M65w1qg3HvQSKzws5hl8uGuPX/TqeVFgzUA/ea56dcz
5CAwF1XlaylNcIGxzuQvkiUq1n95GSejUrIW/F9FZihPCsT9MtoLkE2nBRn0TEFU
w5st/0iaillPaDDuqejWUcRyxEH21Vgo1nXXqwwgcGyB4cP8laQtugttTzxjNQ6q
QvSoPe8ntmMu9vo3jABGwch0/Fdj1nKSLijWaHkcf4sKtyclix+NwLKVTGEdZWS+
antySgo1PrhrypRYSdDwxRBGblSGM97MEFbRloj2hgcMT6QQTbynitWwgkVjRlMe
ErLPlczGsZYWds8LHnIoB6YyHvssqqJjmcMp4znzE9vBNPc0BVttUsp0YB5veBDj
Pu9pUp+5cFuoa+vCSVJTrrNbhPQKXaOzO1E/ELprQJvUKQ7v2motFg+O1BuCckTU
wp1NzQXd5F78cfUk9NDtVRogBESC8cP8y7SC4KaWkffZ08K/qTReyNvnVQ2Adv9j
oW1nQMnkwvixUW9D0tsJSCmu4MWhSz1DT0uBd8pE/Q8rmflNxjjk61mfBs0+bjKJ
pWw35PLxUc3iKnug4i1SqgsGRJ0ytkCh3ofI+cHbzOoL+rE50LYZMoHzpRde9YsJ
jFihbUvPLRf48agkkalsJOp/yMvffnV+tBHyHyA1TZzo8l1hqcm1yitQnTaaSZgR
+TRKt5FN5GVu02y+jCaTCZpD2zY1sWKOlOFRCXja6X6y2njEdk6kJpp87fTxFW10
+cKozd2P/ON/VXrShVPgdafJWrFxhF0kRuOL8lxxDHJ0elD7jcb6OykVH50Bzu4y
yJmzkmNyihXU9mxwENhp6eEdiO13SZn3gU+payNzTfnZj5RzCQ/1s5UFKm/1UYQE
201Y/nOmd7tVRz7YrMSVBXMiEAItq9VHcwuGBfqKPRADAHTdofS8rHWtwf3F1kwA
dj0J6wx+KUK5ZvKU/DNpBwodWg4bQoB/crE3ys1G3P04sXDeEEAxzvjOTq/AMyHj
bQ7vD3dDgBd7yoMRkxbdtnSDXMaDBuMglF5Gi7W4ICx0aN9R5/wpl0TBgLWIP+Kl
LXCPGTtBbw+/3zpN8/ZEgdG82LJctPUDQ0GIIgTmYXCz2v4PA/8X/S9FCHNiA7Bf
RVcK07yy7bIlHNTYPH4Kdn85dEx9AZE+xpyPBuaE1yKMxLZhkIKN6Y90N7l7TRkm
dBOJ3aGLZMAZuCB1XqgX5TRi2i9lot5aoRQ6em9V3s6qgkqdFfToBOl4KsVou2dd
Tqx3bHs2gzymu3O+bCLhTCaSgXhL2TD+YvKHc7Qz44hfABJDAJraUuxOSLhTEeIY
TH78o7v9nFR/hQnsaCvAw6TZRDRhJ3MCk/AS8LFGzPMCQDtFTXaJUqRXZW3iAhX+
h7k8/0gn4kEc7HbNKAjTcQ0+/l4aBUqvE83/YaWff3LYJ4I19frH3G07tTHpAo4T
Fi0Hr12EIRzS66Opa2HtQMrBNFfNLIADPnEVbmajWISRQwPSK9jHC+JC1doeLCx2
O/zv0qbRHtvYTjQapQ8LHAzFm2Uuiok4kKt2Agm1UZiBLiJoVrPaBn//GSiYvg0X
SKHlTq+L6YQ+fKBvamXcIgc08u4NMooWZ5ytPDM+zrutw48tPQl7iHq1tOSy2AUX
ZSr1XHQiCkeJmF5ZQXHsXGwOFRrs92Q8quc0ZdUIeWCPS/aGT4xfvsiwT/qq1phU
hubJaxwLSOETtcnswtsvII7vJSvwCLE+35y/RYTwAV5vXWzKlUI8F4CMg17igMct
it7CL5SNrab8eM7P+QWdxGNZ30/fBFYr0X2x0bWs8L8vp+4IYZS0C4GS9hogiA0x
5p3s0610DgWpc+qBSE3DRhOUydMJUFLJCKxTFize7ax8aBCdtMhGii2qpLPuYg5P
ZWklZZDm3kyxevSMN/wz3pXl0cHT9etOQEBo8cnCJ6mmOGA+TsqJhd2zYrvSHdGC
ol3lESS2R7BOwJOXLbsqhq542D+rUgqSYUADdIVP+Vk5joB6NZnUeoFYwfoddXD+
jI0kY+/3jKmKZGRNbjl7rtLVhUgTfEWauS/KP7UYsxLnPKbTeewK4iS0SSffePXY
op10h4xMwbF3PLTl5xxWoCfyOWQiWZhPrzW5zl2blHrYZyZMLm19PDns5Wiwqc90
4yM5dxsiV6fIRXMvZkXAmTyCrWKoYaSM9aDj9/qFy1l73FN9ZjLLYq1bQOL+pU8n
dLAxXVemZmn1+74I6rtvptkR1HvaGqKm0g2HDjPKht7XjghbaGb58/4B3n532TZV
L9uJCQI7XYmF7n8WROy10rtTR3WmEBjtUW7VfGN4ktRy+Lwxj8NuGEpvNiQ2ULjj
TjWm5ThNqAudWJVxOD1imPTl19dy+gnNs2t5CVt1xOF7G9AK+8itSp3LQX3f4PiW
6xJx/vnKuFYadJoVAR6BrIgBy1qfl+XWzgtxjCznoJli3KH94f94wea010bcVZuR
sH1APBwoJ/1cFYcCdPuZCYGxTIL/goib1CRxebfa+zM+9PJSjmRjY0RkuCQIoE+5
+yK3P3eTcPVsyC6Rk6WD/dQA3BUErxuWJvsdIfLA4UdWNcWH8K2K5J1SSoJO6zGf
GwnKXXb357fz/UUHnm1813fq3+0bdXAijltKlV7avIntvJQ8yz++RgcwdWNGJv1s
8BJeaZ5hSS6Dm/MSkSWI6AFhuyM11ePcaN3XlZET+sBEDz0iqwPvzMrjpB9G4Fp0
x9V1bOjMzjX7NdBzIU3d9+SOD6nYycqskan1LEZixQZpWTwehj0Ekd9gDajj0k/J
cqhddDVxxkWDnjicj6LXvE0qt+h337yamRtnw/SsjOXhsa6lB1ICOQw7HiO7Olvz
7e6+6IaNBMsRdRXfYRWIYGASkicAxbWnNC8fLrmVV25pCwyQobYZwa9n0ST1nl2d
v4ucMW6p8TFAcaoSoiPtWi2ur2u0PrwBGPdpynwhm+71dvZMlhPd546bDf0hUWir
pDQ5nW4Xei1Mis/alp0j3G97/kUdQxCTs++iMe3mAzUiX8ImZEv2gKpbqXDiO4ki
GOfrHCJ9+MJswR0o+ffcjsPRIUcFx6GzTEvlfCnVMNff/4sNCUspgp3bCZytzTG6
s9y+AKLVLr30ibhHt7cvZv4eulPxCmGGKTM0kzNFMQF+lumAvIg99Cp27+cJfppM
y5O9LsXNKp8dyCvH+I4T3nRyB63aepZ37fSRoUsEvCFdC808vpS5bC/LUQPJiaBj
S7WOnW4ZPVG1+5bko6JVN974fVfnO6dsGAG0bsUdSst+EB2p9Og2f17CYEw0hcjB
W996po08Ixo2qAUqDT//Q9ip8xkfAoFfZld67Iq/hAz0fuyR1NyjdZGcNaT+69sc
Wyq9tv1Ulq3NToIAYLBnxx5shTh/mPH2oVbj0Ocwd4h1Whw/6Kc/Icnsdr1vmQ8K
SOk+k25PbE6qsXjd63Y6Cg0/dUSjVCbXdlHg3J5cfFnu/QFHMiNHISnToGR96x2p
F/mPKz6gJpcGX40TsgdCnoH9lxEt69ZupUDVFvJiDSwQmCdkD+5W+dn2ZLGhlJUL
oSwUq+A6qUZkwLknq6q9FMLnROGJDlHeYasXkzx2wDETGt/eQ0FArsEK44RQxXiJ
Xhefa/KaO5Wsc7JOrqq3Nlz14HlCRDTG1v4RLMnokPNaUEEzXY94hlvZ4eCA1b7j
ADyX7bp5bK4S+X2RLhI4OsqLze7bjYgH3areeDwcUfC7/eq3hVsDXqCBXoOvOrCY
o212yrCh/PD1i0IoxBO0C5s4pBsspuoz1NdTvzlw/Zqup4yRUoDALG3oh0QSZazz
2uT3xxVjbvykXCDWRb0yiz57+JLnx9QUCm63DfAO5L3hwzBMAv6FLNGsKIdh/KAg
dBCL0g1ZLjAqNk9+vLJu5RF8Cmsy24X3/pGZWsoWCyKruHZfTtiACIWJSGVHeVLD
9EtG26lx751/IRZUgPdFHQeJksYnyaDOCl1iyQO8K0PUoM8AY/R/QLZIPscuRq4T
iWMEy7JOvRrPkmmU/LD1wedfpcl5JfvAibhy56egNpzgLhjPZS9ccuZpzYvJRPNQ
nnWg3OdZEvP/5f+KKwt6Kjfe67u7XE3IA9K1J1Bmge0czDhL6BwmXPWabFBBd1lc
SCV8Ld0r4/NrrKHRTtgbSIhRRne2UdBMU18dXNgYgQ8ZH1prSltXrGpSCTuZHSQo
sWq547EGDvDkx8bPauOXu99V1ilq5tlPTDd9SyriTsyxKVEikDYtFR1rZYSo4u3H
sxDwrsBVKoFmYIUjwLTE/zr0LiLAclAgHqHg3v+Icy9BKBjGx7eJJ2Et+Uoh2lQs
755cHMwdqUJ4xNBA9Vdp+CsHUNRAVFUYvCcmqvGpbg4uCIXo4fbWJYjGaH12J9Sr
ZQj7Lz7MPl5TY/dOgNuxiLGHAkRyvhztOVA/XVJVNpfYzCjFUItkW8AZQD90FxhT
DLKFt6oKS2SSU5TB5KRhg15ZVuEhkajBiCGlD9ONvqg6J1tZUXtfeuzSy2S6ffrO
YWOAGrZCCjIKLN4dN/hb5nYORgikxJyFJ/dAMeXMtwceNkJKosTPfdiutCXJk9x+
KaB5Y/pEJgDKGuLvK0/HtcFUNU7gKwDZzBbsBqk3krzCsulwAq0FeUJ9LNkNBOAe
gk9pUC0QhuCGQmSDURnKUHala7QnBLEEbVB3EuwzD5zJEOS9Rr1NiMYsZzcT6QR2
pj4UmX3bGSCEipxki+xpZ87jS3XkV3KipXOx8IH/sMHT0BgU8yHjdb8MEHR/CLwa
B3Gk9coWouVgzNwqynPoKKXo4kGsAk6pxgEKyym5IqD7JuGAatyqROn4uK657/8H
pep5PBBHoBSaym/FDj2ZALMn0wwrtQdwWfb3DOdSJ1lo1neGrDG88T0+vgeMpFLS
3qCIhrmgx7ta0zu+ypJFks2oUrslRogSGEPpBChvo0g=
`pragma protect end_protected
