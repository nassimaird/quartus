��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG�V�����3͠l!I>v��c������{�^J�ڸ���V��P��o�&k�F��y.�ԳS�o�~�w��L�0�")���-u���h��a�e6�a'4V �X���%-`�Y�i���5�w�_�M X�����z�\#$�<:@]YL�67�6��7&�O��Ǝ��&�(�Lt;��LڌYI���*�Ē��2��%�IK�

����%5��`�dˬ�J�U}�E����`��K�����
���1�mnw���\��Ic��f�=������|�p��Z���x�&�i�
���p��0�\O*8Ǆ��T�^�nw��2������i��˶%k)�t=h�P�F�g h��0���p;����db���뜃�qK�eI��N3��`�|�ޯ������E�"��^�3�o��RTBgH�:GM\�6�Uy�1վä��֞�
w7��`ו�zs0������C�"�Kdq��/���{BND�o^�ץ3J�@��Ŧg������_Κ��i�[ܧիy� K���	�	����5�Fթ�H�����e���?&��6O[���bJ��~�K�l�;�J�L]Fa���ϏH��MĎʡDʑ�A%Ep�٦���qط�o]��>�~o���CZ},�̜PR��-�cA��A�'�i^��,��d۰9U!�o+��
��� 6G԰k1.ݩte��1�/K��1�祖��$d���PT��nh����=�
U=sK����&�Q�I;�b��9��f��yD~�p�����z�;�qK�ZM�7m��~?/gC����ˈ�މ��D�0z�Fg���Vl8�Ռ	~����������,��v����AC��{�,5ĸ��Xu�1��j�I��%�gڔB��q�Z�hG;��Σq��ݽS�����Ժ�'�nꝞ�����w%���P�����@e���P�ATGt0R�.���*�7f9�ۧ��b�����D�Y�*I�0^�-�)�f)�E�����#6Dz�W`	���r�(�=�f�o�ʠ�8�6DW?89�N0���,� �G�~D#�dl��A;�֜�ʞOp�I�talq'u�Z��l�|~Bg�$S���`����	f����8�/Ǝ�
�ݼ�6�
�L/��������Z�4�	߅�I$l,�6�*�j!�AQO���������<���1��_\y;����Th>�A���Ù� ki�*eN~���V��u�w��=�J�~4E����W���A��wՁ~r�@���6��g�;!k�����'�:���b0C��m1A	W�c����(�����z��orF(��>-I?����uP��_�C��R��?~�~�Y3-���0�魍 g�~�2l�ҔI������W(�妶����F���ˋ����(J{s�DaR���^����'��<�(��lHz�P�T��Uy�P!��ʛ���}�,LB�l�������ڻ׎���4Lhu4�-�a�;�Z�QӘÖ�@���%q����YiؕY�:��ri����;Z}�֛� f)8�g�ќ��:�Hj�e2�o�d�w�����_���	 ��f�=���_M���&��&�ߣ� ��m��
�
��7��t���Z�L2��.c1~�w����\�4�Hݷn9� �Tֽ�{��w����5�L(�7C��u�ּ������!����e�D��6��Q���O=_.P��I%
V���Ύ�D�Q�k�A��n������\D*n�3�[�2�O��ª�"�7�Z�^�h�җ���kZ�����u��tVc�K3����z� ���c��XN�%����XQ@u����9v�|0:�X�ya9H��-V)m���Ӕ��Ä|�mm}gy�`N��$�T���.x���`J�;�*��O��Y�$,��v}!����6�T=T&����}�&�4��5�6�3W`Z�{@����R["�$�����[HI�	��.�nj���}�xf��l[�e7z�Vfc����]K:
ޤq(L�³�1��y��ј��c��,�Q
'��x�n�ҷ�rNސ]	�S^JhOL4v�Sa+M���v��P� D�����¢�;����A��<w]�1���ƙ����9ކ$������L��kj
1���œ��b�Rf,7���7�3�n3&|�-î����>����{��GFKǒT����j�}ɜ-yM��pօ52�5�$���j,"�]:R� ��� P�=��}A�_�p�)]�8��H�t��z[b�~l�A�ՍM{�tP)f�??o�)\�мȓN��*bb�N+p�W���}� �U�F�
O���q���N�>>2H�<
<=�ޤF�#U�B��z� Ike�2ΰ���'|�0T(�I��ip�O��YE�5Vk1����:j(�j��s?���񬯤P��^�L�R��ɏ���i��=��l}X|��7��fч^���!I�p�pW�f-y$w�=l�y�8/�o���![�jl}�cS%tO�Z���>}�1`]�ǉ�Fq4�h)Ľ������F8ژ�?ýv���%n��H�IF�����5�y���O�H���WU�e-:�xKf�?�͡]���ޙ����IPC��n��wL��$'�4�~.���'������` V�����kC���fT��+�	ز��~�#�����T�8����u�z-���/HF�����Z0{��>g�t��6ܘ�s뾒�N]�݆����]��Nv�,�1�R�]��-��{2%�+��� ���3p���Ұ�_��;qU�ԝ�pΨk4S��O
͆�<�I�Aw6�3�<F0�ǃ�p�z]���&��w�w���0��	-eH+0AY1h���f��f�v�eb�� �<�#��w��.��-z��5��r�
��Rߎg�\���ڰ7@&-��taT�Jq�C,ϐ�.3�ѱ�\�h���-�|��t�A�g,	pD-�f/=و��>�ޅIb��i���9�h��ja�t�Z���-�FX����SԷ�T��&^�����oL�@j@O��AW��ɷ[��<��;�t�̱K�~�	�ǰ�s�Gy�OZ��+Ɂt(�c���5�m�x�1R|ս���2��@��D�~�:�}(���o_��Ŏ��e�U�_� Iċi����&Hߝ�c�$��4aa�A��W(ކ��,�A��KwF4箙D8=ෝ��MwZb�!�_��*���=��$*�$KX���yo¾
���d�9�8��^"���6�܆n<���X�+��M�\�Z�mEJ@"����p;eL�=�%S?:ڟ��~&���_\�v�Aۥ�|����.�G�`���I���1���Mh�}{~D�B\�<�b��)���P8�TkDvݪ�7�^T.��[[\�
!U�����M��� ��f�6��vy�~kPW����\���f��>���&P���Y�o�:�Ҹ���i�h�7+� ��`hǱ�z7_�B�R��pxK�oA�;taY{�vJ��3i�ƴ!U��@��E����X�T�������Ⱦ��p�:o�� ��wS�#6툇Q���0+Ǎ��1�TBT�����/��V�1����Y�@�a�����T�"Ɓa�Pj�SG�Gϒ����/9�Y��v �@9e`.�C.S�8oL$H�*,��1���k�a�49 Q��HR��bS�"<��/f)����H�9J�:��O�ů���P�R�KS�֏HE��̬x�C�|��|�����E0
�g���ɹ��Y�����T��eᥣS�xH����a��C�߼Nkw�e���`R�X]=��{�.�∫`R�Q��h����*C��yeVR)�\%m|3ѹԋpO5(���\�)]gt�
쭩[��fF;��!�{ �~�mk��M��h��cd9���8�u�Ȯ� |8��d����IE!�nr��^��_��|���9�e8`����u�<r����j�Y��F�g�M�٢��������~��_P@ 8
��`�:#���1��pٴo��/<��@H�IV1�VXt̘�PL��s��oƍ~*�A��Gs���ĉ���g}�F*\_��?�ZS
�h�|�,�ɘ�~i�5Y.�2��`����9�j��)���@C��N4F�:(���@�k�=C��_'3!1h9�[�)u�aK�g?��(=WeL��l�m�U����i$ ���)�|����
���疗��N��h1'����%g'-�
��"�-�ʃQTu�k#ٌ�@�h�69���!�ȧ�HgQҋ��T�Ԑ�Vw���/(M������zu���qa )`o�.uiç4J�r�r	���BAhTC�vU ΛZq�Z�[��(��)�*c�W:��k���dB �
�V�A7���Bܗ�� J|��=�=����R��yiwe'_��e�n7h��pO�C�3e]���v*e�8s�d���T0 ^� t�\����V΅�S�����r�$B�uSP*|B?V���sdl����#�vq���%$�rY��?�u�)-֜�t���p������:ZwAmX�x��ђ+K96ُڒm��ԋ�pw[AGX�#�IN�z�_t��K�D0b�V���U���	.kxK����Q���4=�<V�k�%2����}9�|�v3��� a+@���1
/W���沀[OȊ���vL3��S�O#'� ~L1�+X����]8�2�0��̠�P���
^|z#�J�W����]W?l�� �?��eԥ�/��TuL6��?��4r�7��7�ډB��_�1k@]��s� �	[tӓ�sU����Lu� ��R#q$�i63Z��]�u�0�Ս.�t��ޟ�_2�4GqpL�S�:�x� �zN�9kDb�������Z䟽�$Sz0C��?�2�k4��^^;}�d�Y�vn>�~�?�����O�;���vsz��6��Y<�N� ��=1~��yR�#ʭ�p�� ]�Sh(~��N*�e�	;�gs˞�>Y/˟�)��SLt�=�	#��J�C�r>;\������kG �z�c-���6�3\�f*u��,h�W:L�����U~Z�1�F=��4Y���gg��e���r�ӕ�(�����c;�[�^�X�wx;�{W�B����%�����/�i|���FϐǊy��]�����r�h5ms�����G�-޴b��շ�ҝQ|��ã&�F[����Ɓ��FN��>�8@b�gsP�&!�qٵ�.T�/�9�����5?�(nalL�O-�U�h��ec�fz�˝,?�:��@�!:�3[�d���}Z�z��9�)�IL��Qw3WZ��~ ��Ѣ�K�`M���|n�E��I���j|*{�Yٹc�y��X�í��؎�)' �S��΄�	�aO;��:ғ��Ml�yJN�ݜ��	��yB��㨡.`ũ@���#�����b�����?��4�����HK��ŝ�c
\��G/�Bh�R�̂��j�+`�N�&�~����-���{R�.iLr6��$�M��#���<����������X����"|�