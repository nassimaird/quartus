��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_I
y��������k%̜S���9('�X�@�'�X��m+��G������g��d�:]�<'� F��-!�k(�M�u�=X͝c���/���A�l�8��'?nZ�]�,�u�������k��ᚘYڏ㑠ڲ]��L���s��F�N��o3KK�+^_o;�_3B���'���f��jI��j��ŪD����8��3֓��p�O�P�hD�����ץtT��Wp��ZӰ]1�b��#�A�H��,�n�ʫ�I|�_T#{i;��5�$mX��b�"�(���<�B��p�J�O"R���Cr�7몈K����r��K��ΐ*W�`� �s���2q���k1wA#���k�b>����8��0~XӋ�ub����?�\;VQ��!�o�U��u_3��7��"�o r��-�ڙ �j��}��q�4(��jbu�h�b)h:������d!$_���E��FH� �%��?�V��o��[M#ߕ�>*8N�5DIba��lm[����������)w�3����#Gk��y��~�*�s3��£�9�eC��>��U���.S���u�_��D��1#�����\'��v���O!��M�,$�* dM��Me쎶��ʧ<��p�9:�`��[5�^�`�e#5{���% [��Dnî�]���3^&�'���l�z�t3�B�Y�ׅ����r��Rc���O;#��#B�j�R�&@3|N'h���Jޒ�1��j���%�
�on�{�����}��.|"�R��.�ڮ�6��J���ℳ�l�\�jS�f=��LI�gh�k� ����4kUϮoe_�8������e�'vSO��Oh$'�8�`�y]5�lL�����w�Hb�%�u�B�:��dL�>N`k�\������Ǘ���'K.Rr��
�yIe��   խ��tW���b+^�U��`���wK�WMn
�Nf�ص�w�o߹/|{�Ƈ�
Uf$)1tF}�P̳ ��E�4ֶ?��v���$�wy~]����zY����DQA�1�j��e��A�����9K��-�Ms���U^v��V�������Y���4��]z5�N�,���F��[T���L��4]����$�|&ڿf�Җ�`��*s֗ n�����x.� C�+HM@=��ޞYS!��P�HK�f>���=�S��a-�MY���0�?����=
Pv�Y�$Ov5$�m���#'��W4��$o-X�ڱ�
�ew	H��C9�^Vo��C����
)�JM'3�&�N�z���Pbo�=6��>�$0�o*IP�f�q���P!�Bn��p��ؾ�~���������'��:X~v�1� ��Zc_�˹�H�<��pk��vK�$A��ڍ��y4� ���P��PX����:�z'[̊f��?!`]Z�o�sh,���<����;Z����q��?`	���(���� �4E�:)P��I ���l��(f*ͮ6�����������)�9��វ.�g��;j��o��3�ʭ"�I����lž�3y���K��>��#\P-�(,�	�qo�*@kS�	�v E��Em`���Ґhk���G�iŸ	���x?h�(�K��B��FdO��]�2�����4s߽�*�ysO.K*G.��w����p���/�`�������"h���@�Z��p��sSn���B����W{�7^��k�Lnc���X4��My����J�U顺�r��q ��$��5�3 ��+�=s	G�wN��>�B�a����?[�X�3��[��6:up����,���̈ߧL�Ô�m��r0���qϩ��a���PzU8��n�ڲp�:RS%u�j2����	�+X�3]9�aE ����$�m%9}ڣ<�2��0�m<D�	*��b�DB!&���=hs���)7l{r+v���𵍡5������H�ES�k���2C����%oV9C���	dU��-��ܵ+��_ݕ�"6��ǅ{�eɂ���-�k�u�.A���Y��Hjپ��y���rr�*Y������1��Vpz�k�Ρ�~�E��sEA+�k��V���Ͷ����O�WjA �ﭛ�KԱ
1X�?$$��@��-I���vTF��i򶘒�qlFB���'sYN�a��A#��Y�V恣J�Bz,�C���-�2g\1�D���.V�JWq���:����:9S��y!x��d��S �����`���Y��>��
 ��F���K˘䱠#'oemw�#�M�����H*( ��?o��uD����|pjxP�ˡbjfʞ��5��o[ܲ��?o��(�u�-�M����Ri�H+�%�g)^��}o��L�^�ɐ��� E�W�`܂<M�s(�t����[u՗`j��i�e�
w!�I�rf~��{��kL�^Ϝ��Rh:��D�\�.��u�q��!R�Aw��3��&�\�%���s/�E��.¥{�[�����9W�P���=�@/�<���_�Ղ(�h�_���wb� �{��;q�~��C������r�A'1A�1�g�y�=�w���R���Ȥ��/��OL���|��w
�oiR]���M�ˬ��ҦG�+�'r�nKؖ��A|�0�뢈䫄ӂ� �Id�����Ѥ��D�T1e- �G��\�����E�d�7�0�J���J�8�6�e��Kg���" ![횾��Xǃ�3��s�a+�?��EC_��ιhn����1��I�1�12-W�j�NT�LL��*Ip��6x�}�c۲o�`]Qữ���!3j�yf�Ȕ*w�d	�C���`F�S��p�gE���7�\|m�e�Bj0c��Y1���?�~��B���ksyK��i����ݙDΪR)�F���Hwm�<��ϖ'�w��X�/m�~@�Kl��&" �ڇX@��2_�� M����DY �{E�����d~u���;�~1�S-�PB-�������t�����I(bD��x��ᾠ�N�p����'c�X��Txge����W�Y�u�����J[*F���͈��,Ju��h���KiwC��Ѹ?(��-o!��i����)�q�^x�@*��{?~g²�c��- sR��b?�r;n��޾X�N8�?<KD*�xO$���l�� BA1XM8�E���o�(�F��e�+�z�K�cE"<�rG�f?D�	GH���Ԯ�Pt��b���b�E�9��\�uX�	��tZG케�G	��6	�Zc�е���N����>�:�9�]�$�$۠��D[�i.�^��f{�D�w#c���Y�g�o�Ʉ@@����Ye�����$����0�J�6�$����H��(�ɝ\஡�E	�<�о�6Hr,�^���sB���t
�ŵ��4�M�����l<�����	륛�xac;���v^E����>�h�G�X�^|ġ`��I��7����QB-ix��dO�e3�X�\X��C�^�~�tq0m��9��3H3;][�I�n_����z�b��> �ޭ#R)l��S��$���w����+8#���n����B��p��kc��0_���h��z����
jz�_ȏ�E���eA%�g}W47[6�KR������o{L0nq3���h���[�<(��P=����іK��Bj+RT3&�,�:���K�a��E��9�[�j��Rh������;���k��x*iw9�wIT
�4��K�1�+[�s˗7J�2��S�&���'�-�!���^&��b?x����==�̸��)ƨ����ŀ�(��-(ZR΂w��>J����4�1��h�:k��K�������Hq����}��r�nᛄ���f����|` �[t�hP�X�Ut+O������h�^{i���=�[�M��>H)c���y^�B�m� H�>�a|R���|GЈ�TMv-Į��$��F/q޶�k��˵�-���&�	L:��N���4�Q���j Q�a�$���J�� �ږ��W;+��֜�4G��U�xu�i�����n�f�9�b���!�b�F*�{�/^���p˫C����6[+����\"r1�T���!�o�B�s����so�X��ߛ� �����ڠ���1�Mt�4B��un�y�TU@q(I�s��`8��=��9$ߖ�1�Ar��sP�&�K��C���Äٱ�ti4�T
����`��Ч���݆,��U��I�"�FA��^k���1�3�Sx�ɮ��/�X�,}h"����n	��:�1A�g��=�I%�z6�;�m��z$-=�o��_���U���m��7��$F:"�Y�n�('�\I �����#���O1|}>nXG��� ���[aHr�D[�0>l�<b{Yb�y h�!�����,RĨ��0V��0��,��Q�_$ӫ;W�xT|�s�*G定�D,84D��&>9���r��ƌ�bU��v#��V�'���v�����Ap������S(l9Ex��uXV�B]t�\
�؄:V3�}�<E�$���qF5|�~���W��>���!'���<׳�Z	�k�=<�ԼV�YE� 8�azo���ɌX���?��eit:]�s�?��_�ڋ·����ٓ?�%2#'�s�!��7޶�Sz!e]A�}o�
	��v�	x�3$0���pٶXڱ��˘e�l�	�rh�!�bb�`?!���%�]���A�/2��5Q��;��4�R7��/�_��\����e��4�$xA���K��y׉\�����?=���7��u�[$р�t�6Bbz�H�ټ�l��=��DS.�~�L:(�57�g������M炊�����M�1�K�A����`�s``�I��?9���\�=��M��z�z�k_��}��������m�f�c	^�ݭ�|���»�-q�)��?���I�0,��脶?jc�r�+xm	4������&�nN�{EYR�&��у.�v��YFN.�Q���[�"=yp CZ��M��M}P�W���%�I��B��TEWd"��I��)��T	>�Ό��n�k=���4�®g����Xx>�8����f>W�*�ҁQB6���O�@�-�Y�޸��������)�#;	�xGR})}u\���U QȸMMʰ���&Hֻ�+�"&/n��z�^��Tc����)an�J�S'b/� �����m��$tb󑣞5ۛ+=���<���X|�S";38�D}���{	le������{��� ]1|�!�S�}�o��ovq��`��h%�x���0�G��u.�L��	:I��E� ~GS���P��?p�7�$��.�eiR���5�{�Ѓn!A1B�M�M��D{T
��˼�~x]��Ũ<^�Y���}t���]㪔的�wj�|[�ō�G�~�}_�L_N��?F��t���
�M���ߖ�$�D�����c����?����5���0�y�4Bl$�vN�[�I�A�׈�ԘQl��**����2���\��L2lhJ^�CXa���4�� B���

_��ӻŜ�Bl�H���p��pॵ��J8��HRDN�Z5?�W=^ҟ �s�(]��b�#�x����4$�VG�2u�_��@ѝ(h0�0!�d����p��e�&ܪf��j݌�(&��:� y�G�$��Ӑ��00R\u9�)�f*�^�^���"e�� d�BEl��;��2E9���T����� �laaz���:�畣���ӌh��Ű^
˃,��7�<s�o�M��Ƽ_-�]�)���u���`�w�;�y�( @τ%�s_��d+��Ǧ�8"u�B��?��
���2I~$�\L��K��	^]>���9��&/�a��uʊ�+�n�ѝ�O��{,�_�?[c8�3�O,l���7�X"���li9!?���)�FT�
N�7R��o�����b�4���gO��>�
�����R�?�ܫAs����F'+��[Q��~�$�uq�����/:ju�s%�X|t]�Q}�w�llx]�)�(&3���Y�OY%Dި0�h2vd�����덼�?�*�L7��2�qA/�Jg���<�u3Uk���~K�T�x���M~����A<���8g�D a��5�Y	�aV�G�1�z�3d�$3���eN�쭲:�9~'}�˾��7?��]��4%�<#��m]?��KO�8֐�1�:���g�1	�U�FF۔�Z�ɲ��:�(M�:�Y���4�{�%�s�gd��@�}[�Yo����=��r� ����I?o�b�*�����L�j;��PE�Ϣ�KZ,��X�?l̸"�bF��+�Ut�,�7/"x�-Nxz_[} 1�6��Re����W�W;�\E�ݓYw�f���ܮ���݈N��N�vp��~�C��p�l�>�3�1���s�WPhp��"$_���T0ʭ�|�2x�KA^F�	�����w��'��'Ğb����U����<|y��5Ϳ�ʼ�8�<�Ey��) �dr[vo��CS_waU���U���C7���3욾e��?����z4��c�}(�6�b����.w����m.��K=P��3��]�ߋ����Py��>�x���Y�T�#mz���p8kiJ��1�l��
J�ۋ�0H���?�aD�GE}� 8�Т6ģ����0��`�L�Y�Ǹ�����x� �'YX�{�m��ӶO,��O��Fwز�����=�H�3.���E'^������/��SP-��I4>�1ʎҙ�}ќ�;�tܲ��o�Ae�n7"V.� ��z�HME���8;�Q��i�{ߙ�H�� 
��/���\&�cu/9�_%r-}�RG�Qӥ��#�nm�j�_*��>�2Ցd}k��8X�m_�Vb�K�vmn��b��H9�8����ͯ��xc�Q%+�4%�ǻ�J���L�RC>�_��T	\����͵M���<�쏤������ڿ�D��N��tj�*��bz�f��to��bӨ�qT�����+G$� �����.
�n�i8n1)�	N��u�,%�rt������ӫ.��M(�"����-x�>
���h��P�UEZg_ג�g[O�L��q�/��r\V�����50��E-�q���J�-N'�2�#����=4C�=�c��y���@/�)Gv��6�;��%�ڞ Y���%�|5���%7 �)�ؼ�;L,鑫jo�y5��Kz�ڞ�D��0^�CI\uu��˸�r�@&���G\��}ilԢq�=R��R!��^'�a�X�T_��g �d]`/�<5m{�j�Q��^�T��qR���K�b�6�A�}��3>;�3���\��P��}���Z����
��x�XJY�j!�q�m�� }���V'ĕg����Cj��
�)��͢��Ap�ܡDc��C T`Ҁ��R���hr�����ѷQ�.$�Cѵ$�+�v��>�Gw�p��Ȟ�{�L�ċ��E
߻�����`Y��B��j+��<τ:_�U�=�y�S?\<۟ v���<����ݐ�8�b:Rs��%!�>
Uf��N��}� X ���t1��x����7���뛬!�[�Ws���^��q�ă�+ &�4|O�\	2��a];�/?x*��h̲@��ْ����.�X��E~mA2��θ�����tQ�������zY�	I0�Baw��+�� ?�{�HM���YhԒ����~k��8��[,����LVz���y+{<$֣�/s�n>�6_�Y��
el��jU��g�=�u�yY�iE�����Љ�5v��௜�162?����U�Ŭ�s��:�T�Mo�+�&d\�NT��窏� *7)��:� �i^����*����G���а<͝� ;�X��8�<e͙Y�?@�-@^�W{��x�;e ��8ׂ�R�V+�zg+�vS��5���1�#�ٻ<b�`V�xn�� �A5����M¾Ҍ�Ǌ�d����#j���q�6��vtWq�em�vHD���6����`I�L���*x˲/��T�+4ٟF�T"�� �,��j�+0��Qhq�{�@�bF�oɭ�U�?{&�`d�>UVK�ű��+=�;��M�Y�.W^�/�����_?���4u�i0[�J�ʝL{�:1ǧ�{~����Q����"4r�Xc65_��r��<q�l�M���j��ӑD�!�e�*xԑ�gGŏ!�[틅�k�h=|�ܭVfLpRk��@�@�~���T~�*��h�UD���dEPI����Z�]V�@K�[U-ۅJ���\��/l��%���Y0��P�p���+.���L�Zd�PV�>�~�22�1Y\�`(��&�SD����r7hn҇`	�5��3 �G���K��=o_�Yi6)vP�o]9ݟ����&��m�
1~����F�Gۢ�g�8օ0p���q���Wxs�'~g�� W;�w?,'�ZE���2�e���>��<�%��L�G���5��CNY�*v��ȿ��-��,d��(�p��8��:t�y� "�#��� i��مļ?��k1�V����T~���!�X�Nh�%cΖ�B�Z�n˦ʘ��2�&��s�Ǯi͇�2؛�-����k���5��������ή -֒�Q��]a|Z�6Mb!wB���3�6KQ{�j�� �(�Pb(p�� M�x=��`+��E�?��J�4,G��rZ˖��'���N�|�E�r#;�D(M%9�y9�D����e$n����t�̊ ;�zO�-µ�cv�5��P�������O�6��;
,m�[��=0x&�̛�!2�s��{��~Mt�Po��W:X���b?�2���?>o�f� ��i����ZJ�C�V"�Oũ��
�2�GY���bU��ԗ��v�-)9Q����'��ѫ[��җ�&	�'K֧��}�Q������B̶s$J
k����ih��G&F��]y����7R����16����*����b/��,?��=��&![t�R\~)%h�>��_c�QHc0��Kf�&�2Y���q�1�V�{�3L����T�s��YX�E<Lm�3M��Eo�"Odٷ�ģ�t��)l�O�r��YY�*.�Հ�6s��E�3�8^c�>Y�VL�'�.F#\�R��l'����*�4ș\��!Y�Bn��h��+�M�qc�.c�S>i����q \������=Ҿz���s���'����5� �VJ��	�$�	�V٥����	�������8���[y����҂��;�>r=D�ǳ�1�3���?��3eיּ��<�`�"����i�%�iحXO]�8�$>䫸#F���RsD1c�Z�QfV����-<?��z.�E]HL���=TL�����V�w��B�ǒͤ)* 6�Vv��x�2��e=��=R��؉N9И��}�
[�O�~��4���U���ݹ���=r� z�|�O���]�j!s���i`l����@���(��'�@���q���a�vVp��{��S�~�(��0�I�i�;i�w�L)@���,c��><3��sU2��-=l��z���Q]��*�O=9<åoƁ�ƌ[�"'T_��=\D�1��xu�Bb��A'��O#�\�~��O��/t�ƃ(�
w�7�byX3 �Nh��(q�RA:G�I���_�t_�y`�q��v0O,!�A$LaxUh��A�o�	��`&�&�${K�<�C��m��V7VK�O�D���<~�F��f/�A|�@�L [�ؚ�噳#�ϘDso�,x��l��pPƆ��k��*���_��,�҇d-��FP��g�����#��V��as~M�T��xi�ʏ�"�w�dz(� Z�֞*�ө�_UZ�a����@X�@h�N���6�����B�y������u�8�a�B���C�X9bknb�^Je2'E���m[:���t�g��k-%���	�Ojز�m���!�TPO��S��%�2��l}���|��6g���~S��bS��pR���	}��^�~]V+P;��`*d~1fB±��O�r� �}&�U�7Lʀ��ӑS�U�xcuÎTz=�u�}�8-��f���@A�`��S��kӴh����=u��+-��Uo��y�
��=���Lf{Hdq��w4L%g�tU�C���^�P9hg�t�nb�ꦈ����m1R�y5T������v��"RҀ+�d��V�'gV@�����C�[Y��đʈ%��+U�-��B��>#�!�L���8yZؒ�ps.���G�Q��*<��%\���
@�h������F�$%���� �T�L|)�J.�W��!]�F'�Of��]"�7�븫R?����ɪ��;�3(����⧽���_{a( K�}���2�c�S�O�l�%JS"�O���w��a��<��DC���`���6A�O�%��C4U���_�'�u���񪔍g"�$����,��YJ�2�
��|_���Kˊ�ԗ���r��kv��~�v$�5�8��\����͏.�뻱��5a3SԂg����ECH22k(�˟���)	R�6"<��֌��n��E�IS��m�η����0l��"��~�~V����:�@(_��� mYl)wt���r�'Xl1�}��
��`����_=o�]iؙ3u�[X�橅b�$k����^+*��\�G��Q�j8>Sg
�1�j�{=�{���||�GCI�#�6����'�;�'���g���pnр;JV�ë/��hee��$5թ�_v��N�^�l��ع�]F����a��8`�K�LaEL��\5����-�g�@��j��/
���1�#m�2�21��s�S�ɭ�ؚO"����1K����z�=��jKm&Z�Q��&�-��Wy�aQ���M�jpn�C�����I'�B���H�H����%p�������ijTN��ɫ9���s{����e�uc+��K�s-uT�Z���#�۽)��0>͆h�6�l��=#���J�72S^Y�O�t����;���R@s��h�s��P�H�5x7i��CN�/$�}�
@if�s��C�+��V�OM7�j���A�3*����H�����O�o�z:!��Y�����A����N�/�f�ʿ���޽n
�F�7p����m�b�l7��i�#�;@33T��Δ�5_駕Z�ڝ4�2&��g&��F}�<�Bj@k>z���U�+��7�3�i-������V��H!�u�XJ�m�K�О�X�N�pҪ">=��Ѝذ �:1*���"�G��B��lu~f焸i�����г��E�2-��-:�㯰��%�&�bv�n���!��� ��s���.�y9�B�pT��>!��J|mD�bӁZ���k�R��c��E�`�HB3��� ��a�y�8�1~F!ďsnp^���o���׎��ތ�b��oiw�_�UE�;=k�m�r؁���ֻ���2e�{����C�����U_�xIb_w���̺��r��ϦtD�|fvxB��qG�0���I��������E���	{����0��g�����JX�`� �21뜖I�9u 3bPS��أC�7��A*��5x��q��(MS?5�	J8,)B���p�9�a�����Bn�n�K�u,bWF�s)����@re�841Ab�=�h��jِ��#0���[��w,e@jش7=]�Mipm^{��~���vè,6�*9� �4Jݬ�h������V�3T���.�}N�A�T��N����S��/���탤)ci�HIAK�ψ����L�A.���ň�:�c��L���:�� +�]z��&/�r���KA}S��{
Mo������v6��]P��m�J8/�2�YdWO������[�~�5��4s.�XDK�5�G1�)����;`�#��CIG#�5��m�3iM�m6�ȏ�&�9:���?}���R��p�$�RFY��^���@�N�����3���Z�+��sP���<O��E$��7�AG�T֡E��%�
�7k��즼��Ӧe&9�5- �8c �r�Ⱥ�P��X��ޅ�%�X[@f�Ai%c�^"��0����p���i�ϠȘc�Aѥ)&�g�����?��L6��"96| RH�^�E���
1v�=ٵ���$����(�}#؃�^[�tU��3*�8���9f�Q�#)�=w�9�R0�Z:��|k��%���V;\ �2؈wRV�GŶ�Qd�����5�Y^����F�cf{e`��Ơ)W�5�{�4D�zX�<�nkN�vNq)�b�+�k˓-����1�"��ņ���ΐ�f�^y��d1a���!�Fki��J)�0aG.+~������K�&�?$9}��z�8���x�>cȔB|�ܸ�3Do}{󏱋�	� ���C�
d�"�>�ǧ�=$�}2���:��SL׎�]�2��6e?���yus�edY^�	�\�I@J�7�l�*c�mE1Y����U�zſ:����&�7	WC����s�U��L�_N����P�OA�Y�N�7�KC�́���2�ĩq�+�l`nq�ԫrgP�G�� H���	��֧���L�OT�??��ى�l�0�1F<Ԋ#C�U)K޳5�B��>6�$�q��3`T[��b9E��T��b[�s�1��Z������GT���Nq���Oc1ݎp9Q���_�Ed^4b'r�5��)���Җ �K��+���� ���i���I}SM݇^��u��k��O'���G�X
�0�P~�����ru�j��P�t��+wQ�xQ��I�g	�X%N���~{�����Q.&�� �z�U�^b�	^��L;ͣ�LH�[�T}|��=���C��Q��NT���/�8�H�!�{o@|��8�@3c�����(����<�l0��2�]�����~��'��o�����0y��{ꬂJ�k���i���^��M+�`µ�j�:�]HvV�$�����m�c�;M�Iz ���Խ%py��a��A��#Ò�TF��mN��	n�o}b�G��-���n*�S��6̠C)�N����PV��K�$hh�����\'�VyĶPۓ2����-� �DE�q?%|���Q��l�Q�c2��T����<���'��[���nDgB�|�O��7�¸"������;��X��Y�3g��_�2���G�y,c5�}Em�Ѐi��k�#��� ���wA�eF9�<C.�$��l%��Kan�U�B�AC]Ȇ^�i��t�ޏ2�Y�i^��Z���U�� hQm�{� �E4oޏ�<�n7���h:�~�y�큢�McD�s6�uS�����fv��~�����K��r�Ŵ����fA�z�e���4_l�<�y��=<oC�Z���<P�tٯ1ǭ��a�"��qE*|r�'�g�qka�y�H�j��9�/
p.�� k���Ԕ�=��@}�6 �'�o�p���+ ������(v���B���.t�s��4m���$A�*tU�k�?������j���,���!�P����]�nf#�#���J�L|O.�eK����Y��cR�?�J����bx�4w^[�ed�=��e�	��4 	�-�Zd��U`(uc�C�@��L-u�zuVW�Zb�2X'�G7��Lx�,��z��c�N�R� ��%mh��C*:x���I�ZcґP؎?|՟f�O������x�oB���WV��p��Y�hT"�Tpi�f[K��e�J��DVQ�Q?������-Eg�^y���C��в��t�߫��5��n̯�K�پڛ�|�n˂
���ߧ��K�L�O͐������AgH`�ZTy���&xͫP
��aIlK4v]V':�|��Wr�-8=A8�|AX��8aY��u��!��-�BC���
�̢��3���X*pE�ū����|�(b��L�'��:'[��I��~�.�[4���la�IU���_v�cπ�*���U]�N:�o|/���]R^C;0�?2��Q;�P���Fn�v>]ȼ�� ь�J���=��es�t4L��b��^����
�EU
]y��^Q�$M����áx���	�ɯ��6�_��A�Z�����'�$�\wȒ�D�)l/E�f��HV�˯v����u�<���&̿���,E�GXr������oR�`��1�!`^ƿ�_���k���A�Ѹ�MP�|�:��9z�X����2���(^�T��`,U�3��4���G4���[q-஺	���
�k��s��/[koG��X��	�@��r~��<f�C��.�Y�~�#iС�lf�#7�jʈ;Ep{���wW'�jxm�A���O�I�2g��y����ci�bM�ׅ�y�`�PF��n�&�;�8r/���޼ZЊ����;��zOÕL��N��"�E�I��B��@��XѢεr:&��uD#��f1�òەZ�ۜ&��a�]�N�2��%7�����p���ʸ_�?o���r;�/WO%��ָƥ0Г�3i=J'�������jܫg��?z��������c5 ?���65.����D���8\�S,H |��-^�q�~�BĊD=��ˡH���K��L�p�2����d�f{��`ÿ��H��_O�#=��-{��,�m)�̤�}��J��&k��	�tV��q|7������l��E	���-�w<��Yx��Ddm�4%�e�LdV[�	fl�s�5E��3l���O<��M�A:{-r3B�'q����v�6h�\�t���i��v߰�=���"O�[���ˀGΩD�؏&��n�a�I��Үw0�F�b��9�1���$G����Q�Sz�߸�)z2���0x�q)�~��)��H3q|#���h\��G
�;�T����r8֐=���TK'��������Pl��;�h���K0h:�͢���z�XT�͞����vY��c��]��H_}�m�⮍l��XTz	X��Wh�����'�x�Y*�'��z�}��v��pdM���4?�2��	�iF��]I}�'�6���d��[�9�Y�z�|��@h}c�ي3% ���ŎSr�(~�Y�o���\����i��<�퇴Y]�X�e(��F8L���0}�3�R��aʮ��\�2V��n �uuY�υ�̊{�
F4���P^N�;��? j�x�퐀+5%�yvo6P0��ϩ�e��"�SU��]H�-r�#'#��?L�ï��0�l��9 `X��,f��XC�j)����� F�\�����z��`�HT~�S��8�Y��^._�J�p8���}���*��z����2�jo������ͤ򰀣H�ᬡl�x�R;őq���\?69���N�_J�� �Vr��=��ѳ�e��cv=v��ߎx_Q	6%���f��.b�Hz���j�\)�1��Go6Y��������[e�@EW���(��<���@�~�T������1�&��L��W��� H덟��Q��~��ߵF@����0�����J^��=��[7A��J�(A�qٱ������̡h��˶1���f��GI?��1���SEUQA�[��c��]+4	�{�1S�N�=fvŎh�e�oJRθu��}*Đ^�wE�0��������8�W1����X��֩���\cF{29�ɏ�˪�j�B�F���M�6rt�\�b�>&�Q^G!:*tƹCH��|�rj��F2���Pf?� ��r�� �O��Jj��Jf1f	5^��1H	ʃ"ZU>X�x��ft�<��x�ã������J��L~ �e��FPN�9O-<�i��^��D\m���Y���Z��L.V�I��H%k�t�5J���/��vw��5�� a�:5��T���j��<y�`��'S*�
����+�{�{��+��[��\�O���kh��n�,��`�3��0�2�W�L�:ݺW�C� ����H���^��Ǟ����ð�e�/pI�D�u6�!�^�[b��ܹ�Zl��f���|��g$�ᅸl����m�[������'�dlMH/�B�O�Q���mh��;�p.���1���Q嚃�G�?�|��ȱ���Ox���ؐ�Z?��/���]6�/̬Ϋ#��oȖ�����mE�IqN0��9�����KX0jXG��-z�eE�Ha��:Ҳ�����!fΘ��ܶL�x'J�ne�.5�ë�GxL`��[�;b�Vo��ms}./��.McZ`����2wQ����X'Y8Hhg6�΃�x���>}TKi��<���3��D*�Yo��~l�
�@��
l��D'-��A�(j<[�5��YJͤ�)�(�G�(�Ifϼ,e�B�j�3o��tJ"+�~��lf�"k��)���.,�h/�cu#.�>82��!�⍌�%�$O�X��D����e�p�`_L�+I�NZ�(U�I���֟��^:��H�
�m�t�'��~�c����|����7��g<h�%��VJp��Lp:V���� e���%��	&�G��2���W�C���^�
nQ�� '�0��j
�9K��NYa������4Ϭ��5n�q��Q��Y�:d��p��:U��2K|Vmj���E{$�y��v>Zu�a�`i&�!�}���_�\�N�¿y�="���BX,�mn�R̥c�9�O^��|̜N�Y���ֹ^��_��q����g�R}�~����z@$z'�V�g�qh#:��p�R<tϡ��&��UQ�Wx�C�	��*b��F ɏa1�R����y�ӎ��<�ۜ��E ��9�	t��u}�{��((�r�R��3�[�'�:�ob(k�}:�ҋ���w���
᳓g�ۦ�ǆG]�2]7i����Ikx��\�y��U��ƌ�n�o5,'�O�>j@�9r��	>�C�A�=>*���'�o�����T\�NmdO�K��ib�t).*AH՟̀ӥ�C�#���~:M�����.�y���Z�+��4g 7'9d��D�w{Zbr�da���=**��z#x�N�
��1�E�R�4�� �Ӯ����~��v�����.%/>�����\(�		$_�� J��jyX�ө1CO�|%�Ӥ�V�Ah��b�@P�Be���+(X�pp�������8}�z���\�|׃�'x�y,��E�D������oAgB�9�1���N�P�;��r�`��J��S�x��W6q:�]�����|�`���B0��VB� �G����\	|+��ˤ	������_���*�IG�h��7��s Ϛ�Q�&����P�ͳb�T���b�~=,o�F5>��^5T���
g��t�G�d�O��Rx􇰓VL�x��+{����S����A���Hv����Z��o�� SQZ���)��w-��\���* �V\dp�3Ք~����F�Q��۪��YTӸ�m��A�T�嶏���֐�Y�^��<��Ծ۾ɩ-�<%A�C�p�H2V!Na��0��g!�( ���M�p�F'����ئ1|����"P�m�/�,�y���Ȕ@��JD��ZM�9���%��~��W��,��^J9FX;9 MІ��`<��������(���R�'GC㪵�o�tX��߮�9��?�K���dJ̈́)�����;�l.è�*�O�T���3�,�c5�f=���@���.��k�7qP�\���XH�w�O"3��Wk��r���Q�;���=葆����zaր#�<��\Hy�;��g�?7�ށ ��h_OR��j�9���6�=�9�_��M�|͔ D�h����A��Dojv�{�0����Kr��]���RV�cr+��0���T�6�G�e�s���0`�f3�#�0_�o����?xD�����'xNk)�z�.$�3ۅ1��x7?`�:=�C��9z��=+to$��*V������;ƕ�	6yD�`.0P��;B�\:T��Aռ?1����3��ޯ�EzZ�O�S��=��?bfo���z-\�w(h��m[���j�:.���o͵Z���Az�qr;�#������Y�ۈO7������n���8�3T���lQ�U�<a���jA�@j��!��?��uqkS��p.^�%�X����Bs�[ۆ�h�M\f}~pw��t�
͜�d<k�f9�_�A��춰vo��dD<�����E.��ԣ�#p�7�r�7�qz�1��UI�2H�e:�_�l��`\+6O�]ܸ=RL���h+�0d��1b�966�t�c\�c��L�\����^��cUۄ�*���uu��ZMQ���� ����w��:\�UA��8�%Yl�BT֓S�z#�]����i�&C6փ����x@� g����I�-������T��(�(��]{/3m�YKhU��e����Th����1�f��n,F5>�<ܞPd��5��A��6������h�"p�M����wY6Ǔ��-�v���o}�O�MyXU����N27
V��aګ�:���^N汶��]���$*8L���>!Ub YUE
���w	Ʌu��R���O����P~D��,^.��J�v�<HR�R��h>,��OR����-x�O\��R]��ԗ=��O�ws��܋�����!�J}�/���Y$���DaD0��:��.�N-��jā�#˳oz�jY6�أ`�(7 �m�G >(��Y˖�Aأ{��<*�E�?�t�?ܷ^��	���_h�ۡMN�⪧����w�~�����|�P�h+&b�W�㠉+��*j�_QQ��U7*��33c��F��A�Z�4��B���({@m2���jɡ�x�(}S���)KZ��v�^S� r�(�j,i<�a�k���Φ驃�?M��Rj� �|���O�_0ƈg�/��ivf��ȇ�(Gfw9�����)���s��z�tv���y}�5��'���&����lxD�|/�9w��/=��ࠞ��	D�l�,��s	��ټ�"^�������t�$ôaPd�K�جX�(���e)�@��.H�#"�]�����Dr��q���R��u�h�;��|99�"���"�U�3��a~)��4M� h���(�W�.���F+���
=�1�%��_ɒ;��C_;CV�e�g�qq������v�.�;��	��S6q������n5�T��_��to��S�x�h��<[��n�m�AO��_�@�"{R��qC�Ц�F��ㅣ�4|ͼW���5C)@�@�O�R���Sq=�&6��"e���d��w�w�%��:�6�K�s��~�j�K.�<okB���s��VerAe{	�<��H-"�+��s� �U��w�):���/��OpE1�n$x8�{Jb��Yт0\^�8�j��0]����yA�F�5$�a�%E�V^!�~B
j�O��`tP�UIL[!�L��������4�`�-�(ÿXa�p�\/gqu� &��tM�;���ȸ��~a��'�S�j4��6�hJ�/7�hҭ��d�"�!�_t����JB���ꛧ/�yC'�K����,0��������F9���O�� ���W5>>�l����y��|�N|� �I�a�ؑ�$�ʇ_7<�l�W��EY�H'\x/���y����ȯ?�dÁU^D�R�č�?�i?��'��Ȱ"-�qA'�\�(J	=շ��P�<ؚ�t�<|�1M��"Ԓ*'fb����D�DW@��%�~�K���k���J?m�8P�ON*
��	��-�ֿ]���/��Ǐ6e��,ϱ��������4�	�
R���$ف���<:�	Y�-�� ��Y֬�x��+:ST���M��\2/�UPc�`E@��SG�u��i"�|L�0�\���K4Ӟ�u�U���3�+�Cn�f&9��ZP��[�Tj����>z6=�u��{I�MYcL�<�}���s�60|Vu��NmPM��c+�`���,�},&X�s�}��R)x�mܴ�Z$�d��Ƕ�4i�� R�T%|�����^�|̂��@1��jx�dI�߫2�uTMZ�l�D٢�mل���'����
�n#�W�5�x:̐��Q]B&^#MB���+�M�d�
L6M QlZ�0���'�F���0�3.�f�k��f��A�c�VKTY�+u�LpA����;�65`��2 �� �$�!,!3/�"��V`�z���V=�Z�WX�N<����D���l�C"��*5��nq^t��Hc���q�&��k�㺩�ˬO6�P�Hl��ר�,x�����=R�L�=_���z3X��p���7c�����R���;I(��E��A���$��Ǯ.r�$�V!6� ��X#��v'������ƙ5�N�0@�&������2��j�钉ӓ���)N;#1#�c
����X~�]'�J�2�ߔ��ӗH%r����uM*P��ŒUp>��~9�r8%��s���ri�G(�D.Γ�1���B�����{x��2�٨0�
��:�]���C@�_/� �6v2��.$G�S;��/����@����:�b+��B��Z�B��}󰺂�b�|̢��P
KiT�:�7Ƶ�5E�ᡶ���j|Y�����;/���z�/P�&/lF�W0s(��ߡ��(�z�O��H����a�	s�t(XG��R�@�� ������>����ڰ�� �"�6mu�{�#p-��҉��T� �*f�1Ý��#6�.E�֬�o�=�9�wv3{v&C?��r~�b�R�e�ub�}���o�a>����3����~���� �tQݬ�9��R�qs����h�.�1YB�Ȏ�k�?\��pA[��r�җDa��� |�2����Ι�g�Z����V�X��8<!t��D4Yio���"��fdM����*�	�
�d
��dD�@��-<�N�Tt�ׅ��r��}���o�ۮ��/x8�����̬<���r쏇\�m�O��V:7`c���SD�|A|�,ٸ���;�Ugf�/�O��3ȯU�管� ��Q��w�/������.��z�dϊћ�/øAd2gI����L�T���~cCd��5���#E+�_G�/�62����E�r!Wo*�wIX�����T\h [�$�\�v/TH�Y�j���Q�'4�,l����^I�G��F�M�d��m;�H��9�y.6�q�#sMJ�M~l凂�î#��ƿq�����	A;L"�v�n�)���, C,�l��R�E}�~@( q�2��j���gY��ܝ.$�r4����x����'���3�>ŉm���j�ю�;5�]MZ(#b64q��О�Rgc�ru64��&(��V7��&m��.�;4��f��/�^�0�������m�{��e�|*����"���ԅ"�ǭ0k����@}�k��B�-:|(�RG(�x����q�xx�_b'�#4ρ>��C =o�q�ՋqjQ���vPGCnP5ˑ�e����S�Җ�}���$}�[I�r&p��c��h��X�$�w'eCpXZwa�&���z'�*]�`��!	��̵����+*r"�֥_�s�X=���1E��5cy�&�`�)�b5g�C9�D8su��h.P�qNS��[�d�E�2�q��z$�s�j�W5 �N���ۇ�[�×�z��:���o]��q�+�a3����jmګ�|	����6�;�ɣla�����'O���y�b�I���M.�ToM���D&�I���
� j�q>�f��9X�6[ޔ��οo�.��Ba��^hZ4TZ9>��o��|B�lS�*��Ű��\��i�k���`j�eMU?b���M9ݤ'Pw Vk���m{p��������Se�om�v(@ ݏ��GQR��FA8�ZN��#��eWI�����(􁐯�5���bR!2�zU��=eI`���P/@��]4�9�[�~���d�D��F�HLK�~�ZM��z�������>���,��i��bަ��[����*�f�p�~�r�-�1���%��F����Z���@>�^���@�G;匴����ʴI�m�O����AD��y���.2����"ϥUD	)��w>�"ra���;�R�(��?u����&XȈ`���,ZPk��\N�/_A�?����0�1���7y�U������h7�w�3s+[ ��K�7Yt��r}.��IAt4���4�R1���X1��_�{.��Lv��}̢��kB]�)} �!jpW���o���2�V��XtD1j��9�k�)(I�ܮ�Nd!!l�@ p�G�D��A�3�	Q�r_��k�=�Db�u��+�~��}���!70_RX9�s?�Q��]�.�i���e� DIXF�h8_Z��	%-��;�zt����Bt������JH� �ܷ���Gg����
�U��iu��:�^.��Zz��ϭq9�k4�-���p�Z���,T����Mv��d{�[KL��Z�H�*�V�5��s8n>���.e���!�*y4Ff|1p�>��`A>�z3�G�g��fs�~�tY�[��.K=���P����!��z)hJ`<��bk�K�=�m��D c�+�ָ	��Xw��0B4�.�G�i���r�������(s�XE��X��ÝMP�(e}�@i�J�)�>dJ\m_���Q��m	6�HD=:��7|�~��^l�Y�^K(�ֲD���E�U:z��Tcz>*T�ӧo��\i:��~�~��:3|�F�k�d`5��/ !��X=�kZ�J�x�nU�}{�g7�H�0^{zA`��0e�0�1@�mX�Iř&��V�@N��K�E�|��X�2�nG�������@ɒ�����%���?�ŵ��L�{VR�Vؗ�ն����w*�e{r,�0#��R+Mi��i �O��x�L�ȫ ��^<� ���-g�=By��g���߈�x��!��^}$߈h�-�<�1-��í�R�&��t�h����wR#�w�ሇ�O;���s6�S��E���C�bfzhV�3~�`6���e�㏶�k���p�i�B����(�6�SF�˷@ͩ�S��!��ÃɎ�K�B������ =I$��!��ݥ��D��?�X�����m��C���!O͹�r�H�L���;5I}�NŞ���T0���k������~�/�9�}�3ğt�9.�	�L��8\�頓���3j{y��a�He��=Orv��a
bՅ���'�:E]���bJب��v�.��8r�`4�������w�/�u�:q눫�f��И���/���c#�������f��B��5'���}`An�+h�$�Æ"�g�̝���q���:��f/6j���|+3(����qM���ɻ�nS�,��:�L��h`Y6�
�d�`�c=/���2��7,ƞ?�H���M2�#����?������x��4l��z�զ�}�jye��t#�jM����"س�ᎅ��� (��Aa��wp��'���'I�j��%rsO��|jTe�iʐ��E�1��üO��7� ��`�F5�u��U(L���a8�,g�N;;5FBdM���i*	-
t|�)
F2�:���
�����e;�s����c�Ӏڑ��a�s铰5�M݃�v�|���g�B���u�Wڙ�3T�]���a8/����}�Q����r�a'�Pf���b��K2�F� �?I��F�e��	O�lF�LL��a؆h�gx=VP4���&Q�+�H��V�}U�!3`iiQ5e�=�$\?���gܵUv�2L�:��U�L��(��b�:/�C��R���P�"$#<�����p��h{V����D� ���:�xCթ��< jE��:7�J
�4�3��g{p���.�X����q�t�?>f���b��ꝯ�����,����ꔄ���Uǿ����N%3���
��1T�t����Li ٛ�d�O)��8�s��e�tX�i0GPk�dM�y4��_���C`�����7��#0f(��w�ѓT:]�3Hu��n6����3��L��� �-p�_A2l�K Y28�����ٵ�\�Y�]�)O�u����� �vN^l�!����</�4�d��q�n�@b�FU/����Lr��+��9��W���Fn�Z`T�9#2;`��x>F���2�b[sR9&�$2e�����U�r
���X�=�eO�_�M��z�,A.�Z�/��^T+���b��O�':��t��:�B+ώ���;$��;uj�x�<�8cۊ��]1=kU:|��~�^������5�H�n���Ҹb!��+�E�c��E=eQҴQ�m���X�������R�kфՄ��B��o�����7���+0-f���[��Vo������e�o�Q($�P�A"Z�Փh���sm6��k�&����D��L����v�P{���q�fꊝQ�V\ц�|633s�[����ը��l)8�J�˙��"筇J����ugd��BF���t��c*#�{���{��?�3ӱ��i]�X�^ߩn�hj�"����Ͷex�PU�'��� 7��8S����;L@�(�p;Q�+Z�F��6]C�S;*��5䍱�*(
����k��k�gz�3˳�B*�����n��bV�sx'����.�_tx�T��������Q��S������(���iɤw�d���30�\A�OkH��Z��B��_ ����H�K����~����*�n�o�A.�)�ᰬ9�ѧ� �V��{�Kdr����8�r���t�!���K2�f�����-yuk�]�&SC���y�����s+���MWՙ�x١��ј�����ۺ�7L8�w�����ϲPEĎo��q���c=���U+n��__]Lw�B��ܹ�B�M�UF�I%O}�������k��2!�F�< �s��@`ߨ�Ir'=�T�	��8j���ӽ KܓU��0|L�U@��P)K֫B�K���Cˏa�GJ�HO	݉�9�"w�l�H�����r.=�&zҝ���^�H�dk����`�}{��]6e�����2G<|:��lxk�V"�H8��)�&���h:(:�B`>���R2e	�{�Q��B̌,�.n�C-U3�������Oq�Yҝ�r�<� jq_��-D��{uk�skI���!���P�7K�$ �M��6N�Yn\u,+�j��.'r'��*��	����5���0}��(۸��h���֛�l(賀�]�o�� �`
cCJe�FҞ|��Ȳ��r�L�!mv��?_)��fn��uvF�����s[�uϽ�4_���
��:���R���J`��^|[���1ňq�jWU.,^NB��)>^՜p$�6����c�_۸}-=F��Ue�� �ـ��T����7pq[�qk�F��IĻx��2�ɆW�h+��.��s����4�`�Xnu,A���q`=��0֟��:�i'n���]��4j{<�a��I�[�-�~Y%ł �v.��d�Tz���Z;W䣎�R��/��J#�,� >�M����RQ��!ӫ�F>j�O���$/�%�
-���r��o����-
2׎Y�����'��G:|�]���R$;��;�i�
^-&׈����|�,^L�
'5��L}LO�,:C�D	�{`��̯�NCFű�� �蚱���Ƥ���w5t���.L�~�R�]e䉖�8Ղ�is�g$����f�nՊ/��,>,4�ʌ?D-��/�����g9K��G%~�6��)�f�Sf7�1�F����7���w��e�q�ܨfK���=c��sM����� �g����v��c�����fV�Ee�rЏ-2�`E��b��"�_!�%�ڦ��`�J�éQ6K���oN���Ew��!ۂz�`Q��`tN6��'-=89po1!.���DD�28n�b��RSDR��=�uw��x��*������;g�=��-����M�I�EQ�!2��x�Jm��)k���դ�qN9}zTĿ߼HN��*�q!<��	�"�"H��W��CÙD$�@#\�����3�PG���-��������Һ��K�Z��'�j뙭�nX}=
&t����OkĤyj��Ǳ�A�gʇ����'�#�ބ5�j�I����$�yM�r�3����������kv�x�^��'�^��tꑪٞ��\��z-���`;�jo����pb5�n4cE�L�6`ȮoVulA�o���t<�lCl@�OhJ���V|g�j��s��t5#�*��'��'z����XM�8�j�r.���@y�Ȏ�̮%Ul�	Y[,�zO���&ī�T����y����^H	�8$��Q!L%����]�u"�
��;��84��Ԋ�@b%)��5*&3�J[�OTԣ�RL ��J��y5N�Ý�_�S���9X5�~*I���� c��)�/�[&�
��	���yJ�]
�/Ľ�b���s[�A<��mzX�KƩȱq(
C2B8;��Qw�M�59b�Z|T�pF���U��N���SyR�D��[�_].n/���a ���s����%p$t�A��
s+�W�wc�o�5N?I��f�g��_��@��XZ��DC0�]|Goo�C4����(Mç�hkb��oGe��x�sX���TJ�q�s�3�Y03$�����f
�^W_�:��]:V��/i���+���ь*�����<�ΩreE.EwY���j����R6�nxJ�wa�������05x�,��<� ��Xo*�N�I����⦽���53�zf�=v�����a!�d��3���(����rⰍ�ҁ#�^}nPvHaaÞ�;�>֩��AL��]]ڒ̇�c�8e('�ȢՆ��?n�#�3�d�3I;Ѹ �.��ܡu3ӆ�oBčE�]ʙ��]��֚�E�\�q?k�a�7:D�A]����Kc�����4/b�ܼC鱤�y!�)�U%���(%^Th��6x��Z0�w�cA>摋����P��\�=Y&P�{��O*��U/�k����"f1/I-��אan��߆Y�GTU��I)�ęi-`8 p�(�B#
���@NpV'��/�{�Msļ�4!��: ��o�]�����}D_�P�:՚���$d`����D�A�Z�Œ�?`����V�P��������>�3t��c"mܡ7�Pش7����ДybFL�㠧�F-C^�Y�I;�E���T�4���؛y��d�~�c�ą�`[���R[AN���"��B�M�)���Rp�˯��<J���pq�{��c(D������$��Rc	C�s;�p&����9�l�Wr �~��3NDkKq*�@SYvؤ*G��N��_�Q���O��v������>�rb^]��j�A}�l�]�S�@4�{-�0ղ�	Mu{�jg��A~�ϊ�ls�6��}ُ*�u�V�A��3�G�^�>�][�p�w3���Lwz�"��t� ����1���MPBB�#�}GEV���aT�2u�	e�}�i9'�'��Ay���'&&�*���� �>������?�i��6�h�\���Zj�jsl�Rכ���M)�����mb�S?�#��Ur��ђ$n1(�����W�#e���(vv�;�qxd��\d�Ώ��	vM�F�J]���������|^ܗH���vײnP��9��ϸ�d������� ��zq1�4Ձ����������_��2���� �4��2C���/���V���\�I�Uyҳ�V���:��r����kI���6̷�A ��,����ف(n8aE�k��1	�Ƣ?���WU�6))�ո������N:��m0��
�t[��*�i�P9Y�����θVh5��L��7f�&`�PV6R�"ޞٶ����M�2�#�ڊ�z��I��Ύ�C�� |%����WN�Q�M,�9��bp�KcԴ��$޳[q�B	��8a�)���?C�v+e0kl�	~ͣ�cr�Y����	��������y:{F�Ԧ+����G�~vB6�
>����'p�"|�J�wrX-P�;���(�Ќ��˖�h��C���l���������W�{�G.�C& ̦gO�ޛ1yA��� f� p����A�3;���
�(q��� ��_��g��Ryd�b�����1�D{=����^��W�
���kP=Z��{P�����;N*�c�P:�gK ���E0�si�������H�"&��gJ�a�Sh����AM�w��!塚�8$��?�7��8��hغ�z��w�u"�*�ѷ���W���@q�% 
8ǲ>���O�z��c�B���Q��BOY�x8\b��CU��*^�Ϸ��:�x�׵[WsY<������f���vh��P�o���m�Z�v;D�����O�ޙ���5�c����g��ur�6s@�3*��l;8%h�����2IN1�y�A��
�CA�z;�35묯�v�����$
]�.?���S��<�k���5�`]���D�ٖl��i?�N�Pș6 ��Lef��,�|WHLO�x�I�UT�1�H�L�F��T��Ȟ*%2�Z�CʚnQ�F~j��H�8)�}ʐՐ��s.��}�#k��[���jZ�~�o��;���u��s+��]��I8�۵A�
����k�d���{Zg�u��26O�9dk���ێ,X��o�6k�3I�H���4'�+!yև8d[���|6���$�tԥ�O[Y�Zю��j��r�8|�Qc�G
�j��9�	�3������'7�J|���Y�ތS5��U�u/�1�t��5�]]���v��i� ��F�ivV�1	֟�)����! z���@8��yދ��o��I�7�H; �c�g��{Y�'t�_r�'��X�A(_�UY�
�0�]>������9�mtH��0�h�6N�\��x��%���wc�@C���=���8�v޷�k�Wh_'"9vv�2�ħQF��Z�nq�]�muz��җտ�n�9��������4Ky�ʬ}C�$VAR��I+wlc+��\�IF5��k�A�)tkRai1N����R�k�"��+TU(���aHsC?�y�����&ڇ��6�r�4_�v3���q4	�E�SJ>�
?#;@؄C����~|zD&�XU�2�^p�/u
Q���".y��ZO�`T�EU�R��r�#䢇��M�����(���Ogk�J8cBY��ox�������d�66LG���U��o�IH�)�㈬�O"�y�R�t.����Mg fK���1D?I�l9�{�
>�!U&����-,�SŔ���>I�rd7 N�2�#�Ѯ�wh���#穡��6��[�O�_�g�R����>���&^�0��Ŗ�-L��
m�H�8����M��	3��KT�Cˁ��bR��1�1 ����q�ء��]�>�5�H��w�#���^��.T8Q?���3X��[O��\�?ARf�	-��1��� �i[$�+�Re��n�/.�
�Q#	s'Sn��O���.\�0���{!�\t>�����c_ϡ�49f�0o^��o\��o�E|���7j4�$C��g��>���	�ˤ��&`�s�-��-'��~�t�����Z�/N��:Κ��7eZb=��JH?�3!R� h?�$��\���]]��_�S�u�^�*B_-�y�6����޿��57��a�!W-<xN^l����[�k��������{3�Y_wD� M����D7݊���0�oӛ���W�K�㉫��p��˙Cߩ~�0���&#zj@^gt��gw��L�ΰ��Ⅲ(��Qʭ8��Jo�yx[����h�M6D��·�<R_�0$"��Xw�޵ �nNm��]�C�������H	��"�s~e��\�&��^\J݅D�������B~^�}2�f˧�1ɺ!Q\��`p(��'١���/�E)3/=��5^����
x�}��M ζ�Q�,���
m���{_3X�,Z�\���-$jc�,�p���z�D�v���j�6�g ��gUT����l�e�9
/��H�ЫmAmuQ����qs/�哭����-���ft�G����z}<Z	�=7���L�(�Xo�Q���3w���`*ox��q׋�^`Z�VW��ya�]��:�u�_����Y�QP�"��������F�_'������:�k�M��C���i�-�^R�F�1!���JY��jg���Lt\�t&6f�_O+�:��Nz�q�<F���Wb�6��q˺�d�{�������DB~�]:-:�~]���1莡�@E�n@����r���=�-�׉]��^9]�6TQr�-Y-�|5��,<�
Du	/p��8�����0��4��OI�Jc������A��L}kݶ��3Z�ȄiL]�%'�]��V�ⳍ(��nE")��ȗ(���ޭ�ڊ�DvL͉t%
^̴:2D�����a��J��
zB�23��sm��;׉�q���۠
U�^������R`�L�obu�Eل�,V�����Ӈ��0�`Wf��$�HܫO�� 0�I�{��.�nǠ��{��JB��4$\"2*��H4Ղ��6�Ҽ�c�u�N�W��t��Յm@��2/M�&+��*�������P�<LUɱ��5۩�	���5|�`�9��g~dNҽU)Ijfo�(x+6�R�8����{�/��`���S*�O��|OZ��=F�}�8���f�������tk��T��x�wU���7���ďQ��˄��:`v�=���un"��&��LG�-X���W-@S,L!M��p��=q�J�lI�&Z�q��1K������H�L�_�J�T����o*7���_�#-gP��JY��d����ב�f��z�n�U�A�`�T�Cvka�0�
�v&.��A�͗�/i�j���u���=JAs1q�P��1�eM*���=�r�f�eg/�f�ʺ럡�x�������zܣ�
aԬ����(s�4.�O�YKS.�� ���ZL����l��R�"���I��	װ�mX����ɿ�F���O���:*��%�Z\�F+��v�t���dԢc�Yv�f�{m�s$�S�v9�B�JY�4�f����
x�C�$\�2����&�}7+��
�����C%5w9���n�B�7dVΏ~[���n�8S�c����d�/ǅt�j�iw��DO��\V��$4l�KE�E�:�>����w�ix22C�*O����_}�<�e��6+o�顶x(j?0�t@��ɜ�S��4��F�^��wZm�o^������cH�k9�Tj��(%r߳���7�ց/��~K6�����S��=��(���P�@���]�M�uo&CkZ�
g�.�`�ӕ4�;g74r��4��4y���wb,��"�YG�+z�!Evl��$6Ťa��U���3:`¸"M�c)����=�g)/�fKpBK�,���+(�u%��MzlZ8�)��z�����Y�@љ��Ɠ7%f�����C]t���4ԏkw��DL�(��(�l����F^�3�L?NĤzn�h�)�G�|�bg%^�yKX�������e��D�z�)���ķ��ߝ��׈р�T������kA���bf��N��cⸯ���/���@��0/����j�֧W��<E��;2#�O�:oK��&��V
ə�ѕ�@��>����h��I@���q��((�}[U��A�F���6�1�*a�&�3������c�/0ɃXQ����䵊/7��3!I&B�x�Eg���_��0b���d��tc�j���"aR���]�Nj�m���t�,(�\�K�*�B�)	�9�G���U�� 0Y!�O�}�o�Xu]���e	�݌;��	wٲ�l2����U�qVQ�
�<~�B�����1�+�C�f�p���!6�c��7͉\��z��_�}�U�Yq���_��!��? ^�g{��']A��\A5�7�Q�~c=2d���լ��Lc�L��=�@�WS��o5��&�Ob\u�%��]�೤���q",LǛgJx���y��	�
6�0�c���Ý�;�8+�[f��T��CRYu����H�����S�oy���K��r�8N��N�ߝ�<�v ;pkz�hP�5b>��y۞��B�Ðih�� ������%��d_��O��'�wK슩��(wP�����>�����D�X����i�8w�u�dX���ޏ	�l!���`���ʨ9�I�z����6�ܟ ?nK[N�Z,0�C�O$��ur�v,�]�D{�:����9մg�O�8� ާ;JӪ`���n�SW�ܞ�2��o�;��'g�?�<.��g9�{�p��	9��sj�����W `��5���SY�#Y�Nc �J���v�S1X�tSQg�(�����[-A���h�s*X4���F��>t�4_xu�ç{��Y�YAc�$��9NH!H�� ��	�@Xx��K������=G�%��m�F��E�:�N_�?��:�U�Νcs�EՕ��Ե������ ��x���ʴ��/�E|��^�H�,������a���ő�w�����8dL�����UvF��wq�"m�E��P��!r޸�솢�ٺN��͐I��5/X���ϻkox5���e$�AJt�J%��� u���9�5�R����O>_�&Uz�ڋ6����x��W�-����Nʬ�l�NpޢjF8����}��m�!תcE��o�Bt��e���o�0��J�������y�?_`Y�-�l�i5a�q{��m���FR�d�~+c�.)+��pww�7�X])��=�z�5BV5�Ɣ�p{�Ƿ�ŏIf�%|��X�_��$%��+z(����\e����ce�g,̄>�d��}������"y��J_�[�����X����O0�_l�&��r�&c4��F�D<�#Nؗ,z@�cQW�G��w}q��P���s��挀�
x2���O*��F�Ts��'æ��ߔ5lƈk��n�s9���-ϑQ=�1G��W,l"T�dw�%R!���ފ[���(�^p��Gj��f��0�s�i��),�~�ޮdlJ�����v��f�L�xꊽU��HO�V�>NNM�m��F��pJlE���X��읡��9�س;���T��XO�#�3W�y�[Q2�Iaz�՗{p`q��Xa]q�btU��9��L���X�v�5�Q���>�J���4&���}�}���>�n�&��O 1�D2P$'�ݳ��K�(���KO7"���^] T�v;P`�V�yd���NR��Z�v����/�˰= d�R��.�c�8r���3�3�ܷ�ߴ_�/���\��
� L�jGJ^���P�=��ʻU�;`��I*�M%8W��vz�q����ϒPP�
�
���C�/PK���8���/4m�����/c!9�ʜ�54P9ǌD���G�(�X��߿a���Dx�k������a]s���U�q�|��yй��$��J� �~/�"$��#�8�c��ܱ I�z��"Q��R6�H���o�^��~K	>��^4:��ݍ�O���e��"��l�Rp��Gc(W��V��+L}�,�,�[�g;�/��+��þ-��ȑ���P�%i�~gE�R���@��O>:�m��n�~�4
�Ҷ1�%�T�(Jr���%W�mT��Ȭ��D+5��:��`{蕶m0J�M!���!ރ�Ҥ	�).sO�	�0&q���B�l�%u[�}B"ωZ|~�%������ɟ��u�6r}����%�4�%�=��$��3��2��'�X�I?=~���M���GZ��;��U'1�ˁ�ռ^jc�3��$,!���d�Շ�Ǥ�+h���N� s�r�ǻ셪���9pZ��%oJ���g���?��'�9z,�ɵ��@�r��h8��蔓+��uCtE�X߄Ih�j�|M�7G5�"g��T�ޟ��j�u3�`�䍗D�������hR���hҸp��P#��F��Eݹ�\W��ٿ��uT��o�b���˩�yYC������� �)�It����6��G&�93�B���:�Ӽ\��EUW��%�^]ݾ^��{L4��MB��(�M�f���a0�](�0�����gH��ֱ`��!ti�5��B���r�����#��Q�:��lZQ�u���pT�'��{ߘˠX����N.��a2�)jeg>6x&r�x�BLC��I7���}y���7'���m³1�����{�A���K�#��F���,KR�>( �`����A�fg ��r��є�I����������g�Ea����cr|���(�6�zW���X�dv�[�"��P��@#Eت���B��K���Zi�?������dd��4�Y�' }}6_�O3�Q]�̴5
���ױ�mm� ���a��w�G
8�#�p�[a����_�O=3��NvƁ';�	�o{��q�Г!�%P�ӑ��|���M"�an�.�"�~�h6��~=��
Fz�K�Hↆ� ����*���+B��N�G������o;syim�<��ۗk]G�����:���F������Ҫ8�H��Z�݌#���֯�p�.A�G��&(� ��7�4�$>g��h݊����E��ℜ9T0�y�zk�^)JB���$@Z���Ȭ�<�<�#�[Ĩe�*M���Ma���gr�F��6�Hn�}}�.���+7v�������b5��*� ��gw���Z��Z)`� ��M"XL�Ƥ2�DW��~N�pы���z#��������0p�:)�@t���k�Q�r���ۭU��o�#�����_���T�����U��8��/�]���W+�֞J���5x���Y���d7���go��TvRX��:�g��<߯�v$�����f�^�p��B�$�tl���n��W�$�4���ˇK�`��̫S7��!C����r��M/�̟�I�E*6*I����J�,�U"/A�7l�H����N+�9^��y��9�8�1���<Ґc�yM�_G\�	/n�+&5h���Lq�gw�J�s-���EAf!N!�b0�)q�gU`^.����+ǧ$o�'ڶ��C���J�r1W��jtJI�r�O?���JF�m����b!��X�RU5<���z: ��͞�]%�'#(���p4��'�S��K�v��;�A�"�m�"���@�}=W� @��<�{"��(�>�C��~�eMU�(� �x�˅A)ūq3���i1�}T`��`���e������%tKi��@Y#�g�{�Ŧ�D�Z�*؎.L���|��t:t�gE�o�'�����B���@E;#��0	�û]��z���8�l��*W�Tp�=�k��<�GĊ(?n��{��ؤ�V�bHEA���*�1�|F��rh�=��y�@�TE��1����?����3'��R�?��w�7��|��2t���o_����[���"E3���_j��i���<ɔ`MIT�D������
�@�|W��&�33�9H���d�v��Xp�
��$��R���p8_�N�ϡ9G���H��m��s��B$:k9�O,�l�Ak��h��o�5��1ע���>���;����ԗU���f=ZQ� M"y���X�B<��H�ݸ���d�'=,T �@�>���u���,R�%WuU�S�+c��Q�c��D�����K���]Y����Q��:��әf�i@��p�P]Ac9p�Dk�D2��0k�@��������P�����Ե���L�䲔Ś���@����5æʍ��3<�$�W�单X�рf9ʚa�q�3�����#�~J�ڧb�X���m�v@)d�Ʋ�H�	܏��B�9�Y�=�ni��|�����".�d�2ǣ��Wb)~�:io&-��g�i݅��兲��ؾ%��,4�����8���ڲ������Yh2���~B:�A���h�r�T�Kd��j!�G/��K�Ė2i������e�s�M��p}<�,":�6�'�2���3�{��`Q���q_��R�`��LF;1i*uT7��'�������P�������\�U��C3�j�VWI!��G��)8)|)_��Òʢ�S\nuk�KY�A�P�j
��:�")JԨ2�(��b4'#GB�ix��%��ճ[GW?
P��Ъ�����*�8/U���X��$х;q�	�����1���ds���}����i�6Sv��uǜ���
+�Ο�QƘ�AaXhf��pܸ�����)1!��I��h��EG�s2/��UY�&}�x��@�{B�^���cv8l:a��k�ٯ�q;E�e2��SGF/P�қ*���N+%���ťnb���.�b�g�4�̫��$б̞C���f�:Jޤ�J���6M$�,UC��Z:Ț�z�(D��|�IE��X�ʆ�k �uɮ�0+�J�=\�s��אak��ۑ삊*>�X+>��h��ȿ*�,�U�/�E2�i�2Fz.'x�ƞ��΋	n��K	7�I<�[�'��i�$z��{�_'3��K�e4��U���`����7�[�9����ٟ\���3���j�������E ��9wwe`���e�4y7���.ۊu>����H�0�#>Q�
Ug���u�j�B��J�w��꺼:����c�d�xb`,�	Uc��{�W��=���Egll��S/ʎ�tA,(8����4�����<�:�8XG����r0�n����!HA�����mFW�!�p�����S~�	�*!�����D-�!�2ȷ�� {\G�s	�4�h���f"��u�3 d�-�o��74l��k��ʽ]61��J�C��I��d�&AD(M�=	��[�m"~g���I��Ѩq�L?�HO�-T�t�<��!މ��%E6�^A�k�?��[N<� _�g�Lh�Ĥ�*����`�HL�Ca`��<��7{�2�A"o;+l��U-�'��Y`��]���j��w|G�Q����DqbHPy�+��ݰ%���-�U�/B���5��T����#��F�,�����V��P��錥a2т���W��Ե�?�P�8��_��o��$"���;���f'��Y���^g]l �*_L��ꥃ��/^���@����t���漣*i�2�>�Ko����P�U�$�뀉�Y�ˉ�=�d+�v�0cm��c����t�s��w��5`=I����rX�Ԑ�Q�*�}y��w�� ���p>[�	���7��ً�i�4���ȖK���Ȋ��0W��Q�+'ss����2J�jʾ��rS���H%]4��u/��	T�I�w�hx��Adi�0�S�=b��MV������wKG���)�N�$Q 􌚲�2�F��0Ȱ0
��$w�m) P$ m5�����]$�o]O$	:��~.+�"���۞�ўru9�g���*���Y�E�Rt�A�x��``Q/��$mM�e�J��Y��RēdS@��Qׅ�k�� [�����LF�S|�}�������ME�km��e��'rd?����O�렽�(H�X�D�W�aNo0��-���9:^����&qs#g�a�^ إ�vv������׋�à�D=�S!Y�OT߾�������֎N����xr�n�Z*^rE-C�1V|�:z��L�fȢ5������YI��}!f��m=G�l�V��!���6��K�[�B!�J� �+շ?H#_��?�.��� 	(~�S��?�c�4i�)�JM_½�g���7}��gD�`uc��̦�B���#��F�z��c���i��`�Ix��Z^s�D��I�E?��w@�'���֒
� ��u1��"So$M���T ��D�裬�e��*�mS�Z0�}��
�iߘ��˧�B��8�S���n"
߆j.�xLh���f�7��p��Da�+��G�
vO�0y��#f�@��2úF(J �Y�,�to�{�M3�0n��)�_P�<�\��֜5�CU�Iمc/�^6�O�*1Ԙ�#�|2ᘥ*�}8��Q�����jԲ{JL���p���cKb��,���哣\RߟDm��x��%]���Y�Z�Q:�;��kh���'c�z]�̟O.	��;䧿)��2���K`�];��y����CSI@��Tٍ
�NB`�����BsSv�&��26�^g�_��`!���6t��8
!�Zw��r��i���r�xJs��?�Ƿ��Fdu�����_���[\�d4�c��Z�p�v��H4�%��H6�:QZ�yJ��hj���O(���VD�ct��"���ID��[O8`���)��S��������n�T��T9.b1PE��7<�L^�1�����hƄ~��P��еF1񭙯�]��,+�{;�����x�P��U�Q���p�2?3eb_8qu�k"��A(PCnvU�DR��䭾i�^�ߊ*�����Iq2�B��%�378;�3v=,c�r��o��^�a�A�%�ސ���X2�-,H�U	d��0-kB���wK"򲣵��&��ϯ.M�-z��}��3����٧��Q�����Ϊ~W���)隑D'U�
�r�>/p��z.2Ыu� ��01)�l׻��}��*�@���>PFbґ��g�'�ԧᤈr��:"�QC-Q�)j�.����Kэ�5�_��i��
t�k�C�oc���`���q�ٟKG)�)����Ț����P{�-��x�Ūv���*��f�ڠ�� H���?�^��*�_b�Ul�[���[��uH���)�=�NeS�sJ����6t;��E��FHَ�mJ���������F�^�hNMN�4�h>мm�&Q@��AOtK����ǟ����=������7�N�����g�I�5z>-��`d�W����3�K>`����0j����p9VC���}�*��DB!'L��IHV5�E9<]�/�R�� !��D�Ƀ�8��;�[Is��3�~;�2OI�s~�0C�P�x~�Zm=ӂ0���m�����]�x���`����Q2đ�`��YaW�z�ya��e[��Y�?�*�:����+ʚ�'��ZDv&gߩg�}����̽]\)�L����o��3V?{'��'�cd�r� pά!=*n�	�����16h��`����i��T���/F��,;G�	/x3��]�&[;����
��	����q�˥=�J[�F�H?�Z�/��j��A�a9�I�}Nu��}�$ ���1�C�VK�$������x}�d�z���J�z�%�v�+WZ�6��9)�{��h����f�24�;{��Ô򽩱� ճ�NIM�^s���c��3�N��P5�)Ni_9IL�J�G�V�=k�V8:�V&�2�Zz_��s�.�t��Q��)a��f�B���L�5/�9.vB9m� u�A�),K~�y��#1�����EP���3F���08�vrF87$6�άXقҔ�;�q�aK�Ԁ��?^�V�qG�Tf�翫��G�Sg��=��X@�l���°�XI��YƬ���9�̗���E&��cFX����!���`&�D���L�&+��9�G����P9V:�zs8�F��A�XaiX�m@ݭig�8���L6�0��̲�\�÷���M��3K$��gEesm���nD(/�PG��[{��N{���Y|��J8:8p��>&�]��^��AD���Ͻx��y��CT��V�|��|�Nm�a�g��2�Z�ZV��6`����3nS��f��|'g���Kc2����f������Y̐jXY` �v�fJ�������(�N�i���T�u|��Sk�k!C��G��ڞeת����ū���n���������K� �O֬��q<2���K������
Y��< ÌPF�bc�i0A%�I���[�nH(v��t�oL�Lۖ�|��X���q�,�CF������*h��+�B7x^R�3	U�I�!;},ro	3��������
�O�V�m��y�5��f!?���S��.����T�9l���I�:��=k���H	)f-K7�k��qgs5��/�#��1-`_�A���j�0�L��B���q�	�u;�
U��]�EiU+�V!Nt���������۲�g���,��>9)��H��������ԖJ��!d�9#���.}و�kf�{���*zG�:+W
s��>e"�x\/�������(��{���֠��c��2��� gb!�i=�2�}�?��]��E��=�4L��[�����t1;��C��Ss��4蓟Z��\���[H�{��DK6����wJ���(���r��.�d�;�<˘.��l{o^�<�M:hzJ����h$�'29�Ti�O�PcLJFO�,*��|��h`��|Ɠ�O.��o�2�g�.˥=�&9�?)���gv��0h��U*�h�خ���/ϡ2X
d�)�(�ޙ���[ PD�A�����P7�H#|P�O������ڭ-&�e�$�>	�)#�*�O?�b��<�E�~�G�H�ђ�nH|���"y;�1|#���DZ�G)Ͼ�����QQѭ'Wf�^PzI�ܖɒEy�f���:�-����&^��A��`LF�C�_U� :�����&f���^m��60���i��p.K)@���ۅ��R$�"I�P�[��{Q�Ɩ
n�J,�:.��p����ޥ�|��U�S^7v�53(���F�89?�	��&���[U���حb�0p�N�-�S���Emo���O݀�Ί]O�Ɵ|�a��Ж>l�%�;C_��� K�b�?S��3�Pp���m���!����!0�����\�쒐��s֔��_JX�*/���muyn���p���ՎG1TR����RH5�4��Z�f&���I��8�A|a�P�/�$r#�Ej��#RJl����%��[3�a��ݹ峕���c;�$�Si Sd7l
.<� ��#Y�{�Xi�-�QaJl�t�ݽ��if�wP�F_ff�z��h���r�K<j��1 ������p�Z�u���M���8̶`4�I�.{�6 V�n^[H�w,�cʵRB�-!�b��;��?X<��x?y�U��=��{:��R�M���i��,˜�r�
8|CГˊ?iF��v1�g⪵��_�޶��x�EL-�󟣺��1.R��m@��qe����m�9bcl�|�܊�|#*4T8�[>8`z��S���#3³V.Y�C���:\(��(��1m7Q_X�"�`&���͓����.]zЂ����^�7����t�i�liC,AX#?�"R�<���}�|����2n//�:KT{h�y+lwHg�ۯ�Y�*�Ȋ�1x�K��mƎlP�a����Ӂ��@Yo<	�n�:6�9����ٌO�&t��[���a��n�W;�����
[�?�{�P�Q�F�45Kh��7�SN)�qZy�L�g!����I�[��b(/����p�>N�E5��MX��(���j^�	��������Y ��6E���"�̌ N<hR*Ht=ԓR�:]���G��B�h�׬TI�U��l^c�S�Jp�%U�Z���{�_��.+���u|�G�
R��]❆�eo�yf�}�ԡ � :����Nkoz�;]�B�sM�5����Y7%2��}lIB�Iy��
���1s�u����y�<:˗��6mAKf���n��nhŧ��|c����ʔ�%b��>]|���V7��5z4`�8
T�\�����웥6V��S�����B��~����ib!/\�.Vf[�`��D+�ÎA�W�����HX���z����b-|@�lj�A�4����X�i���7������}?j�1�<Z���/�n�;m�O��{�������1�ں��^���,��k�ԓr���i9~�'d���?U
?�T����#9�9���.�JY�V��p�K>s1��\!�ě�a����tYH��y^�wK�0[q�ط�3�U����2⣒�<M�������v�	�XM�4��j�Zٌ������ݜ+]�w	OsX<N�S*��T���R�@�S_��Ab��x�m�}u~�g���Jf���]��w�T!�2����7��-��z�,����p�
������0)s~���h;# s>9��e#�I��⇫R����O�(������]F#�"��v�}5��P�ݗ�||��	?�`L�T�ފK'�u�%z�rbb�p_D����X��'<�Ĉ:A�#�~���Z�	Q��	8B�直�6�28Ud��R�fx�4*�Ȏ���}�=\�<�D���K�� x��1'c)�����g��2�����V�<�dM=n�"wKF��,���ca�לwC�撳t�g#@�1�SV"fŶ��TX"��rm���HƗ��l&� �q2�l+�z
:����<�^����.$�N����6�oΓ�ʏ��׋ph�X4����>ʡ��J!ǣ�n=\n%e��Y�M�n���t��'OC��U�-ً2̳o�l�����s����̴.��L�_�s�x�@���˂tQ�݃]=�pQgk���n�$צ647xvO.�Dy��g@�z��&����k"�S��Y�p�=�\缈�N�'(�OD�>BU��.{s*���P��J��r�g;��[V��LnA�H�e��o�x'��%��E��b��8�ĠT���θ��(L�����ŵ"�I�I�u�Zm��;8�l���D�:�\�r�E@�N��wBD��SG5����g&�G>CP��9�3������R�  �*�;�/���v�7�<�,��^@PP �����7J֣��s|�&l����G��#�+-�/��ê�%�ɧ�.����Ī�o��������C8lrDJ-�^�LF�D$M�F5�)��I )
Vx��Ђ7�E*�^�)��j��M�i���nw���OQ�����q�����)�E�S����N�Y&1���% n��ZMxUo��kD�F4��DluY������s����"�j��`0�}tֶ0���'�aD��N�ۏ���=#3���6�܇R����*�쓶�rIì\nM_��(���yɥw-`9�׭�@�T�(F�@�h�oo�8���c��0ß�d�%�n06���G�kc*U������=sm��k7���5ی�C�9[�a3�)6�l��1��67�;����VA~/��ezn�m��Ծg��`&b�Xz����z��{��9P��Rf*������1r�ʉ<fJOd�����}%�|��0��ae�[ pͯ�o8*7_��|��	ʾ�d�#d����(u�YU�"�eC�P��H�M?����:��Z<	r0�|��C���	v�{g�_u����]r��ܘq�;?��~	A��Q�	4���<jؖ���P5���E����M��a2�В�Ks��2nY�j DQ�Bbr��ezYid�����J��Mzd�ˬl#�����0�$��R<|w��[��3�1��r��4�ѝ���C\��G���D;59�([�㐪���D�����_���P�ug����p��
A>Y
�`!�f'LI�*W8"��=q��B̌���|X��ҏ\g�q�^�}{6��o9x����Gb6G�+��!�l����򹭑@^6��Q���h��S|W�$��1�b*�" n���F��J%��MB�O��CS��ʝ*��W����=���	�'���R&C�ʻ�I���H>�3�����2���H�>���POmV�m�E����mY��;,4�$5���z�W���4nF;�����g5]�����$1�
ه"�H���������A�X�_�^x)A8���À��G�Pj��Ϡġ���]����&K*�q��z���� �d6`qŉA$��f��On~���+ߗ����έ|�tl��~4�3�nA4|9L�*����좃Ё���گ{�1�$~�ȼ��K����Ϣ�E�Š5m%�9�A���E�L�#2;��go���E�޼){�̰����C`s�BAB4�.]�P-��U��aF;��F�UA�v���ld���D7��W	[��r̞��u?Ȗ�8�#
tX-�6�,V2fӕ4�Z;���NC��p%����p���y������}���!��sj�6�ö���u�FGЋ+<|Cq�}�� [�=��	n1��]��J!�8�U��ΕYɽ��c��(��QR��Dܲb���)0y�^�����_��g����
��X�m�C��i]��HOn�;��ޅ���L6�6Gi�����|tIO��xX���ټKZ������r�����@^f���%3�9�J�G;��)xE��5��xdGG��#F�N	N֋.�e8jiQx�/��lAfP�s�����lI�ή��
��+�˟�o��8�^��Z�y���$ra%����|�I���T��@,�N��u��dh�x<�2գ>��Cv��%~�P�(�^��P?�\Fo �8tPGQ�Č��W��kM�n.����M*�9޺_��൝CrkX�z�{L�̙�(E�O$�ɚ��v�S8�Ge���$Z�
ꎻK�͏��i���H.a�%��ly�G6��(�gٔ�"�ۈ~(����Ӊ��Z#��O�/���#*C�^���ƃ�҄?���V��"�Է�5��t ��dpzy����K�9�O�gn5N�
A!���@�V#/�Q�j���<���[��!ܪ�~.`�o N�h5a6}}��=����v6�f=��km���N0C&�Jܭ��r�%�iL�c�a�)F�Z��X����o�U'�U5�N�A�c��Ƙ'�t��Oi|Z�׃��+���L�����#M���6�PBp���
�EO ����EU���f�U���pe�X�̽Bi�h���QV���޳���Qa�ə�Θ�n%ܾ������NC]�Ȅb�a ��]w������=;,}{$r���[
�]��8�:�?g�_�*�4`N���-�q�nbfܽ��M����X�?�:\�s����!7fy�i��E4�_saYp���oJ�-80�?�3��Y������$R�#h��$���稱r��x`ݏ���:_&�֌�(�Y$�qIjD�C��(���f3�؂�C�#K����ԭ(�/lh����A\�)+�A7����I2G��OՏ={�".m����mXW��h	�r���X�����p��Yj)���.���N�;Վ9��Qn�<�Ag�W��X��s��n���qL_.G��Q2�]�r� @M)�(����6(��ljL�U�m����E:�a�<��~�-���T{M��jG��׉�~����6�5x��r�?G���,�o��e��C
n���%��!+��;��?�6ez?hW<�1��P��t���B�DC�<)��c��$���D*,���!�:���Fo�ǒ���e��>���W�<8��+��$�I��.+�8�%��U�7B8�jR��ٰF?[�9�k�2��FVe��xĞ�;���,"���`?a�&��u������	(jS)A�T�C�8b̳o� ei-���8aG��~ƴ��ŵ&Fi��zm�؋Pɒ��dP	��P�Jj$f?��|l�����񃱧���b�d��a8ڴ���Aw]Ø���y,�Ů,߭�cp|L�W';�Wn"մc��!Ɍ��Y�H|�O3�V����T^���*(r��1��Q;]�Su������S�1Bg�bb,禵R�e�2��e�3��@▔�+k�*��L�^�m�
οBO�5&~_��G��x���%K���y�99�^�sR�a��J�95�b��3����텈�z�|2��	�Vwi�M�$(��Ý����)�\�c���~��⟄XzuU���׿*��J:*�]:]~~V����w�L���l����f%�`�x��7���䌓	�/0��� 4h��no����x�����:SӨ��Q��<P�A��D��deF�z)/�jYX��(��/n�҅B��� 5�XT�a�G��xˡ���U`F�O��C�؜DUh�=t/��S'@�^�)��x�n4��N2��N�)�����KF�\��h.�z|�6_G6�� T�*I�Եo�B �p����O����q
��r�]Q��</�O�m�G��.q2uÜ}$��N�"i�=)����(�s��P��Ν(X���J��?"�U�!��{�r��O>AUid�.M"㖲P�7�9���{��j�H	R�rj�{!���=N=�Y�F��,���P������Aә
9lyZ��4�č�¬�CX�{�Y'�Z���)�?✜�5ؔĊ!O���v�A��J�BT�-�:����N"���S���Uj��13;C��'�5�<�W���Z��Xս�q�z�ə�h��C8�X�)'�(���3{�{�����.~�L6%�JI�7�o�VA�ݛ�v����Wy�m�g�3Z�Н��t8ݰ����� P��Kͥq����5�GՌ��L������anU{}��}�B�^	��,���[)�vw2���+��lX��@1�"m��t\��׏�
b2�?ܝװ�z��i&���p�4�n'v!���׈��e3�7�z�!��3���#� ��e(D����V�_�A-3H�e�0�2�x
"C�Q��s���õ�� �����[b2%�� �ī���Y�d&B����D��gw�����8�Z��C�)^�i����� �.�B7veF�-���~k�g�wP�e`�<��I�ܫ���Ala������L,nU.�2�f[�A�"xϽL��2�(����s�	�����C�ߗJ��o��V�Zc���Z�ăO����
�����B�ɀC2�p�2���I&����9m�G�����5i������N��A���ˡB�"յaa��[C�쑤Z������t1�:�ל	�je��Y�vV�>g� 5ИF
r�]_�����{��9��qb��%�=��i�w��~M��9̫�C�z9��� ���JA�d��e��ښE��0�܈�k!��i����`�� Y���ȖƵU��C5�u�P��[�Q�sc�>�f�f�!nf�T���MDmK���7��T¼�d��*pLe~�v�O�¡O3ڿ��a�������ox/f���]������)_���Z���ϐ�w�H�~A���;���+�3bTnAzq�/�W�\戧�H�b U�����\:��:��&'�ďWf�K�·
��r�����/".�c�4�L4��+�.e���eS�ݻ�i����C��bԹ(M%�PN`4�5CX�c�>ڠ��r��}^,gfcş4���kY͵͜��.�i��*}�})-d��;X����g���5�QG'C��	���O�~���~^N��OgΆ��q)w�	U$ؐ#c�GlԨ����؅����`v�b�1�EF�q�c5n�`K~VV�<�ωB�e����Q�~Y�	�Ạ3݆������X^ ��F�1dL��;�Zrf6�Wݬ��Aɞ����a�W\�&@�"���?�dOL,�\�س\�e����\��Z*҉����l�(nl� �	°sEV=o6u�jcƋ~�H��͙�8b�;�y�U4��lZhpU0ä�(���Z����z�Q_��Dx$	jIHe\:�qw'n���1�S��W�E)�sT)8�(�VU�Z#��'�ҧHJg��y+WH�i�-����=�?BF�$`(�|]�b���l�/U:�4��/u�>]ϓѨ(�x���iړ���}>t}��hn�G���xzI���_��Y4�T
��41-�N�
�}=��`�X�;��!�"�