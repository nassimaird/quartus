��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�˅������d�xp� �5��B�{�	e��Hk�Z�徒��{��\�83,�p�)V2V"'������'v�{��A��L�J��ʖsk�eRGAO<M��a.p�b��@�@a�;Dep�r�p	1��"32G º��*ڦ���ƫ�r`�c�}_1������	H?���}� ol4,n����������\p�kх���F�y��f�T%���^5�����8
�2j��pVq��zK۴N��@� 0 �	��ev����m���z_ws�=����#͑��]�Ţ���FC$����
�4o��3[�Y3�v��� r�'��̷�l���S���W�v����E���1��_���Ѵ~���;�ﺴ(ܢ]9�\h-m蹞����3���Q�ó�?�A����Ƶ�̟(|����g��~�Q��6�tg��}Q>�CW��k�9����ΨˡI6I���OS5No��k*�D��p�(ޚ8�5���6����I�0�~����ǏFA�2�;ҩ7^&�'UNg7���ZE(�����
J�E��B�:w���'���W���;/�R��y�p����r��Q���Ĺ�х��9�v|e��E��(h�,k�NNk��xL9ӌe�9:-cJ� ,��[��.����r�A����eA�v�)����8j1�A�ƨg���o��������Ƨ[cP��^��r�Qfm&�ؿ����I@��3Ml����Ɗd/��gčZM��H|,*-�r|��bo{��@C��P�eV�c����C�u�μ0�3�,������N�X�WBC-���2St6�8� �7Uƃ��rX�p����4�P��V 涱�P�n��)\��*՚�S
��V����RO�����d�׾�����P�䈾��*�A� 3�b�S�|�>|0�X���w�g�g=/�CmL�~q��4|S"�p�Ń�%Dd��E���5��@}�n4��`���/�z4�5@���Y��R���ѡeM�t~�ao�r]�4lQ�4��e�ެ�A[K�����>?���ʷ�ֹ�X0�v�n��d�v���� ��~�VYH��& ����+���r�C�}El���E=Lj��٧R��y��\�-v���\�!27|�HD��~����s�5�a�zh�����p�0-k$�6Ґ�����C^Q[)�_���4�1�饗�x�A�ϱ7S&h!��G�����zi	�;$�ov=nY�r����#�J�tL��|0��ۃ�H�����;�"1��}0�J�YclyFN�d�PŌ�K%���{dѴ����(΢�M�4�B���OJ��M[=L�#ϖW��45�	�e�K�k�y�zu���X�8�&G��׳�>�7�n1F��!o˽�5Z?�A�t��I�L.���B�yt�[.(�Q� ņ������ `�ӵ���G��!kn�@S�{X�Clr`l�H]�V���.5������_{=��`�~gY>�8�⾢o�\�A�������2't�eV��(Ӿ�x�[y�gbR�4e3ޙ��<�KA4����oȅ棛��路[Z��4�T�k�X �d��>Q���ڼ��ol��n6��,���ꜘ�⭐23���X�=��8Z��q�ܰ����� (��(�aH1~fb�b���W
�$���v}��KU�}Y��XR^19~o�qkx�T��5�eQ"�a5ǆ?,�A�x���Mۀ����#�0�����3�݅���1s���.p�d���|?�jz*��E܏ �r�j�Qȥ
�"���u��n��$w��5.,e��s(��\���KU�R�e���B���5�����侸��b.)�gL7�E�����^�s`�|����=��P�?T��Y��]�4J��^�Z~�j~����8�w_C�.�{w��~�^�0�	5���V&7�
[�-��x���i)���@��(d[�R٤�s����;�s�h{�((}��%���(��j'�0�/�[y%�/���.]���0�3��^ޗ0(5:��K��%O�Y/���U����nq�~r=\��d�Ü�N������{�{nܶ�Hw��� �����Z�������;�8���w��_�Rn@y���az�8W�"���W��0�%��3:*�1I7a�2Û,�dd�����'Ͼ���Z>ʁ�*Z.*R��dj�o](q�Lò���������<�"+��.��Dz8�I�ujl�|A��uF�J3/ ���k�&KH�u�Ta�+`�c��[x.]7}�k�{#�0�M�w�3x^� �ު�ݢ��������m}<��C�	�29���/��*�P��Ñ��5Bg�Y�XdO�׀J�����Ib5���Rk��K6Sդ�Scm� �ii�Ӵm�14�'�vE���|㘬o�Ց�3"� |n`NH���e�ʾ�H�$���weY��rʱ���Ͱ��������̫�+��ʓ�IY~^�uN��6�k
�ٻfhy
dI0`��mׅ�D�V��v�"��G=S�I�����),��0e+�}��{���9s�z�*�*>�D|�ft9v����N%�H^�~l��؄ݥEL�ޚ.�qvG8�p`�@Q&^����Eݴ���]~��	(*k����Ÿ������ya��̢�V���F�A���_���h�WP���(�_��o'�(Hn2�����E)m��[7 I9K���	���/�!1+?:x�G��_9yX�O����7��abM�O��l#��P|D}k<Hm����E�J�ӯS���X��c�Я��]!5�����L@2����(���7�7&�I��yR�h� ��8}	�S^�1�x�3��3��d_�LC'��;��n�8��MǾ��G�7у���WiJ"�Q1�γ��;����*�B�JU�WΈ!H��f���}?�ɻ�OE2>F�LtUx$��S ��n[ �u���Wz�����a������\6��$�Ȏ����<Zd����,���P��V���t��P3(�S_�N�7��r����3PE�����˺�9`��/$�&�I@��6�Q��Վ?&o�����z����9Β�M�.��4-��[f��\���&!���2�A�C�z��fJ��k�;߶_�����qG7�9�3pw��@aN��*B�i�,��Z6bՈ}����E"���57�k�`�1��4���'B\�s��Vwj��4"ʮm]j��*4�b��A���f5j�&�zZ{`i�:� ��u���?��Ƙ��7�����m�?��R��K�o5}PT���#vd�C�E�4~���A�vǜ��i���<lP�,g�nn9�;�t��LQ���;�39�(:4��Z��i��_���*f���������*mh��qZ�QV`ޯ��T/�;�E�/���W�]�ᓧ2��E��-ļ����'�kJ:�Y1[������1�sD��o��5��=؛�×	f��OK�
������X�$���6g!��_��]����cJ�Ԛ�^��UM��m����S���N��\���:?Y����c�� �Fk�P_�S�w�Q�SJ+���cR�SNVM6t�\��h:7��al�>*��[�q�pn�[�ٌ�D*f�&�3Ւ��~�:�!�
�`|~�6I����a�:���?���\��c�YC&u\����Y�t#�Nx,T`ee��!C��k�ꃆ)���<�q:�h.���%t���`�>�0!�Z�>Y�kT�_���_��u���-��ev�S*��PF��(w]6������l?f�q�#�']����?g���ф>�$􀖭�Zǰc��D"�P��a�=�A����-))��[R#�;�04H��8��Mc-��:�0F�l|v(p��k���uDI��A^�Ƒ�vj���K�~p{�-��]���K!�-�)Y�*���D��	�o��{��lq&�@����B���z�H�}�. E'�㴀X;���|�Iz(�"��l���CK��Ft]��v̂B�w�e���m�b4���0�᳣JS^�!K��rxV�I���������񺁫JU]]���o>i^���t���:���8A	��ؖM\�dE��g�%��}-[u�j�kn^����OE��=�#���_�@?��	�(I7� 0����],�gD�&a��o��	�<�qi�lo�3�#Zdy�?o��G�F8��)K��[,do��p�-k�wq�8	�:с<�A���?�]�9Y��C��lS|�x���i=;����Z
��JlbKѯƨ(;��/���v�E�moC/�P��w��O��
n���̓��[?���e.�!4��DNVp�7�Q�/�ڤ�ѱ��\t�đ,��ʖ����w��lj.g�Ǳ���	�ex������Ǆ�iS�wrYg��ߜ��ޒ�$q�b�1�ע���&^׆ˊ��6�5
�AD����!�M�m2r�B�$����Bn�e�OC�	T�-¦�d�5���ׄ���^��5�_
�j%�8^�xa����b�.,�-�r?�jj4ZL�+C���g(9��گ�xO���:-��x�k}*ME_�Hm�{����ۆ��G�����Ԫ�'oM֕��GX������[��(x5�J��Q���EC�M��E@����eJM�-R�oخKn��D�9rAX��P��l�µ@{J�n'{S��6��~��������=<Qq�[T���D<m�k���ρ��r`�Qp�\�M�#U/�Mxӵ�l�4{n�h6!�T��E�b��uG u��=u��j}o�-yj�U�~� � U?�������k��5� �ۢ/��3�%u�o�!�j��l�I@�~&N�?�h�C�N`�ߜ8���z�S0���)���ц+ ������R�����@�]�jA�y��$��ę�7�5<%7��}l9�A��gzyZv"7U�Z^�Ë�޺5����`��4kA�/�>����9�*�1�
5���i�"f�꥜��I�J����B;�Wt���!�赻r��U*�͂�+ݵ��2�
n*{�~t]o�+�D���V���ͦL�J�X��b�����^�i��H�Zع)ޫA�3�����R��X��,m4,�?��r���8b߇�n�ݷL�t���T5� �.ۿ��y�-�CPg�d��`ht���cBi�����0v3Ҵ����2_oB�4�؞n��J5���g��2����r���
bG`���ص�F�����h���UҠ�u��w4�9a���ŮD�#��` ��K�e���1�U��dH����e������u}շc�9L�oΐ��5����U�7���*.�N��PF?6�7�H����bb�>�)i�s�u�j9f��	+`,�U͝l�-�KPkz(�ċ���(O�쥧��%'[h��K�+��/�64j��]��i���נ��V��B�i��������T�����(b�Y�-]�O(���� ��%��-��Ռt']E�P\G�i�0����� V�歫o�<��M �T�F&���(��	:kn*_aW���|zm�֙��)�I�}�M���UI��$�ZV\$�Z^+��]Ty��6���|���.2T��	OȂ(�%
G���vj@�#�©#L�ס�݌E!gD�� �/���	��;e�c�G��^C@���J�Rz��(P=(s�!�Z��4���?ߩ����ED��%�������š��4i���b���OQ�P"H'���-y��2	��ʗ�%�q(1��&�>1�iL~d���ͶӞa/�pm�ܯ������U'�]�[`ws�t�$���7]�8�{I�̥D�4�[��|Z+%vt ��(؏2���cڻٻ�ϮRM!ky�s�G*�̀c����RVwsR���ʽ�����9��鬱�++�.��N���xd	� NBB��ђL�J��3�{闪A,.���˓�0sv��E֜��Q;�b��ؚĕ�Ӿ�-��˘�R��o�p3o�rf2:��o�{��g,D��*X�`7AQ�_J7���n`%�`�.��0����_(�5�ޔL"( UCzD>΂�}~b[ںJB�p骑�ۻ�D��*�����,�q����h�x�`�����l���`%�w�ߐ�3�������:�^���dmw�_����O��1�8#� 0�C�KQ��v(���*Mm4���q�&��"7|�+���3�V�@��û�Z��ݮ� �m���~�a���yX��i�|����VXo��bin���JL���Yz���x���u�C�|��֚���J�~ ��ֶ%78��Zb�ǜ�8ͳ�	t��03To��` ��Y(��)6E;d0�}fr��y�G+�F�_닉�,t�mRS��	�� }
�,`�wI+�y�UL>��Q�0��scE
�H�
V���O�`�w�U�˙��)2C��"��s"�q�P��&������vLl��*��e�h=�c�����E��r��� ��8��xEQ��Hz����at�#������{d9@�d��>�֢TA�oph�ωj�<U3 ��9���-a�B�!�f(�(
Z���6#g@\\�f�:�}�������������~Ƭ$S���G?)ޥu���aQ
Y!�qi���\�+�Ȁ)4ԑZ����*�ӹ�ydSsT����K����WE�%x�䜵^m��6zz�d�K)�)�V�z]�k[r�	���k�^RE�ɾ���=PT;�j���w>߮	�����z��l��q!^w^/�L�ϵU.���)e7� \5���T���3o7��l�B���pa��gl?�8�f�k-��|��=���Ꮊ�#�_ .Ej#�=Y�t{��& �ѷإ�kk	1[�*MD��c}Wj,x;�R|v���q���;���a��U��I7����$U<��FF��9ö�z�zW�`Í�&i2̬��.iկ3��H(��3��Ձ<�gpv�Z͇��z)v�L�'i��y��x��9��~�U��g�8����@9̎]�<ң+�U\y���#��
U�2}D�*ܴ-d2�"Ew2E��R;r}a��zt��H����k��8�#rP��KtNo�*�����e3�Yeʋ�=�D����0���%%؞�	S/~��Ю�`�0+䰌�4�V'u�kX��9�y�v�30��s�Y�Z���\#�v<�+~�{��ܛ�y������0H��Fn�w`H�_ �a���M�7�0�aw�[/ϰ�xZ�y!��1v�����kNJ��;�#9���1e���%v@42�����oc#=�@��ވ��� b}=�m/�ʽ���7C�ZN���(EQPߦZ
m�v�Q��z��򝀉��lw�v}��*8���)�D��@{�9J�.�۬��Lʺ�]?�	f�#j컯�sFYՓ�cH����`�P"x�ɿ����w�v�u0���3O�'@#�ˡ��贤����*f�кx��0�c��"�ŭ �Eo�N��Ds�m��b�����^�":2D~�ߩҙ���Y{ig"��"�^�b]-�װ��S���*D��ʣ]A�6� ��L*i���<5>���q����8�:;�5g�����h<g�ę�tϝ�frQ����cʭ�op��S�F�S}�>��S�FrX&����m�z��Ib�i�4>��C�l��觧>s$C��2��L�H�_����z8q*t6`4���W:%r�^[�;g����aj�ۃC2t�6�қ����X���� �b.9��\�Njb��rq��p���S��ѧk:�g%������I�F�ͥ1v��z�%t�}�3R䟬�:`�Av&=���dv��]C͹Y2� C鞪C�����*$R���D��1���NECe�7�^ב���7���_K�$�w��FX|���ED�%�"G81FNla�8I��'�40�_���K�=W���R�#�v]T�1CMo��g�	X�s�xcZV�����S�01|���O�F�;�Q6���C_��V�vW�D)��&l7s;˸����<c@3<�yZ�`ڵA��ڷaN/��k��'���UMP���j?�:�)���H#x�GX����k�T-�i��
i�o}	���ϡ���l_/�Gx���\����&k�Ն�qu��>M�2.]�0ը����d>��Pƃ�@\i�]�Id۶���yZ�:׸z��ax��������9V5]��!W\�v�u��cP �m�+��æ��r�i���	;e��A����~��z��ca�1�|�v�"3�	�y��k���c��\v���R�U�z�S�Kz��n!������#��f���`^��
OMP�b�`�4M�t^V��/�@�y�Jfo���ͣ��K۹�4|d撫��Y�Jj	O�
���K��Ʈ���Y�{�J���e�Ct�
�}.'`&�uސl��&�$Wn$���|���Z-�o��)^���NcxsBa���=����GtڲKgԂ�:����gX���N�����!x]�Z���#���ƛ>`�)?���/o��t8=COs����d$re�h���u֖�r�!,�A$g�Nc��xE.���E��.�S�V�*���U�Q�{�0��Pz�=�?т��Zң�e�Ǆ�Q�|��M�?���A	.D=,�.��<p��в�j�Cۦz�S�Y6KH�v�ړ4���dfV�Q�.�zG���pH�wY�	 `�!+�.���U�����D��{E ��n������P0��h|f�op�2�[�O7_e��]M�B)z"�'A��DW2y0Yj�=(����_��.Pɗ�^���g�:�9�l���Ӣݵڹ~Q 5��I;�!>$�tF�'�c�籧jH1��H��U��o��T&P/����"c�'��38֐�s�����Lq�uֿ=Aa���>k6W2
�/6�*�"�>�Z�ɦ�p-[|��VT@����q�p��rJ��Yva���e���Z�Y�ى�R&�l��M1�a�1f������~eu�"@��^�����/\��ԝ�E��t���m����e1�F?�g�A��"��^?�|͆��IKJ*�C  ���9ԩ0R�`w"U��b�e?]�;U"�T�;�q*5T�&ϞEܥ�eջ:�(���Q5�)�T[0��cw�X�tȲ�@� m�Lr�����/~������"���Sd��4�?p�	V�h�R�o:��<Y���
�>|y�+Yo����/*��f"o�f'���pde/qs�-�3`~ظ�7�P�+�Z��\YL.(0'�7�V$UR����W�g�e�w�����M�8���X��/x�)"B�>�U��׫-�e��vu��eV,l���"��`ԝk��N$����v��&k_lԝ�����~��sl�i�Y랐� �SWf�=!�B	_��.�F�<��.�OFa�B��;�Q�F��9D[���������
��T��9�����]�z?V���]�V���ZG-�w��]�9{��t
�NW���S{e�.,��I�l��_��q�����3�xpc���6XsF}Z�n�o���%�j/"#.�l�Ny�}p6��c��h��?��gM���e��t;k������2�Wʕ�)Z�Lԩ���:H�,"<�@��l�\5�nܗ�I�0@���`��^ fM��6�j�u��xĴ�W����v��CW�����7}Ǣ��|��O��6�/� ����
i�&�x7L��S(w�	�Z/�ȹ��v��H��<�����VU�[����Y$&_/���wp��1_fU�_����YoZ�ȣN}�>LyO�@��8��P\J���;?z��s{jj�iB�x�JM�N��<���*�¦�Eㅺ��f#<t$��wb��k�4�撚HD�)���k�Yh��t¦�*m��t�D�s�aa>D���8t�[�|W���[ߌ\���a¯�/VXL�9�8�`R��f;�y��}��~Ѷ2K�XEN�2�r����o��C�C��nk?#������W�qƙ'��r<V���8̓����3������E�f���$�^�N~���Ԝ��.�.��w>a��?#Rm���k�����Za��0��6&�+�sZ>w�&�Cb7`�'1��ݑ]�,.p+�)#��*����D��	wY��K��~ A�k/��e�+o��pznU#���>d,�7��z���/[V)H�#_Xoڦ J�g-�=<��_ц�
K}cL{K����L_#��{nL� )�d��;���V�\�z|zl@*�@���/��Z��	�L[?�ƹG����ZӅŬ����c�_�g"�*���g��rW�$�t`���c��j��f	�Leoc�����"�H����V0�4�XS\�<sMda�&c�j��M+ދ���=��6x��z�º���lG�U[��S���q�crɫx6��)$�^HT���{W*q��L5<	7�=��@:���}ڠM��'&ov�oFv�����R\ÿ_�Py����M����*O$�U���o?0=�N]Aa����]�y��p�Ho؟�([�IS�XX(�5�m�w�R'��.P?u�4;z32E�����b�˲�5i���#`���趲ܪ�ׅ��d�_��-]�_�d���X`�6�#}wyu�,G����� ;�a��b>�=��hrV���Ix�O����̊�<���&mM�2�B���+_"�ڤ�_h;T z��h����&�A�	 Q:�`�Bq �H� ������Ev$�1��M���=��v��2�%ˌ�2�Ƴ��G)�}�G�h��x}���0ڐ1h Zf�.�Z&��b�vD����s�3p/��{��
�<rVgyl�m��(�N��fr$D���wc7^L'�\���"��,�Ip�f�>��7�<vpRX��yiNu��ܻ9I[DL��vL٫���}���^��m�[�X¶S>Ct�Ȥ�o*x�"��r**Nc�����
�o~ڦ��7�
0G�N�~��G5H!�s����p!}[z��菡�xIE#������K�sH���ZD1�$�W���x�=y�&?pz�({�D��Dː�v7��}��v�r3ӛ�֓����9�tx����Y���T\�A���B�Q�����r��L�cգ?Ҳe$uqv�>���8�!��Xj���g�k߶Wb��A����Qm+��#X���\�F�n-)POB'��^r'*�'H��W=>P�5:�E;�$�b�-��ʯrJOhz-b�nK���5����=ۑ�o��^[�N�����U�yc�,ƾ?N�^W�����!Yد�YM��M��u��6�����޸0���o��3�=�	�ۇɷ�����Ѣ
g��nX��u.�Z��+���Q���:���:T���c
���e��#ԩX~�T���9G<#����������}�3��P��������ԭ��l��D��Uo�~r?jd�wr��*%��e���<�6��c<&��[��ibf�q��묚~��b~���u ���-��D�Q������R �7���֐��]F��]�����KE����,�}�u�V�v�UFt�SǒQ�qZe�arD����zCXL���Ux��G���W��QP�f8�~	��+��RY�N���r�v=������4'u�����b�S�U��GzB�^�)<,�����d�,#�Gc%�!�T4�b�+�Kܓݑ׸��9Q�ԟ
Z{|������kn��?�b�C�:���( �;:���S-��w�)`��{�jq�Of0U��E��jP���<�aCA���wV����-�-N���O7%��C��ض7��9L�ԫq�R�k\D�X{�#��6��kꡝU��L\�u[$an��4�Z�� �����5��w �m`����Y���|�wy��A����Ȳ��.��|\j��vB�/�%���;e��n���Y��>/%���۽ЂM�c1�����i��O�!�'M���้ϸ��=�q9�r=�t@C��ԬIa��4%3+�WB� 7��|o@�T���,�w�2���V��:Bೢ"�d��X#��=0�f�/�4h�zCW� ^��uf�띉f��.8���R!�9��v�RYg���HU�Ng��YVr^:����&�"$$�tQ�,mI��1Ű�=N�&������y��g��#��N��D�m���{,t�Hq� ��V<X�&�c8�[�zwg�<zyu�i�4:|��7:�e�5�c��L(O��5�}����!���wM.T�[!��Gj�7b�I�I���T�d5�l�*�g��/�$�@E^ᙂ]�b��Lq�Z8��;���b�����������8�dA��`���A.G��o���-�<�M^�vd2��^f�ѼȂ�$���<���6��:�b�����������=��_�qOʾ��~
@��	4�H[$��ȵ�$i4<7�V�
�/ѵ��澃�1���6��Ǳi�
>&���B����U(,���ח}�bNNn���S��c�����gڃSŊ�����-�ܒ^���6�B�P!�1R� �¤͍X�����]���h��XY	�Y��Vz��\dp��! Z�t�K����c��8�����+�U|���v�/P�j�O��z׫CG����z�W0�:����9T�xФ�/y�)t�o�xG}ֿDDAv�z6Z������τi���</��r�_u�npB�/r��&]�ڟBo��O��T��]?�
9��Ö�<�?�ImQz8W�ΖF�A�f�53aݹ�M�����d�kZ�dal�����Xa�H�T�����<1A��B>�d&�����C��(L?ar�Z���ݣ��*���sF�q�wdvZ]������[�n���h��q*㟀q޲���4��$��s�^,��3���k�4�/Mr���M+��>��EC��~&(�mC���!���g����{�t�2�XQ^U"������0JS6�x��<�Z�׸v_�2U�q���o�=�������#�RL��Oa��w���fj��q�9]� ��i�SSXP[v��}(i,d��y��
GS�K�'���H�����v3�,�Z85��7:2����Y��(]�F�����H��ƹ�gw���������:�@ˈ��?C���\�������;���ĺC9��b}KL�Ǎ/�����hI���V���(f�s}�N�|�I|�c0��M������V1�uT|�#��D��ㄚ��C8s�m���:��{k���C�b�幗���	ג������C�I�ϲ��c���x"O���Ԡ85��E�6�K\�1��W¯��.�=�d��������[FR��$t�	
�� ��n�A
1��3��̘ŝ�8�.���Y�ޭ�k��b˨�ig����&�E�t)0xrՕ�+tD��y@�/��Me�s8W���+��w��Ѷ���ӻ���I�厌@s*RN�CS���!kO�M��T�E���ó|����;x�����uW�à�Ꭵ+�Β�!k�G�FĲ~���W��=�4�Mܓc|ߤ����{�����;�Ʃ����i{C�����\:��S�M/�{Jp3��y�"��hP��b�qQ���Yh�g��;G�K�x������� �R0�I��TG�8���e>+nou��yYf�i�Ti_�'�'2;٣SM��a�\ic�{�4rd|���dX���!��*ξ���A޻��=/S'G�O�1�S[o�Tʲa�M�v�)~�ͳv4��ۛ�1h;aڶj5�Ss�+��>�*�v+ш������-��W��Uv��s���3/<޷�2'�q�gy
�Nݗ�xj���
��B���,�;�m���A���7�J�2׫��=r���A��}q���6��&N;�(�
�B(���z����s��������E"�K�������e�O���GT��,n�\j��b.ƆX�);�*ۃZek�w��Y��`OKU;W߄ �E�+���~[�#��Ȣ0���k4���;v����c	��h�u9r�\�	�!�XU�W�_Xܮ��4cR��oL��<���ɹEqqa_�Sc�skQH�ҟ�����ڣIm�%�V�@V=�%�_'��&�.�2�
��PT���P����0	���cȈoϪ�zG�絕\>������I���Y�R3��`�wj����O��.ۂ��'+%h��S��a��/L1*5L��S��:5�պ��v�({�V���[&��aC��N��l�3�tIQz�LF��Z���}%�p|9R�;gź����dR\�k�����-<ڎ������n �U���W c?�W]^�߯1_�^fɍ������pJgby}�w�\�������,rq���{>r��0�;��vOr�%q��Xp�4f�������Ǐ��sJ�^R���Lz �o�~�o���R�=�}I׷j���_�5��;���ö�8�2���t["�	 �0<�Cr5#�c�qNrK��r�\,����n�=���Ѩ�֍�	␦_o"%�/���cC�bY������g�1���W6�*N�@g��A��C-�V�Cmv���>�]��z+��.�]�C�wV�
,��Ɖ˛�	���L��Gd#�m��r{K=jƬ�d�}��#��W��X���E���b'i[s�\��
���K��E$��kz�o�ӳ�"8������Ug�W+���Jsrh�V��	y6C��Hzb��h9Jd_�7�b|�j� �j� �-����m�{�Y���8�V��qZZ�y�iw����)���N�b*��U��?�׏�G�`������vSg�e�t��v��Y����j�Nz���R�.A���V<r�'�tŷ���O�X�Mg����V"���_�%9���[`��������֫>��huNl�_Ɏ+T��	�
[�I����)�Jm_���oxȡs��� S��C=���̥k%<��W=�F����dCi2����IAT"n��g[`y�����`Yp���rŘh�THY�<v��7t�3���Q�Bꨚ��*�P����.a��Z߄��h�]�&	X�� �z7�[�6�����HF+�!CLLX��Sz��f���GX���q��`�U��:�����܏Eδ��	���;;��W�}��rn�Z��Fq�_ �`�H^`QM���]��T|b��sO)��H$3��D�N��F#f����3ȳ�YW�<����ʏ6QǄ7n�ArȍQ�<i��K�K�EV�?�fw�]I���Aj�;#EEO
^�	�쩬��D��$OрV�tGƲ���nV�ӌ�$����w���H#AtQ��P�u:��i���m�Hddqh�q�}�	u7-��V��\��֣��} \�mu�Z�D@#��N��&�
��Y���f���"�L��L"���D����%T"�&dM���<����0lv\%g3��A���<��t:
�.Hoc��!�ZZI��j�;=nvКJ?^��
 ��	�g_6�l�ӎ@ʒ���^L_Aw%�f��8���KnC�������W�5� 3 #�r�"s�춣i�w�I�No�vh�c;#�RL�2w����3���Ŀx���ˆAV�y_����D��(���k�4�R�ȇN�Pb���>�B�A�H��twL��qZ�놝
"ޢ`Q#��i"�z��FX�]�?�O�\�B��sv�̣]�ASǏ��˹�� f����g�fVu�������Մ�2�ے<N�(&\�? �i@�e[g�iG�Z�Z$d,@"� �pǌ@�p�D̐���Rɚ1	�sD�ג��M_!%�#5�C};*M�S5� &&G@T�ycӠ)�S���%���j{@�ү���H�W����ry�m`Y������h
�x�n��i�J֘�j1Jc���{&r)�𩤂�YZYaƒt��kӪ�����F9t�6n5�3�5k�����[m�ﺼ	I�58qЕ��{�Nj������m�:' �Zp?fY8�����$@�>���-�nX�6h��ԭH�?͙d��fm�����5�����'�΢�@ǝ�s��q&
����txpK2Y�u�s]h�0l���Ϸ>>���ԱT��Si������db��S������L%r"��IgWu�|���;h��	K��������s��?���xׄ�~kr����)�]`���4`HQ�U�'+q�
�+.\�2K�ҭCݧ^g�21T;R�s���u(�Mp�WKoXD�kf�W��M��1�_F8�FS.,i)$xL�
B��x*lB�:r]�_�\�.�L Ž�`�sC��j<���2�l��ߝ�W�Ή�9�Oߦ��W��1�sՋ?�Ν7��	I�p���uNR,�$��[�¹؁��&�:ٶ��ؙ֟�՘QG`�(��s�X�ёC�׋ȋ�j\��!.�S�O�I���*_,r�1�k�a�s��!�v�ik�͸�v��q��_��Pj���z����~�R�?)7���B�^8wpì6Z�X��o�o���(�t�1��tb�l�_ӿ�i�Zr)7� 85w>^/Ĭ�f����9���n}��9�c�s��SK����3d��Sv����p�G�wa�W(�te!�֎Y�X-{���W�Q���5!=��]D[��8����J�+7������V@��YQ$��������뤏[�ʄ��5n�I&g��eȄ.<��­pSfH�(z��`���0D�e\M9�5k�u6�l��<��w5�߸�"�ͨ��a%�|E�t!\��Q����T��{7�7���F�'n��5�?�~��YB뵇�2o=Ͼ=���_���m=$�Wٷk��V!d��C�>�YPm��l�ƛK�U��L-�CQE�Ƥ�<�G{���v�g�W��0؝�l>�+�T�?=�1k&0�B�ȴ�Ѕ@�1�8��z.�5����!�#x��4��ב��jn�xR�2���u$8�Ѝ!9��f��*O��w�	x9���a�����Lud���,�am�����;�����T�	��;�!�=��&	V�� e���:|�\Q�w|�<��y��7f&q���_���Ny�
�L��C�H��6�m0ć3gH���W��j�����_��v����լK�$� RK�X���㷴(�Ƚ��/�����sǷ(Ot%��u�y��z���#��B��KBHT�P��i��l��PE����%7�j#1����d55A!����qQ�S��H3l̷=WQ���;�s �(p�	<R0i���"�����a�]	܄�G 񝄿M��؟��N׋����t��=}CP`�j��"b0I��6��f�RV���v#K���H�8Z-�]�e
�C�;&�k����!
��y'P�}9rL&_�F��M�>V�F�!�e ������|��9�<�B�G�Rz9q Q���xI1H�ϐk�tagyTG�k�*�YD�M<_��=66H��� �)�n�a�^)�J�ܮ��Il]�N�_��?6L�أesGH��Y9_��Y��zW�à��Լ_N7D����d��H��
���y /,9�1��3I�Q��_/�:�Z���~&���V&?�m�H~R�K?�&Ϫ!u���ꓯ�j���kV����D,���[��M���@�2�?��O����O.X�a��9P�~�Mml(��KQ��Ӂ}�	h��K�5��ĳroB�w�6��A��B��ht�:�0�I�Q��8��LU��UG�t��|��[��(!_Sc/<�k����hXc�����U��L7�~�E�Ag�~S�pv�ѻ�c��-E���"U�.�e>!�6Wy]ힳG�`����b�W�!J2VME3Q��-��x�a�NH�j,j�ct5XU���M���z����(����[Y��<R�#���z9����h�3"D�[�C���ś`���9&��w�A����d�
�e��8�!�*%�!�f�~�"���G<犌7'b��/�a��^�ਿ��� �	�S�`���S���Z�j7�R�
�!|�/��}�������{�f�����m�X�ɕ���^����1p?U3�IcQ�,k��`������8�w�c��X#O�Us�Q��v���\�_�u3|-rʚ0�"�>\�������9 ���S&����>Cs}|iT��_�~$�A�T얯��BD�$��@���f�{<!��Sq>��jlQ �`͗�T}:z�	#��~�|�Dic$���IZ���*�MW��������`�z�<;�nf�
ˤ*�����-6������lZx&���iX� ġӞ�evL�[��@f&␭3��0#�*��y/+��M�E���(��*\��x��P��R�	�|<�P"�1���m��`Rڏ�k"i�l��ʙo�[sj�3׺14��C�\3,�u�b�U��j�}I��;h����N�ôT�d;����y�,�W��t����w݈dD�.o�?��^W�D]U�o�p�U�?�c�����W��
,)��K옲�7@	��������*�u�uz0��2D�t7�'/��L�~o_}_�ND��A���|��c���*���}�7@�/��C[�8*vO.)!X�C�k���5���X�WJܻǃ�(� ���C�R��й�a����?�?tX�#Wp�R��\`8�9��h�^Q6�ɊM�Ω��UU��݋r��� G
�������J�Z�E ���J~G3f��7WU\�ɨ�gC�9��αFHs{K�d.������\��Xp�����@xb���2�t��ZBLf �����M����=bz��V��6�On��aT��{��)3���bj����H�e��+��d pՃ��)���8v����K]����Z�W!���%�啈{KIj	�{X��8�$sE�F���p�)�Ɉِ\���W;������UAn��^���J+�	�Q�y#�e�],U�UP��-�����`��U����;��<��W��Z���и[5�j����ky�fúP]��K��
����.ᅽH�	�,��_P���}��뛕?Pu0$�7�+����k|����KN�ZS@���v�3&*���-��]���,.Z�w6Ki�X�	�;
�~�
i�u���q"�����N��~F�k�_��(]�9<��J��F��b��E��� �^yZ��`?0�,��˴>)Pc���##�w\�ڿ7���n!���M=�#pm˸���Z�E��{U�Iz'5NU���V|�j��zņ�%b��\���9�<��[���#jRi���*U������i�J4ga���sb��J��PB[<5g4���<R�)������u��\�=ƖI$�i�ƨ�x��P7��m�S͓�V`���k�;��Ķ�S�G z�01M��4�z�UXg�0��S���j�nF��T�������N05m��D�%��x�HJ?����Z��mr���YF���o=���֨)}��|&w�íN��QPٺA_ܧ�3'�2�쏇E�B��QXbǬu�y�}.,�s$��7��>}����xHR�͟J6��O|#��jb�ӑRb���-3>>��߆X1ݰ!w�����O@��hJ��ج���@���;�~��.O�`�xV��u��[#<4�mp����"�J�}�	)N���,@��kN=�P��-um�ƱA�i/��Gj.st�i��S���KV�6���rgk��} L0�/�78�EqV���R�krhL��1l��Y���^��`��X;g�����l��p�.SR�������<y�[�D�oDQ3Y���q���8ֳԣ��b 8� o
\`*m�
$a;,�h*���I��}KF�Z��|2/�V+�d�K���y���a8g^����٘�N��X,-;���v ��H���[�cU��ZEJ��dv!��x-}wj�*H��������񫠊>�.��5���PF������	V)�5��u��0i�����%j}�)u��	m��R>��@nCnn{��l�,ň�	��)c����l� 4���!��������rr�Y��-��aTR&^�(��d|E蟉����.��9��E?�B`���]B��2��(�\}��(��*���^m���g֡Ƈ�t]��s�r�j�Q����_�H���& J��ɿ��x��d��� ��Xf��/>��9L���\�ПB0�ǙO̓ut��/�p��kSZ��C&G�4Q.%يsl���H�̈�D��Oyh�?9{W�E��?c�C�Qe���Od��b��+E��ShJ��f���o#����c�����Ɉ���Uf@��o��2ܸݸ�PlHps?(H�ݪҺ��H&�Τg���y�Д�	�F�~*��U�N�d3�$�%K[�b�0}��@� #]μ� @Ba�+P���a�n]�&Cd��!!45d+�T��-��?{ղ�`<Q�;�1<�I�B��c>��>I1OM��WV���Ap�s��4P���8f�M����I�[���yN�R����?�[K���FJ���
���;����A��>�1s�u�˟:4�}iL��rcP�m�'X�%"Lj/��@�a�5�A��� vc^!@�v�5F�y��/�H%�&�ٍ�6j@?{�TY���U�휑/�3�=��B������EW���@�T�v�3�3�����ժ񾞵������Ju1r\W��9��t�a5�H��>���t^�)!�C��P8�[Xj����I)������b�����H(E�%�%d�h���G�k;�A��֎��;k��㪍�E�����l�1Vp�5�5�Oދ���bR��q�Z�aH��e�q��r~���i��ɬ�R��}S�H�8V�(�8��';V�c��̤��9�dB��ed�4����?q�+�1���_xA�+���$4[��~����e��*��_R<�5a�#�1)����i �y2�Q��gD6[+�-�A!55�~�l�a]�P���, ���͟ࡪ���Y|;�X7��ӝ�%�q�M�ʜ��=��_�5m?�
vr���ϣrTg��v�7��Z� �W�ô>�T+hO��ځL��3숟�m�mh��Lݐtz��V������ƌuKr_�ӽ]��F�=����)��3T܇�c���Ј�lr����	���D�Q��k�Ϟ_%}��Ri�zFSъS^�?Ů2�;����!
kr�8+����`*�6d�T�LV"K�����*�7�� �����Ŀ�q�����j7P��h�M�A7oV�d��C��f�qX�~[�d$mv��-R�p��E�����>>`��}a�� �,|�����)އA?��u���S;+&!}�8 ��F����d�Ɣ~:xު�����{�Y��1��r獎#kR<���p�tk��k�%��u�Uaty���_�˒��X5.�b��|��R���������F��������k�@>���z��(U���v.��)�I3�xL;u�y���\V����3ϣ���p\!7P�%<�5g(o�BP!�c��h鎠�DVW�����A�B���l��<��C��7����V�a�Ca�!�5#r��r.�W��_D��xSӇAP��7�S����)��Mh��*����q�"�Y/V����g��v�ߢk�R���E�����7;*؅��u��'�Ly�վ�z�'�$k��Oo琤l��]������dUF�;�x��šp��'�g��IMfMg� WL�ݜ�����=��'��s�Ȼ�7�}�i��%�Nn��L��s���^n��*V�͆9�i;�p��C�{'�X�'�q�$��[L�l�!E�]f����|aݢ�l	Ʉ���gJ���fV.��ic�?���T�]��XY� �u#�g2�
AKg0�De�W:��0m�)�a��fJ�Е��c��{��<�h������*�p�L�\��i���}�ރF=�������VU��Y�^u,���7d���ȜR��)5��Q�x��K�R
{I?)2�g����[^'��6_c�g4��7]A���Rg��k�[U-/�T��FZ"\+��5���*S�c5H�-=������o�[��u���P��+NÀ��qc~��^�O�%k4� L�ш��SD!O�+���}��j6�-��.�E�}d�i�4�L$�S0R��9SN����)i�	Mb �=;�"����!���J����L����ً�6)1Yf�;D�>u_�B��g�째� �_C:�^okhH��0q���T� ������gV�W��زXJ�o7��࿞���p+��z��n!r��>>rʌ��L[Vw�\E�?8zR�mD8	��K}�(�]-�`2���Z)�5�5wT����?��C�AJ��:�9Mo(���]	)D^��o, *bg���:��vIt���0^1���g�'�gC�>�J��J��u)$|�<���\�ap6I�W�>�B�Ϲ�XN�K,.��9��9���s�.`�:K�Vp�Ӗ�7�1�&3���w�;��I㡗�<c�`g���p�T*�$�o�$���1��*�aL5|�>w�|���6�.~H���:n���/, �C�[u(v�0��D��s%���i�%z	��ypwo���x��הּm�b��u��n�JN�K�"������E�|L���Z6y2p1�5�3���Ɍdt�����QHw��ۼ�fc�S��=���Da�N�����7�؍�旡�@�Ļ_��t;����Q���� |\�po]��ّ禧P���r���C0nR�l�f�ĚԠ*,�Bh�@w`u�R�C'�0��L�<�XYߜ)~��T�G�9��o�P3jl�+0��A��Ї��@{g���X�@��9�o��z�V�j	�H����ݲQ\�A���)����M��8�bM��nс=B�����M��{
"=�����Ք4�	�i��t	;� �Lhbύ��cu��ӑ���P���kg�o::����X 6�eCF���*�o�`Pn0����� s�B�{=�	�ʣ����	��!9Cϡvн7�j�C݆�GcbC�v� ޶�Pc�l��m2B,1ҹ�S"��G�q�7�Cc_�Y�B���u�`�j~�̴�:TAi9A�Yq�#|'�� �a�j���7��}��}�e)6�.�Ik@[f�U޽�l�϶�Q������2�>f"]^E�,�'�.L3��t�%G^!:���٧��Q�2�u�̷P�Y���q��ru�
�4���Y#j[c���� N�?޻�w1~��D�}�:���8���)��\u�_�����@w�zJ]��H#���ޯɳ�z�ڭ{5�*A�An}�s��������O`7~xBWmO���'�.�T��޳�2�~�\�{_����/��P�L��z6���|D0��	�6}f4cI�5��{��RJ��������;Y�-3;�g�KG1��	��e�o��q9�hz-�*��u�SG�v��q0��c�#��{]xa@��F��k7:@l���_��d����q�~�]c�45�-��,��ݣ����B�+Ћe"��f�O-��3��4���ډ�����"xP ȶ�Uks�7	�61J@�i�����'�f{t%�q;WY	�� �'��ߖ�����,z����p�"�M�e=##O�� �E�ԑ ��8`�'�����p���M�N�l��,T
�о�W�5���?+���ʫ�.�W�e����n~�ޡG+�\f�j�I�4W���w�� ������WFʸo'���J�k�?�}g�2;��h,��"k\~��)�g"���ͷ_x	U#�4)
�G��c>a`s�ys���wp�)A#���T��l��3ԬDĝ�8�LzD�+�mSc'K���6���z���;�����+V���|]g?�f�����S�\��x_^c�
~��K����Ʌ��N�3Z�J)�ψ��K��z��)qB��\ ����{pЈ�Ӎ�߳�"����-��+O�J �g	5Q���}�Q�io���$w�k0�ړ�(p���Nom Y0���3 ��1�&�����h��>��mSO�fS�t2,tÕ��H���e��>'
���'��W]��C�o
�a�	�Ùl��ͩ�6�6��̕������6Pf*iYs̜��I}�@B���)ܟ֕��٠~˛w$��"��g�4y�5�݂���G�[v���Q'F���F*N>l���Qf����W%�_6qI�md_f���GE���)�yk\A�@b�{��}ЋWZdݻ�����	���ɯ�����+��ȝ]��)��1��'�Ն���5���0��BS��7I�6l�{�c~F͕��2wϒE�t��mYЕ�����w��%$��yBMFwTB6�yس������
�v?=��'�T@#nE��U��	�|:Y9�"o�n�a7��Z�
�F�"�`��ts�`~����)ԯA��:���
���	����o�
lMt��b#D}(��
*]R���������/�i��A�<�(�10]'��ݩ��͛��`��-c�g����q���VHi�B���l�i>��ό4�ӊ&��8ɚjU�r��PA�4G��R��\M�
�$3�sx��%����!�� �r����M�^|T�I��c�V�L~���m'�
�
,8w�9����P���k*�控�c�+�󍵶2 ��<䍿40��$e��s��5�km9���3�XUG!8y�bѷ��_����^��W-����/����R�f��O�G[Oݵ�F��E�n�)�o�}U�%Q�L+���-�}"����[o�T�e�{G��D�l氹ĩ���� ��O�>Q�c�O8Z*<a'V��2?dLo�Nͺ�&g%���S��|㊼���8�1)��(0���7$]G#��v#{�Ʈ���
E����*j�;ƽ_�^�~��S��#dS�/�) �\�_Y�z��������¨[�1t�nkفn;���q::�����w�
��\6�cwT�n�=0���8�&	!
o��¾Q��3�//�P[?����9�t�n\,��M�h����LO�:��,R�?��"eqF����%�XZG�(]Ӽ���Y�R}�2��+��t�翭�ŵs���)6,p�/�O�l�|�������$�!N�ut��A#��S`���\��������l`�(6G���$5�Zl��[ʅ>zQZO����X�K��1��U������� r��/[ą���𲣸x؊x҄�ԯ:�5��Y�t���Ө��n���B�K]�����M�vΒ��
�l8^�$-4A'��ģ�mF(�@;qoQ�)�`��pah�K-A�9*GeN uy<Z��"�d7���y����ў�Wik/?
'��Z��`ʡ��5F^~�}3K�iM@c&�$V���$����fH�q'O7�.�nޗS��>-V�2�CN[ߘ��w�,� 0����'���P���F��3��~�05}e�t2�K�Hu\�f�8
KSn�����E���g� D�<u�E<�MO�bQ��P9w�U�#�h��^��8@�䏆z�D��)��uSlNջ�]��rYi��8�Q�����V�Ӈཙv��U���y�5�ttȖ�J���+L��b�L�`��N�r�E���I�UjѨ�!B 1~
��N�������c)i�Vv�0��_>��(����ϩ���N�6�b�L���{@{q8k��wq;I�����J	�B{J|'�2�hK���m�د�kc���އ�*�p�Ҽ��:��N��<J��=޳�{-�����KY)�J�54��y��dR�Z������#[0�ϓ ��F73�z�*�]j屷9�3�bi�	�l���^��+Q���V�7.�%�4b9��9쫰dvcVy� �4�*[�PWc�J�R��ג>&P�j+�t�d������2ߤ�7�'D\���D,�G,1R�e?o��dl�H{i|.�Q��K��2Y[s0${�r�:��erA,.�y�}p��'�1�p�&�|J�{�L��qQ�!��6�x������{��ΐS���1����aSl��|��Ԡ7P���H*&<�&�����[��=�oa�:��+T]9��R:��W���j3$ �<�|s�u��[�cR�p'g��:�:���E���q��m[z9��447�%y��чxjawY�I@{aO�5�j� +f�b��<5�q[�6���	�B~6�hv�b%�х���X��J�`��kl���\,Ȃ,8(�)(/]ԟ���Ec)���&B�
��vD<���`���\���]�8�Ԁ�IiI�r�
�;H��B�\��R�A��0lzq�>�r�'�ԲD����xM��Y�jJ�z���7 �̋���)A����f=��%���g:��i��Z�Nċ��]u�J��}���E��T&�<�W��5*�Ď�$@�ǆ�:�dVn[<��0��|y���8ST��5 dʑ|��r΁k1��bLN.=>C��m����x-<<ۿm�c��"j~�b�u}1�|q��j�d���@��+�Ȑ�cr|�T��ա�"��TAX�tc��$;6IE�f;_��Er�A ����v��E���hG�h��X!�[�wI}��H�>�k��D=t�^o�r~J�W���D�P�ܐ�3hRޜ "��WEs�z���� z��b�vQ����������ztϴ��`��P��-��hgU$x��L�R�q�T���S���.�i�3>�~ b�^"v�e������_�zg���_���Z���E�r�b��K_xV'�I�Q�=O�?�􌟡��"��b�m��/����OQG^�/��f�r1��y���{5����,nIi,[�JS��7Ц�y��#K�Ꙍ2xt3�S�O|��n[WY$4���(C���Mj�\��+�L�|��՜�/:�/ϜW�;-Ť�a�*����eʢ��;8"]aWT< �9�~�Q�" �G���5��MB���84ѺN�H�+��Z5=��v�gD�R���	����Q�.D�����x�}�7å��"��璘��}��*����R�:9�[B���}YJ0�W�\�_m�.�*R�������g����y�	�(���NB,�^FB���6� (�K������V���g�3tk+	_s�-H�$��AB�\ִ#k�	�`����EBC���ͣQ����P�I7G<TG)	Ť�$9ÛM�P*��&�"�p���I\_�hCڣ�bxc���a���Cڑ��2���He�1J
� (���u�<]���^ݻ�H�E��آ� �D������(�+�,v�5��%�DI��R'�{T����d���G�\L/l�,�҉ ����yքd=o�v�.���r��dNޔ��۝/��,6����}�=
U�T��������:u�͜�����b%�����d����͙�yJ�g�<��$�O��5%��F��r6&0�*"���dͺ;�5����u����!U���P�D�	78�h���؄���|����f�{�`U�R@�s_C�.��g�u��� ���h�����_N�%H.3ЮqL�0�O6�LrA��P�c�.u���O(g_��9+���B�#���`E�8�;�mk�I��`� ��/桄ud#&��0�{I�x�Z��&��O��!��pZ���*�*�~�;�f��Ü�o����l��	�S�F�p�J��%O@l���3VOazX���o~8"�O��p��ޙ���2���Z��+��82�y.!��-Ej���LR"%=Q��kG�F~/,�N\�m�M?�~,�o���G��_ ^�M�/Y����4��/�YQ-)�{��(E��{B�	G=��>j@ p*|�M����TD��TZ#���D��/#���3����&�����S"��t59I���m��.L�r���D�L4�@�R@^��97Q��x��(2� �,�oaE,|�� :��Xy�T^�J�ڻ�h�s;E�q�𯅚\�,�����lЇ�]+�����|w���3��	�_���@NdMù����Wv���{$��*R6�&Ĥ��4�"�|�h������9)	�a�Ŀ�5�4��$�0����[��9fd�n�=(TFλfs͚�m�pd�zu�=�+[�"�Ζ��� �%�x�A�q@�����K�+#�ŵ���U@���?Y���(�.�㨩����;?h��ނ���6.Lx�p!����*P��9V�;��+M��BA٦��Y��Tt����҄�W�=�[���S�1Ɇ���/F�	T�֏�J `c�$x0C8�S��2��u�knk��Y�O\���S�<�����U�9Qm����+��}�ic+ޗ�%�>F���	���QeH�F��^��i8�<�N�I�Se+�G�̔��:�;�aG�����ggZtG��_܀kcb'|fq[Ǜ]f�׽�����=�vqY1Eb����k�a����5�9��_���5��d�$����FidNY��&�����yX�	�?��ܴ�(��fX�o�bg7n�g�����ES�0��y�E��Y�D��X3��	�8��y�=�� �p���<�voG�� -�Z�!� ��� ����]aי*�sm�F 	���%g�G�9cf�eK�bNKà%�"�V(oE>W�t�F�����J�l�D?��%x!�����& <cc��e�zI�`�/.Η6Wp�R�m����Z�
��;{�� ͓�+*Z�F�9��ּABn~V�������~b�;qe�������O�Ɨ�>~��:�[� ��r|�e�g�L7HhZ)�]����Ҍ��F�Kt

�/��ߖui��0Ⱦ5�Өs#5ݲ$lWK�D7��t�<���վ��]�X*�)e�%�~L���(��m�
F�Dw-	���ְڒ{��Z��t��ǋ�#��y�Q՚�
���7��K&U�m�p�o�������m{��î����������$@1z�.�:»d���უ�9
�3nb?��}����2:Q���ء�+���C�>#inj�����9a��Ø��pP�܃��|�h�@��� 7M���B����'m�/���rrY��]�6�l�G*~A�u�}-F ο�"DEo�P/�}��IiE��7P/ȇ��T���졎?��"H�]�@G#���|٩���Z���E�� �s���j��6>5z��1�_W�eC��L�ci��i��@I�{��%� xBP��������q�?ǩ	AV�h5�N���S������#"<7W#t�6��C�J�����c{��(�J^^6P��i��1t����d������87�Ȓ�
���r��/�DgF*�n�Z0��
`;`x��I?#�ۭ}��"����y�(%VY�K�A���Y�9[&�ˣ���%�0Tۈ�������#�FS�)a@!Y�P:��Q��di�A�Z��t���q_L@� ���ieܛE�PO��6�`�t��{-�Z~j��\ x�J���Q��T�A��M�T�u��s��Jd���&�K���K�ǚM�j)�Z��A�^�H��_�p:'xcq�V_��;�(�|MT�g�%U}�"b_�� T�����hgO+�ԑ"�e�8*(�Yz")�(���{$����Q��6�N(��:z����o� #�r%h�3���|.�����s�_�v�1vy�p ���"hI�<e��_Y���LȖ�?��y<`|�&��Bi�ԛ�I�f��&���v1vӮ'�h�"�6��Q���Q���� ��-�Zy&��>q͆��S����D��:/��D��7.P�_CER�ck~��NU�ONI��Ŗ�]��ɬ�C�3�f���Rp����'<�f;6��ý��V�����r������h�ڄ��>�:+�p+S�E?r�����e+��X���9߱���:p+Fw͔l(o�ЂAΦ9�&F^��2��Q~��a�%1I+� N��U1F���O�w��)�o�����VH-qr�5�����Gs���%���/�=�F�1�Um�uɼW�{���G>,����ɋ�Nh�>�tj�M��Y)�Ϛh_=r����V"B�� e�����*��f�z�z�w%��?�Uڃz��R�U��|�0�q`�jNS���<����|�=��K�T�����Nm��[�=���!�*����F��2�Ru�~��2y��0O<P���cnbWT��:� ��Ty�)�R!Y�>�"��sN�ͱ�N�gN�x��ә�`�h��-)�i<�e�����+6� S^f�?%2J��Z�pS������0�gQ�,#�k@�CE��3�ؼm�4��{��]<�o��)m��KL��U%?�ٝF����U\��z¢�a�Q!`�l쑌�u~G� ֛;�i��w����K	z�8��l��9B���vD<bp5�~����,~5qr����w+#�y��Z��`۳@Ѩ;W$�����ӏ��Ƽ�!c��5x���%�='��q��PW���5�c��7c�]�T�˷�>HsS�y�m���q�P1��]:��;��̇i�o�z[�������鲇��S��%�ŕ�f0���*�����1���JA{s��ɉ����7�������4��A08 ��͑H��a^��~ȩ�5�%���������u�`�G�����9z�ίv�����.�= ���:(%�L��R���<V��!}��Z)Ǵ��5���޳Y�)��EX����O�YQ�h݅?�<F�{��G��ky�	�N�7��z]���Ƣ�"gP󇊯�$�=�RZ1�aT*rL^V�R5��(�^�f�KE/*�<�H�4�z�y�.�o�)�>� �mh,���=	�܍^�(��'B��^�5�U?�'���k��F��x<�� �x���ͺ1|m����GhuR�^��~Nzx�7M26|�� \DG
S�+1O�sl���\O� y?���l��f�m�k�?B:'��0���fJs nP�P��E߶����pr�VIX� {��^��ſ���Q�m9�st����VI�)�5�m��=�ꮠ���B�C�x����)�Z��z�H��/��q�/���_�4�".e�ABP�˞�ԓI��m޾�S'�	vl�W�!cN�=zZ�Q��d4��6�vԌ��P���L�Iƚ]��h�MR�R_���>#s�p����yT4�g�T<Z�j�c^|�l �W�Q�+��
�뢭8.
%�%��k3/\����ƃˁ*��49g�����'v���[� "�7�>29��y��=`
�-�~I2��K�qY>9���]���P�A�Q�Â@�������esۏ��n��M��<��G�$���?˵�~��:*k�3�[}�e���ǅ��%���R����|�˃]pG�M��G�E���������ؤ:i}��{���$/؁�b�&S+e9*7�0�Q���P��ӮՎ��t��s�;慂�^����y0C# ��5��	�v�鹩�9���ÈT%�R�
�s�S�eW7�gQ7l�E�K�1�` =w�:�r��~+ n��:�� �WIy�,���?��C�:�x�H®�U�n[�s��㷒�E��:�q
�>����W�B!�Ӯפr�j#��
HB����J�@�7\��ESusc�������<~v?�����ְؕyN{s~U�Z�źR�~$��Cȼ���$s��Hc!���4��ߙ*X)� ����ҵpVu͂z��yNh����0����pp�r��i	���H�����>W�������r|QM8�~����Ր8�r �'������UQ�~}����8��<ɋJ+���s�h uK)�Ց��ūRn2�xj%��{��V���e�v�i�}�����:���k�����Q��D����|�F����J�#�$V��X4�'��$�]9��@����\?�rF>���r0|�*���L"�4����/x�:7;l}ĵpX7L�L�/.Rӛ>��w�qo���4�!唉5>d�TҐB�F^JK�3���ڕ���p�R"cj������>u������]�8�&�˂�B��v��M���{1}v�� �J�������G��
[�O2@0:����ϗ���Ah�P,U�T�����w��T�}s�t�W}4�{�9��� �1g��_�����l��U�^��ЩY^Xo�4�j(�"�eϐ�?�����mž�kY��Cڼ̆�YuH�"7L�;�Z�xM_������ԴG'��,i뺥	��t��1�4�X���*c��)���Wf~���z�Ţ���_+�W��̆?�<P �r�h�{S�(0�}o��+�#k*(��4b���=����� ^]V�{R&D��V ������ ,��Wp�3��hU�\tEX�i���$��NPS!��q��/��N2����%v�0p"��3"�mVip�T.	+�#�V�u�7#�8�Fg��#�jGǈiD�~��g�V(�.�A�mk�ܹ2 ZmV��zh��w��~�u������B�p+D}h������N�(�F�vR��������	�닾�c�rH�s��Z~�ЪN�l�uQ���t"���Ʉúk�Э�@�^_`���-j	`����h!��5Tt�3U8�9����%+�^���#�X�$�T:�k?���ҡR��$� o��N�F���t�}?��2j'r�����Ѽ�X�s �<�Ԩ��;EZ�P'U���o»H�"��C�N��k��ں������һ���GP@���;7�F���^�4�S2��.�V�@�'<Λ-s��8�xf�tAɇ�e;,+��#�W�Y�ҭ�"��������z�X�������ׄC����dcNg��f�G{&*$��~h5�(c��*a0�t�>pVy���գa�:S&e�v��K/�'9^D�4]�tP��&{���x�&OT6@�r��=�#U���н�3�v���{g���r$�����_޾�h��;��Ʊ	�pM_Ʃ�-w�L��^�4apG�bs�%b�cE2�˨�U�^����4Y.�������ƍ��Jĝ��+��+d��:8cv�-���N"��# �.#�#����v��i0����:<W#��w_�}
��~?�x4�`a!Ĩq�l��=����r�5
�F���ڡ]8j
�k�Y����,ϣ{�&��,i���g�@"���	�$��uvd��g�,oG"a���7����#+J�]��C�Jr>�@��Cv�;Ld��<me�ض �.F��*-@����Z���)˳ͪ�ݕ��9 �^��M�,����UǼY�(�K��?|ֱ*��.5Zޛ����+	:O�(������e9Mo�&��q}�<�ė������)��hU��xm��N���YO�s��oiO������4���{�{�NK���E֓���c���\�L��
���"�?�Ԕ���n!#�Ä���T����G��fQ��<���5���W�GD�YUu;��޺���J37k��E���+n�3�  �'v��}����d)32���B6����8��xΰ�m�Bʲ��-G&�3�*M��w�% o5f���Z!���B��Z�Sl��]H�C)�
�Ο%�>��4&!��]���˔��e��M�x���撷`�]��!-�-n~���3`~<�����4}�6(9��6�b&�i���O���}�X���N��E͇�J��b�#��=�%���)&�F���eM���������Gb��D�"Zh1{����,��[<��P�6���
.K#�QY.����L�v�u��x���t��~�w<�����8v��4pV��>��IК��b_�l"iu��q�x���oS�>o.�Қ\]�4\���-8|
���2��l(y��L�?�����x}ɫg@P
m�٭��}����t�1�~Cvŀ���a��m��$��X�'A����q�Y>�]�]*��٨���:� �|u2�^�-WNTh(`�?�(_�ڻ��,Y��������൨���JB"c�q�����%��j�]��\P.Jh[��T@��u^}W�D��\Mw\�S�(��R�9�G&O_��H�g����Z(��$�l��j�Y߈o `�:>�5�� �M���6�~t����/ӟE:�4�R�]\`�K��W�h��~�L���������*ob�ڰ�����mҖ��~f"��XF��(@R���z�Lf�N� �P�BY?m����9��O��`��"��P��0'3�C7�/E^K#�)U�0���U����(Lwq����n��F�5�|m�P�'��`9_�͌���X�[�Bg�{��oe�rĄԈ$�������,����,���P	���8M��?k�kĉ�H�
���x��1���lpsp��)�����0)��R�-���M��J���

�Z�f��#.��|.���(Mu+A4�Y���p�Fe/F�g�$�X��@x'Mn�]Zߝe⮥��z��4Ct��4"j��}�πM]Eɤ�M̸?�1(���߰�mh�z+ޒZt�3)�(��
Ja[]�;D�$���y��ǘ�T�kʮ
���t�̇����	J1i��<���s���A��;�2�h6�1e��M���|� �6�=�b	��?�Ydy�N�3�f>�"ģYIm*��c�GByT+�����G���a#ů���_{��$�����s���1�U�b��~E`��a�S�"�9dK�!�U�g��=E��Zv�ц�ƌ�saiS8u ߖ��i�8|֔�b�a��^��})K��Q���]NGP�%9���x��.Ġ�S2���=����+��įS�|w���'�/%3�N1�(����.s>��Z�oGK���"�t�������̈́�"J�;l*����˘L��<9=��g,���_{��k� ��g��Ik=U�^�b���ᙆ�'K5ԺȺ�-_�6�ҋFp��Ju�H����̒ �`����x��:��
`bQLOt����Rl�|�Ɂ)��+�=(L����˂��	aRJz�1�B.#�>���}�%B6hτxZE�b<�ld�5�������n)Cw�8e׏�5�%Ky졈]!˯A������ߧ��@��X�"�с����JNe<�����Opܩ^I�b �lw��?id�WY:'���2�x �g����5J[oiK��>>��T /��%��Ǥ����tQHlS]�t��EB���{ f�8���b��.��N�=Rg�Y��,���/N����F�E�Zf������PJ$�ϼ�}�/�qM����3��"�@~Ȧ�nN�gl	�Yqm�i�k��vA\݀��K��#A+����m1�ot}7��6Q�}�!M�:.J�u�����p�&pU���l�L�z`����}��z������)�#>|;�=/�l�H�Dx
(���O�/5ݙ����1�|O�ե����_�E����A�djk�IRz���-��a>�xpЋY�����Z�r��Ĩ䇆�����LD��Γ��|Xb&	t�ӈ1N�}Ū9�0��8����[��P�z�]�t&jb$�K$nF��5����t���w�K$ڔ��' �d��o�ga�� ��Z�~�ff�j\��1_�I6U���	�iݓ��ɱm�w±/�Z��ռÌ��׮e�Lꑧ9Qp���A;�8Z{ޓ�A�ˋ�GY�
-5yt�)��A��0�cZut�xRb\4T�day�#�
�H<O�:�l
��F�ɗEbi���v͚���R�� ݾW���L��.>_���]�#p��b\�&fIea�\3����\r"��*e��GRJ|T�ŐL�_<��DL@/vB ��5e���P%�S%����� ��q��R�t+�j��Ȇe���Q�j9S̝� ����'��j��h�qϲV�V��͏h�]D�l��k�j_'w�
X,��M��5d�p��ά=cJ镎6?�y�肝�!��&��k��`��W 0�����b�-�Ƀǁ�zh����:��hE��p�˓�ǹ��`��9��$i�=���s�J�p<�����|�C4i,��/�"�nE�q.ZIu��Q��;�̆J~`6������hҔ����9^��]N=�lʮ�p���
�	��Vr�4��rB���(p�H���^v���i��^�s=GKRv�:L���/};̒u,��D���=��$0261�k?h|�P�_ u��`��7dsv��Z��n�r^
���
��E��vD�)eS���ZWa�x �J!���k�_ځV���h������!k~��<{N�1�%z�a�K�a��6P�0�*�B�${LDW�g���zvC?�d�U�A7�$U�m���[r�)�g������Yo {��Xi�s�Xh�3���C m	e/	;ꙗ��2=�k���Oi%t��綖8IaW�>f	 ��k �Rl���/tW;���#Ůyd<��Էu�M���_|�TQ����[qF�	����m�k~�+�3�	ͼ	�zo����z[y�3:=偓����=,�����6��Mtqk������ML^�����h@N���G"�L�ˈ���g�=�4�C�9�R��$�ד��pH��Rf�,�b�<�֯]BM]����2�28ZX���V�����$��҆xT�H��n��!��J}�ӛg�H�yN|��I}ٕ�Z����!����F�ƨO��������ӐZN.�Pś�ZԚ��mr/_)+��fi����҉�g�S4`$�Q���M��y�0Rb��G<%"qe-�U�+�Ƭ�1���VlP�l�O���¿�Kx�^�a��9F00C�X%�a<�d�n7�iޚG�]�d�Y\�4DJ�tO���h�g]_�՝��`���H�����W�6#�A��ӝ5��la���|��	x�`"Q9��
�ӫf�
}3[>傋?�!V�*I�ft^�!�K�P�'���s	��/�"��;���_��:��Hu��)��+q�]�+�%�M���)G�|��n:>Qw�a����Ҵ.T��3��u�<��_�$3om|0�T�3��MlsJ���[���,��t*�Y����?����Ŕ��&ք���~ڍmQ��^��(��;&dР��#��b�X����ߌ!��ޚNХ�ƛ�t�bΣv~n��c��7r�>��L|���5z�zb�n��]��Rg����O!h�)���{����i�O�s����si$� ى���j_�~	5���]����g��r+A��6�f��H0����׳���<~�w�̶� �k���g�7��Rӟzˬ�M �t\I�Ez�r0b�5WG��{(Q\�H��U(BqT4Hl����kT2�P���R _����
$�+�o�z=���F}m�l0j՞������Aem�����Dn���=lI�E�mQ{71� �ٖ������G��.{x ��'�]�Ѣ�§�	�,sR����~��=N#s�^�g��������xV�}�o`ݡ�C4��@p���g��.�D2�&�!A�{喳�֒�JV+N�9ڡ<��z�@s���rx�;���0��`������ϼG�^��۳g�`�5b(���"�I�ҟ-�Ə�J�J%���k�F-��˱_@H�\]?�%Mb�Vh��l�0����SPG���cqo_��EÄ���o�`['s���Ϧ��ê�F����<���=$3F�zqI����&��Wz�8�(=��CЀ��mSg+��Zޥ������ޕU����xC�3���U�BɴfJ2��@�w�����[���1r-8�aX*䰥��m�9��Yw2v��S(�3�z"/���#+�>}n��4��۲��V�S}�=I�Ly��5��{��Μy����az5s�D	gz�����ZF�Y�{=X�y�!�!j,�HF��1�uG���̲�-�jC����u��d�$otC�ǯZ �o/�귣��!�\�?�wze��&���p�(�D�P���K�3��␐�s����>0��9���l�ؽ
�-$�d�8�pq*|K8�����~E�H�Uz	=�b��Ýxyc���t�%2?4(�����u���U��6�v�"v���17��֦�..o��9H\h��;�r*��)LQC�I����b�u-!��F5��>�I��}�>w��.x�������������JV���Kz+�_�ГƓ�3|��:��i�����"\�1�R(4{yro��YP\1�KLGK��|;�jk(�������7���Ł,���f8J��*�T�����p$�E�y��-^���`����L��n[4�Մ�㻍�`h�D�ԂM���F����3���!)�����B�dY��{��̝����~��čr�cm��_��ț};�>4��`�
�C��q�f\QݻT,�˲��g���6Ӟ�G2'$R�����v�aK+P$��2�vҊ�?��fX|����6�{�$����Y)��]�W짌Q9+ݾ�@[+��{vS<�:�ݗu�D�W�20[��N%�Z2^���s4ba�k���;w�^C�H�BBò��R��U��T�p��Xy���
Q���ㆾſE瀁�i?���i�\=�9Bm��E�l�~ �V��xE��� ~%���fI7$ʭ^M�DI'��6���x��>~�fP`��"�H��
jm�����>�a_E�F?���"O$Ed��h�N;ϋ)�]��5;XM�]�>W:�_	,��ζ���Zy��ݳ��Qp�35���Jm0ZS�5��2T���U��|DA�*P��N~�^PzKe�҃N�P��+�&	6;o��}�I9S��K��L�`�*�5�����j���w+��Ϻ����`�L] t��������{Q́�Àt�T�&QC��Jl6�c�F�
qv~�y�v���fI��')�r�d��=����Iz������v���h3�x"�|rﵦ����[_�
�XLS��
N�]���h�:���?��� j;:���A�0����
X�yݜ"ǚ��9�c�W�C�?=�*�[,����^v;��Y�X𒏈�H�ǘDٯNw�� G������r����i^[&�.4�~ۇ�� �X����"�� ?���c�,x\��[+S�D29��Ǵ�Tˉ5��o�ES�oN�Y� *�
zU�k~��5���B~��:}�whB��Іq͖I|�D=`�01�n����Bۨ��w�,�ODs�ȅ9��{6 ^���AM�=�	F$���ȓR��~Z�q
��J�p��S,�s��e����B�E��>wø_|�Q���(	�w��Lc�H����QgJ��g�7)H~k���Q\�/���A�҆\�����n��0r���^�0�S�U��b���� ?��9c���[V�dW�c�7�jO�2��pK"Pn�����M�1=���2}[��TW��Ƣğ��촟�ܨ�c�[�ЫS�Gɹ��L���M\��,���3�[4�i��a})W��]?�^�q���î�ٲ�N�Bo8�Wf�Α�?�b'���W�;@,\[��{�%�ӵKa@��7"9*M�P�},��W	�r�� �SO��f�g0����^q�D���Ӈ��[�v��OfUp�*��#1�|D4��=�5�j�$�~��\E��b���=Σ��j=@$l�)>D�r)�z���~�V]�7�jܸԬۚ
�85ݦ�xV��T��\"rٱ�=t�lpJ1�+�s�W��S��okI��/�?H���R`�}�#�ǣ�|0�� ��ý�P�s�75�EA%(��FewTj&�`oL�y��ኦ��'�L��t �ۋ�+d��j� �Ð��8-�[�Y�u�K����I��
􃃑�8m�S�㨳.[�T�85|�.͜-W��8G*�:C[�����NRa�T����ħ�E!�\�۶���Wn
���/��� '��Tg���:B��m�@���4
$\7@�ǆV�j��)���B!B�(�#>��Ű�J3�O��	L�a�&�(���v�+�o/��1_��!�� �J�>l\�ia��~�\>�ra�-�(xPˏ�Y�P�a��7��%+����ߍ��x�-f����3���'c�gw��
����?�)��O[ȳ�%��o9Lk5�����m?��H��]��΢���)\���xi	|��� �h�y��-9�He������TC�"N�`H�y� �K�q�[��l�Z�������t�6DQc�P�_sa�SѸD���
|y��jbڙ���n��O�o�A��Ev�A�yƎ̙`p}�7.�u��W��n��?�1�:���b+'��R���N;���t�vp;��^�@`�R�e�v���a�j 8�[W��\���],J
h�5n��a�!�u )��.;|1��N��C>�F�m�����Z�]�ǟ�^�� s���lծs4�4Eu�Tf��U>�:�Q�
�@y�Z��A(6@^�?G��*p2�Ӎ��!y+���ji�8%2����(��<m�����?��~�!r_��1�ӗ2OP7�#*�O�J�h@?�.�N�ۜAiz�;[�}�+PwD��_���b2̽��4����b�4��(��71�? ��?�KhMc���W�@�֔�s@_�P��5��'2`�b/��o*0fw�<?0��2��9t�ľ�����?g�D�P�9j���R�4`^�����^�/�����d#�w�n��B�Z/͙���������O o3�Kw��x�pv����6n�=x��M�g����@���)�%�l���&:K���%Q%�Q.I(�4�B��o���@�A��Q![b���r��OR�5��s�;�yz4N<.uH���m�_�S��n���������Zc|Rf P��9|�A9'���g\ҏ��~'��n'�,C��D�q�b޹\P��ɐDF;y���F�[;��h}�7-uM���h��JU�H1Yy�����E�^K٦�m�ӫ��!�Ϟ�@��ȓ�/�w�#�V$2԰��?Q��$���������RDk�1<��w�cVJ��%[�"eW���`��ic2�=L�����t]�*�湀S2�z�r3�(7�W���u�s�@u7G�*�G��Z؉Ts��x�����v�y��h�^�z�������I�>/B�������;����t��DoS�՘
�L����l�1�pM5�X���f��]���<��f����<��Rw��?��g��Z>�ALKƆ��6��Z��8��_d�d5���T�Si3��sF&��b2FI*���Ib����CQ���l<z��{��s	`h�r���	LO�/{ޥ���:?M�]���-ٷ�]��<ǠOj�-%Ԝ��J�D@"j�UDee����fw��
Li��Ib-�-��[.t|.�v�wݷ�)�`T�ItC����,�� ^!��g�1uiM��
L����ə�H�z�p�i�Hj������~��>����]��g���E2��H�\��ƨ��y,G�$4G4�L�7�,��Vp�@'��OBb���D�iy�$���p�X��7�2��]`9�p�=�o��y%�����4lW�����֥�$���O�i�?4��H�T�#���hǄ*����^�1�`;mZl8�^p����XKm,Z��'�v�0�����F�Y�G�o�����D}�8�`�ݥKZ�����w��m۞����@X�Wf��t�{��p�a�߷�B�MP��bl�W�^7�ss��p�JU)�u2j����T�xIZ�]o�c�R��`�������vF�^<D�4@@_��a2���8\�|$O�DB�c]�;�Xr)qO!_#[�Z�Qzʤ��=0x�֟1����6a��v̱�����㞄������%�Pfe��`��o��ov
�\g��~D7޴z T��$�����x
����&6|�s
1����a'ms;�s8��FF��rpI-h3���U
h��:�j=���!a���5�^�w�ۙ��������- Y�����o8�0�P,e�x��!�KZ�l�d!��c����U��1\��}�wr�i%���T��� L����'&(_&Z�j�"�3֥|�c� ��a�ҰQQ�ǁ��(��R[Rе+�6J���]�'��k�J�����0�{�X�=���kvX���̓���'�4���.b�����	:EyP	�b����42�8>����"�M��Z��K�̣��X̽�KL!�>���j�f�2��A���H����C�癭�!!�*d��,�''�?N1��/,IbZ�}�u�bC
���;�� �@N�q.��(���@�aL�ј��W�&�t[/�m��^0n�b�XM���L`�J�\p�@h���濾F]hM?���b5��!��"B�� u]}'��
T�#Nv�A��*/�~�vEeF����8d�J��������ͧ��O͌���u���*�!+����N��7��3#�M*c	�In�Z���������~0�|��#�B'�'��<Q$�&�g����v2�>G��������~7Hq��&&Ԧ��;����0sB��t��)��I�\xm$�_�K��EE|�Q�kC�]`���ƞ5Wv%빻v������ʀ_�iE�!��[m'�[�i9LD��c�J&�gD�n��s����'�{�Q�����.G�T7B�<$���|�Ny]Ϡ��!sw0w�dĖ9Ym����_��Бa��u�4^��π��f�&x3��5�B�������uv�6�8�>6��U(W��?��?xVVcH��\���T� �~o�)8�W��+ � �^�����0�g��u!ˀ^��"��v;�pd��m[�K/A�`i����L�.:���9�	��s(*fcu�T%O�t�6�n�ű��m��˘�|W��t�a<��'˴AJ���p&S�K��~��!pȴ�x��2�i�2q��(o��X���gL�@���4"��'�$m3��O�W;�{].=s�/���.Jg�јm�8�5�h���zH��#�FεQ=�^��K<a��ߞ���`�/|��o}x��cÎ��~4�qp��R��v���c�
㝖��t�~��ٯ���wo���0�մ!/Sf�vda��۽|S��pn����`X�#��e4L�\W�����}�o��¥q�Ǵ�GEުQ��L�:��c	l����-��LJ�࿮�I+h�\�.,�o�\)���
f�m�#i"f��5v;�r�/�q���[�e�A�iX��g�GnsR�.~��)�u��x��K��^���À��^��VT��IT���n�[�mم�)����X�`C�c=:����,���x>YR)K7�AQ�Pz:�|����$��s�`�]�쇚e�'��Où�����b��W���>�,*a��K�Y����W0�����Ա`���e��62W�ABvh�[�l��I���:�𖡊������>ـr���5L���q� Z��^c3�ph����	b�`�Zڄh�N��-IAy���P��0Rl����N@m\��l����E?���Ö���G�%�nQM3����N1DD��'2y�#>~�����k�
G��4~��ki�9c��i]W��Ǥ�؁+E'L�<zA�<f�DpZ���FVI����k�h�Ǳȴ�o��lR.@�_,K*$Aw[#:���V`�X�М]k:DT��f��Ҟ�� �ξۮ��_Q"���D���Rbb"]�f�H�/t�/��(�)"L>�d���r�H/�4�o���f�#�� ��8�����e�ҭԗ��xL��16�5P����oK����e;ѐ|�M�*Σ����;�J9�U�2�r���?��h�l;(��ZB��m��A���YU��駼�Hd�+`�hM�,��D�	���Aˤ�T��ǉ��5Mr<��\^�T��Hͅ}�th/�l��a�8"oĩĿ����da������{h�8�Hvr��㤉��s�A��
����3[.P��z�y���+w��vp���74�t�����0�3'���2�+O˘:�Bt�?Qi)��!*�L�
HK�����yV����������,%��1b�_��KG����g�N�M�cP^^BS�Lv�abM�iz���GJ�۩�.���8�ș�ʽW���ߟӡ�a�SO���3�Ջ��ҳNK�34��Q����.\����z<08�h�f谽��P���E�y��G���쇱�)��2d�Ћ�S��xٌF;�[�%U�[�L�9��s�3��K�O��U��
����iSr�A�֓Hp0�ٯ�,Ge�������wS:�#4y9u�Q�o@tN��)rCD籇�n9����R�׾�T��߁��l�3�ˣ�4�c��i��� �C5�h<��
g �]��(��hZmR���[�w��3w~��~�ƠB*��? �\$>�U
�Jn�b�^و���Rә��k֮�e�)�&�E����;C1К$$e�3z����L:_��}�"����U��sz��+`Id���LS�����Z'�`EB.�b9;����]rrqL��{9���n*�oHUm����Ö����Q8����[:1h�+�P+��s�l3V���;BǓ���H?�8Y�i2Kc�YK<!����-��Gnm����Aa�h1��"]��05�8���~k���+*.�<�e��s�JIJ��e뉓�!���?�מ
�9wK|�Ks�Sdm:i�Z��#=Տ`лXm�޵9*��h6¡؀c�T,л�P�5� c�1O��bf������Y^�ǃ]� Ym�v_L� ��\��gVqڲ�߱4)���J�)��c�o^J{B{�kS��kU�EԀY�c$�N�Z����w%q��o�ޢ�����n�즋%���Zaښ��A���k��J|���Be;[�O��09�X6b�8����ݡ���	�-�n�����7���]jٍ�����7p@s�7�t�@���G���-`\6���`�P-M�DmZ��!�2j9Z{8_�8��j�q���@f��C���n�ܕ��u���/����ӆ��Jυx�Np
�L�+%�0����.!���O�1'�rVUyj�n�qqqU��*4x��}�n�"�Tsh)w�G�I
���8/!�S<�PXUr�¼`�x��V��*,H����圢G�+b��Yҡ@��0v8@rϢ?�凢;�(�κizSy�*��[�REM͢�c�X�u�y�U=�6���ڴ�JHߔ5�?�Gf�T*�u=�d���H�c��^�ä��i�.r;�px�խjܳY�M^�C���l�R[��Z=�[�Yl�T<ĕF���H�AN����k���-�ʕLR��mo�+������ �,��;�ڤ����lV*��%�����g��y ���}�lU��	�bU�kQ&Dk��wX�����5�O&D��,gթz9p�8m��]k���v��cF�R��~�<R���u&��x�/T�d�0��9�}�؏���ar��!F:�Y���;�V?�ߘ��BҎ�ݫ� ����8<i]PJ#�PӬ��zr�s[�����J�_��q�±�E�#J1>8�k,��#3�|-w�YK�Ǝfza5��z��ik[��'	��6	!�lK��{�Qe9��Ô0�ߍdF|�e QG�3^^=��.S���-�����XV�Z]	�O����co%>��/���]�/q�G08ܚ>�%r�Qt�`���:B��r	#]Ń��9b�2aAgS6�`չ<�Sm���9ȑ�y�^E��稓�KF*�M\�S�3�/�-<�Af������,C3�o����TL���ӳ8�/��B�*� oKܿ�,�phM+ge�	&�B:1���Z#z	5����'Q�\$�ܝ �S|it�c��(�2�4)/�{-��!7#e���%>g��~��� 2�lS�e�#~L���_?�6�:-y��1���ݫ�~�����.pE����G�E0�4�_ẺF?"@N5,z&�J������h�UE��r�Y��{?i�M��P��=6��'�h�F�D�t�K�=�������v�X�0���1Դ��Ͻ�	�T�Տ�c��]�S�����>��� I���)=8���:�� �F1���R�ٵL�u�'�Laj11�*�.*Ni���b1��G<�d2�⃗�c�a4�����J'���[�T�}�5scI��g6�kH���fn7&�|��aUA.4Q�$siܨ�M��҂{����z�ڏ��Tp�����VCrOgv�0�+>�'���pd�5�ݼ<hk!��N�.�:K�i٤u�/ǥ��\�'�%�O�I~��	p�S�z0��<;�R�-8B��?KD�4nx�=*�I����Xݲ��{�LB�G��aeY|�Sb�j1d�弗��~/,)\�B1aHe�있J����ފ,B���<���kĨ�<�FƔ�Gc�� *��|q�K���,�,'d,��p�KH�t���"�f��
��>�6p�c\��+����(��y�/<�Ҳ�+��0����1Jql���e����U]�����F\�7� �R%)��������q���]��'y'⍝;Ju$c�G���A��ڋt�6F��	E�*��h��)����J��}�m�}w�7!\���k�r+�40a��n�]F&���K�B�f�yZ��
���c0u=`�N���K��,�@E�u[Q��1𴽊� ��f�^�9__�8��P�7�	(��T��w�����c�pU�֭��*��HZg�̺ʀ���V����:�DL�E�7�$�2�v���ͥt�G]�{��;�O��>��3U����H�|d��,�b��h'��Gg�;IA�v�xK쵅ݩN>�N������w�u͐;kׇ��Ɂ+�D�)��s���[����~�U�&o�;�na�Z=;�AN������NJ؞'K��WD�];i��e����E,�n4�_��`�S�����p��NLm_��pV���)�FH�#l2H$�y!p�JPV�6ƙ��,����՞�O��(D�+����;�82��6>0"\�����G�(
r��Qf�*<gR�+" X|ڢc~��,DϾ������O5������*�Tx�'JjJb���� "�M]%�O
���j�R����7��m+�.��W�ѺNیh�W�|:�����T�
�����/�{+:�ۻh��/�|j¬�F�d�c�_8�0��r�x$�i�Q��g��I�"���r���=�}�$/�J=���O����M�}�#��`wN�������u���a