// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
I5vYEX4sU/Md57QQFqH3Xij7GAMPSRagkt9Wd6Yl3RDzVgEwNAM3/RJJyk3ngJNelJJxFIaBW5r5
yD31jyUO8zEkyywpw9Kwxj3dhJGzv9zdLPf0C9aZ8RAgZoZiJLm/F0rcdbURK6XLwQ5u4QcmPcYE
PGXEAtJ8XtdAqoG+vvn5dY4Usdfc/JDgcdbt8oyKDDg9JRSeGy8H1Z78oUpzrP2KACKpRGcnFXKe
CouXAGD5x9lIGkZCH//+MPxyvPsJNM5flJMYlEO+3go8VSR11zl+DK24o+5jAiHtFffhXIeErOub
kJLK4MPjp04sxjoOEPBFjRbQBUuBq38kKTVxAw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5136)
BrU9qKHzjvPYxEJg0K9vl9Wf98edXXazsFo/ufYdC2QonFi05lT02mQRzjM5J/UTJenIjnFslC8N
UeFaxGHkHefJ645A8UnRwD0r5Kwge8dPDrdc6CWrIWMH27TkAdoxkGfWDrDRAv8ZzR6zDJLedYZd
rIvPRaoTgWFoS/CdZA5v8Ec4gb7bSmF2oJhedOW1zpSU/9zLzYpTAFdv7J+q4E6H+R9/qnq/EGVP
Fzn6l4bXEns5pwH6GncpY6QrqI+8NG2Eoik+Q1RcZPmsKyrA90fEfABdhLkUqLirtLaB5UkVv+uI
1CyjXmUdIvahGc3UKb/HuU2V5f2/L8gQejGpkcASJAP1joNtlFxWWoN/fxSYCdsA8KNhAkKbJSvG
cGoYIe7gGiR1odrkU/w0TCBAYGElkkl51hLTbAgwQfTjjUoJM+gM/AXA6W7eRGhLxRM68qhFEExG
meuHEvhR/CRdosG5Bo9vK+ekdcniwVOxnL5O3mHfyIO3kqpLcLxmOyFUNxwrhZIT/HDlDvo7ygeS
4VJM8Af3YdZMJR5kMMWb+FR/ee/QLO/RttlT3/XY+nyhbRt1DvZ8AqUuDDiez1X8qKR0cHYQWw7r
QWOCaUv+9Keq6yr/nsZgF0sfMUpquhxNG5aWlRJTYsQjoXaUUN9ifZTav8MRslbNPm+VVlaobVCr
WWjR+f2ja6vXI7YaR4XwtpzVR/Qsm+DaiCU883UJU0X2Wk5b/qNoC5CzKF2B6PMuj5K6AqZIpNSF
vDN+8GqTRvl/aMKlsXNw0aXamUzD6OgRx4S7hp7bZD9jSLVKALElFMHtmagqzchVKePfDHvvVSna
ep4MrZYLHfcYwXPu20Jxzs6HDpY4CpHTi/CkrBzcBq2OKJwxI9nzCJJbeZaDRg5Q1YuJ9mwqmMB5
VolqK0rNHijGVxr643iM1MRBRaKMGg0ZvWBR5DRCR00v/9hitKWBDcDrHbYtXF3HKeGPVeTrzPDe
bX7eCBZ5iORbU3DffZS/fKPY2WyNuPGPORX7xkzZjj/KXJ0HemSgirIfP9q6CRVMe8p8+6zxkolM
3XhsULvUxpPCQOvVQr5ty1CMn7m3Erq5oW1iUMQXJvM9RybvntKccYhu9AgoGy4zd77iZ3TaDjqU
kKD+OR+2zgQNOkkZR3LIQdImBC/QYzjr2jL9kUh+a4GFinILODP1Lqm7UPpuUk8X5WgtMOXCWWBN
vkAQp4SquwNtNBEFsqoX5YJa515O+42fYnKWQ7pUGC6lqBlePdBcvueDsuTAjvw8d268u81L1eLy
ehPmZ3qlGNu9WppzNIp1ogH82RSnHWlzPczwCodewMPMw9dj6KYzu7oFDPUmYeki/rBkiuErDPlq
L8MFahtfOrfXx3Kn63abwYSsg2XBhwKgz9ESEq4PobVJk2S+r/NhlCy7j3octfF/jGv+7HejDnql
cbs2A1WUFJoBWU9Ejrvwg4kTdHzG5hPWdO+r3UiFWpdS9i0KQyf7ACMRGMa1v0hSLmC+JVrAMX93
q+ZMsTUR1GPrhEt0wS5colJGXFpDpMEIokvcIDA2Fm+MryefRdDLVNzbWASXhL93LpmwP5Is3L9d
I4wmdFeM1zgpd3zmbzleqjRZBwuj5/f/1iRGQljWobzundwjZ5aKywrv1d4b77u9ckU9kkL8MhpE
NFuGyI/F1xB9AzwFspEBIDVUjRTyXDyQ2ptPvEVg8/LlqQ8KWM7Vo+Ezds20a4H4d2aszQsaNTS/
0ErLdv/FtULgw/m3m1rvrZMlqAYopWZTHoAC1m4hIrEXjCspr+42OM7WUEbfYdFTNEyCsDWdPOFJ
H66v2qs4nCPVhWG+gITBIixeyIfWaqIhBQTVHSV00sc2hxeMNzSDiuuHqf0XhmMYbJqoY5NaGzUQ
5TDB7IJthJX45+eJycnvv23I+xM/4MnMj9hl28aLU+CIxCvzcrZIkHcmp6qUQ9PZX3AKKNxmp9o6
SZF3YjkxgV972eWDom4MpcpMJUMx6x2332V+reaVsp8AD6ZlZmTJUg7/vePVb+sir9FOeJ1K3AYL
hjZ7isd/YnycrCE5sMTkujmLpbnD5yCxfNFoEsxpM7Hi3NiAoxJ447DVKRbcsu0RzTsr9HddPd5V
yZdVo2WdeCiaPhnbqqHstXtV4USkCfn6lDVab5wIAajD51XQqnoedQo3NBmem+eUL+b5uedDuYvs
Z0E1c0erIIfksqJMmX6zG/y2ZDLor1YezI2ZV2J9be75pjEO09vLxgvR6vvSS0/H1P0WdQhACTH9
VAc2Glt0HOxUC8qMbfX6nuR4i/9wI/ITYrf/xbSg9jUwpbTDwXMSQ+nVZMkleBad169u1WvgDuv/
6eAK+PwVM33AQSu4f418vb/zLd3kCpVEaG26tBH/6hBhJsFkZCN/IQ72aDSZaiqn3pbBqCJk8XLZ
5SRgzMxhSdhjfSVb+zSR1UomziXh7CNEMmEYV4y056USbj4soms1upGSr9MZGZqLz0T/CZJTB6rA
2EoUk2Ys2MdbSDPOib7V2SbUcYTe45oogYUlDTj610qY83da1FcUDLkGuzx1AuA/SWla3f3rJnGW
F370GVUQ0PKT6iixt8E/SwkBEtBZq8y5T6nt1vU7rTFw5oaO75iZDcQPZlvJ6TccygcuKgkzxRRJ
D0IgaaY0PQMPuzmhU76WDT6aGKxGROUWJBpvuy66yvkIgFJpGYM8z1Ku0sIuDT+3Am9xmD54VBnx
em9Go2j/K3qWVZLcvfkNzin9jxem0D51tnfDNpQM4fOhcCtG+T2avoMfLaxntev8rSsXg6kKVNwr
MI+wZkzeh91t4o2WNVuqu2twJV7wGfJ/XS7R1/Z8y9d1qJOEmaJugHwM/oDUocLwJQt/gwO98jAw
RFui3wNBtd/Pdxlo1y2/pC80+/hp0CO3PrMAYiPChkOYDIV78Giu6qyDG77AKS5pKoGXK67fYpfD
U/ZK7Q8QrZYh4tkpLwdHfGSKL6yps2qRgSjTaAjgIc75czE94hnaEOZE2UnJf2iBmQ9SNFPpGWNs
eO2XhYchlUXc25EPJNrxU7kyf9Q929PUON8yMDgcdNjvxTC4vad03BeDwSSs/51VXYGXm8pmwo7J
a072HLaorNSkjmUCDSJkQoLBxOqz1ObID5JsOKsyqM7H0z/jwjsfeqWXCaSxFUkgD6ULDM3IMs7c
mvVJmfeexJXjGwbUHhUsQ5k5pMn7rD8zc6cl7jLnmh74uEqLiRQ8+67V+XYCywsM0GyosHqJWWAG
dwnU9aT6aAujfC7bqAuWSvfO9RyFKqvnVCFBGTOAe70rKs9gh6hoY51+2zqtORl5XqL+DfZUDB8a
pyrAVygqTl7XPJF3EhX28RwQPF0o0vrN2z0dY+SJGHYqcpcv/S4kC8fB+92yr28FmkFYkfcBSaX1
ZE722WYlq1BbWIwgE+90sBjlB1kXsJYns8pP626/uAiQDS7mCKhCNinIvIJtQ75Pzwrdpsjc3LOZ
AzaxvOU96YdgsTBMfxFTbMUQ4O8Mj59YxGdchy79v5HRxQTQ07lb8UUeZfPBss+u2/cyv4tu3ROg
IFteeZMV4Z1gjkAxSmRBosE9Fy+Vk6MsgdrJ0sJ0/r+2AQKXoxR5OO7+hRzwkuQN8K5CYGTy2XqU
wocoDhO+rGfbpXY80AoHF++HEnkIMcwPMWn/vLo3r2N/l8r39GbTv1pNI8Bh4m8iJAE42M2J8L8P
Rc/JTuQv0AtKm3tHoJ8qxD+v6rBKqyTViNTlIJla8CfG7P+sUzvyTIEXoUh3Q3MT0y5tTkd+FOhN
4mGsB4zknw9SYKgt+EDnOVbZLcoX+HJv9ydWJ1Pi3zKc98XaXeFgVBHu78vQMlhSpnDPif9B3Ow3
54RJ0eJm/3058K7tXx5xaLZQKHON9rFTTVP51fnyKioiAA/8VbMhCwU1O4LdgA5VHpezOLNFcm3c
OUEmJOm3jpA1tQxqANXN5jQLUy2pXnouZ0rYXYdZaHlsE7HVLCucvSOwRQzKeVO2kh39CviAkpCB
WQf/chel8LozApiLScGWhrqzRbPAJLcUwjpHNJvUlPvkks23t2gZANE4vRQyhLtqEpjREhot3gd7
44XP6N3u42ADhbgRKcIg46HZCtxi2HAfwgwJFI9ocnPEBDpEi0g+eWmCdC3FynpMYA68DDMI10ZI
AVDj0lkDoHOoSBCxOigojHsmZf7fkoHjQQuXKGCmiGceTNCSjLr//MrSnQ1Y7Orw3SEF3Z9Zkxse
t+wR6giE+q0KdnWvjlb43SSbCsms99sMkOixIdC3xiNVAbG1Jg3eUCS9QpBdo9VwG3YuKr3FQezz
bwjvkG8nG5ZVJUxwkbynFqNsNrKMvpWKV7LBJ7YpaFyvjrgalhB3n+uT6XtoI3AqkOCaKqkYLVzt
YnzskIb+xj+Y2F8Zajep8rgE1E7JsbyMAeRCbDPwrAKOnyycxWiJVLMuU55c3q+50UUlRKR4Wvzh
rVygjMOOJLXe0lL4Frf0yAZXKbR+99uBS6D35ZRE0dSVIyakyHlhwpIgJZDl1iUmqWpz6Q0u1IOV
yYxpOzLoLkmKQE+Nmsx0/w4PSF991p6pjrlauP2Yo4AJjmKKuDIOJ+tJOFqMShsOxAKG1X8h3xUY
TmG0sT5LfrR4MLGgCRHuxjNga1ennxcYg43qh2Fnyrff/R6JQ6m7aBC9RuvyZlNOwtb30QEI/mvH
l6DpQp6SDd6mN5CT5P94pN9qvBkwviLv8P++PVaNwLkOkBB0C9mXwyQ/tPuwbfpn9rvLYc0cMMcE
l9giQJgOGKM4qKPFbohyKOvO47sNxamhHiny7RCyXVORjmrp3BHkFYyiWq8DDa/UqmvepfAph+xn
aTc7QC58o/Lz4GrUKVnnQOndvPy+owYhryBsdqIi7XdDwkP2NyJ/Jx208oxF6BCZCNlDM/TRHkG1
vqktjYwBmnkQhGXHcxQDZOWaqUzNNal0dOyhqiwhjSxuqOtLWmy6hN0jLtsvWhuwm6fQQ+oOFyQg
4VXLPwRUwNR03wQmvQPK+f0Dd4Rs5YFm8MTI5sG8EYq9wpzNZj3J41e1Ex/KLBfhzUWMazxl+GRj
XkmXXaUDtrzis6MrVxuVQkahn7BtE5fQxAE452yfczUfnN0rUK4O4H+Gx7ZqxHVpehQApGNufH1V
eILWm4a5a4XYDrv4OEOH7LvqhxbhabUMgAlOCsSWq2E01oVeDNLWFKW1YeVq2T6If3qaMA5uS7xH
7oNxUeOmK303q9iPivn2hEiU/hLj2jS7tfeaFNNrQP7XmwjRU3sIvMtDOh4GBk+qAuD87dY5Pr5h
dUq0uHJc3MpAbhaI4SlTv9YsU6F3humITtU5pbw0JAHUqT4QdwtVh3Q/aA9ahsGLTvj8FPKIoc+8
TboA2lMveHAUZof055uxr5qgj0A9tp+JM0twLz2GOQL/2FhatxaUlYWOXsAVIPjHXOdubb14I9ry
Onx2rZWt8ULeIeUn0msj+lBcDMeVKhhusrOWguITpHJiejfKcG+IQvmqMcTFFKnHppdjSXTkH+Ag
gwnAJMyIdc7B4nXUrSLes7fnXLj7ggUCjD4Ir2c+9AFL/iF7fXQleVl6Ttp9wI+1tylJRY8achpa
yYguZAxATpCb3j57tyiydPcf93XCa5IfSBBPGIvN0dqRFORb8XqQVfitb47xXYdo10LPDKFe8KPY
C3BtERKm6V6pH44MSVr7IRzWF5VZdwSqQa5A+AZm3cBqYsRAepL6nnHPZAO0zJO2s7nRrdF+76Co
T083qrJnySpdutr1TsL6uXa+z6zUg9vdlQATXXsznh5Yky9NSXSpXVPKlmF/JxoItv5ArGLLCJzj
B+k8vFCcKeIB0wlvUT+xWevgc31BaVEfKAgJHLyLRUjEGFGUE2cQ+MBNT/ziIBdTpX0MUzt+wjCh
IutCTdaw0b80yvsYBagNylMbDTn7gmjVI+KW/WXzAN3nUnXu98Gq/nV6Vd1yR15VgSnamfN8oRE0
4xDAdu4JOJ4VDEeYcW30Wx41jBuHrPZkG4aM94MinkGufdTMmrcmOrcT5s1G8TDKUs+TKRV97IaP
6AqFKNW66kOJe+o3doQtiqFy0pzNbcVDLPlIMjfG7Gax5U+61R9WlvmIBVY17KEI+zGWxgDISu66
SKkel9fLKq1MmwOVeIGo/PiVIm2nhuNjJ7NeSf3IJPPiI/6iaJkrafImdbtbf1AJmWSZm/x+/hCL
mmJhUgI2pV213mEGIBPu75a/Ws+Y7IVdY7nPi5SQKqF+jPg9Jf6N4ajtEC8ugLbs1XsiWQrprVjI
hcA4+CaNzbIhuD+o68qcJpYp6lWe8BpgWNjQvSnhC5+4VLu4wP+D8ZuG4Dzs9l0/IbBRCF+Ey4k+
L6H1bI4Xa4r9PGEwA131K9adJqN6StkfjV+a8pjUst7pt3n4zW4qD2hK60PB35rCZLmsI+Kl4qEn
yOqPxrTzyQEHqlPImqxmCTStp0dmLiJVLBQjskAw0UhsAh6Y0AObaqUMSDVq+qdlJwVaZYxE85dK
pBSOsHW9eZuansATcMMrYrbvm04AcejQbwesT48SPk/fJ+eXHj0/xNZ1Rp3GQXKmpchvZcXon+WR
JVTpvOcxnZNruaS8U6HGdiucTkoKAdrBZHOUdT1fLNRQ+oIpUBoPWMDRLMk4aSJq+MCwWbsJJoGb
oEjCiH+Ecs83DPS2SWQXl3rbCpwYm0kf1NWGzA6pC4qZY/VX4Q2Rzs+cxXtekEWei569SwbswaZe
aF6XhN4XZZNgebvJzb4BncX8TmAeeJxzSIWjQp41/HJRcrCr7ruGYmsmD/CjbTz/xHw40fSxQvNe
Ke1zJg/J
`pragma protect end_protected
