`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eFyx+i3RsPoH1YpM67oz6TZ10Wr1k6eumDiffT2/11O2byBbSjlLlDbzvG1riD7c
ZWwF6q7f2jVLzIG8Lm5Z7etqdlhKxzf6XfWA3YIlY1Sb2i/5WrebkjJU3Z87KkOp
8yADVQQA2/KjnS6YUBFgn0O11Kleh3P8uZ0lyXcNIQg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31136)
31UhTH470aH+etQZI23V0RDWOD970CQ8bXJl13JTK6PZXbHfoHy/kQpMWROg8fku
LO0p5BpJWuc7Pfi7iRLPo2tmAtACbBNcOt2NcTp1gB6K1Lxxacula+yQv4MNyLba
oJpQYfTsITZ2vBEOa7x99DJY3v7DEnjji7VD8EYlWMsaMX98Tu3FFtqkRSCRmf7V
GqBhnw96Y/fxFoNhnNphURAw5/suzUdoAQ8pE2fqrwrxiRtMHw1S6fl4WOIilaPz
OFcLztbdUWCH8dW7EufVrCeC9SzwXfpYIL55nOkvJSW4cDObK0SE3MAbaigzzTlr
KpkTXex7bvqay+xWnNWqPf7RPFlOsuCVEB8enBOQP1SmWumzROrWJIhCaLKXxyuJ
yYTMpNba/fiqRPu/qvuh2XHMtJyGn6YuFZ17TZ4ENcbprppvLkJqUdHQsvwCWzvw
EN8KEzXnqunXDrcrEVT02JcZywlItnm9TXqbZRhS9uPYbKIcZNAzEM67vvvn2ArK
fPPO2wAl9jqxtHGt65mSDAMdpLoENJiFIXIEcc1SXQm8nOGtbhP16ABPYzVATdQ1
28wHYtbu3q6C6rbZd7aJyKZSJPNYDjSf+0VRoSKbol42BHNR/wPaNDYpmj/xHrlV
Qei3bP637RM5QgKoCMp7O/0PxF0y4XxrMSQOIL17aei/VnSto+GK55PfGqG/qBEh
02wrItLoSEWxZE8jsLfQ9Eq3+1PCGFrcPcaaCSQ2iB7oomSkhbX/qk6GPPUaMYZA
zAqKRDUBg7plJyrxlth6Uy3D5Z1HytVvWcyRtkRfE6zc8o422pz6y8Zz+vcRKsrR
BfMYQ/QYSvPadhZTC06kbWN3UfF/lh/cty3d5W2IlcUT15GKvlDypGxvy4EIpmi1
2HUVWqG60nY9dgXcRRycehONwCxFUKFtTdgPDHNdFU2/VbW5pN//P17oqH4Iq1pu
w5HE3cLCHMiU6lnOtmUsXWPtnyCAFuVrUXv87yjB/q46XkbsG9cceeDchm2xRQbX
C3qfxhYvupOA3oY4a7aBSUrGL+DqiBacCmkODZIvfU1SI9sbhjpIXdPlqlV5/JE/
8VjraSPzKExBYpEE4a890GMkvCnAxo25yqjjiGgQfuYxA05vnzRY5hhOFImMlfqp
F++vCJwVx7be4p192J2ieHxc9tcFs1wSekKcc2FROHd1b+XXXatiOZ0tIqNWAaRx
t/O+FOQOVL5QFEdenurFAPanmP2m8zK4sC2jxqUC/9/AnDMIbaaPoP9oc6bDOL3j
3Oatk0HYJQ2qjXlKrQxeqFRGeRWNUmBIY8AnUryjtJb+uiJWLVVOs02dV0/0U4WQ
hMjGrChP1ra1KGxJWPZT6cAIaNXdsq5AeRatMokKyuB8dAH1FNPjhAKkGgEWNAtA
7EUdJWx3yX1D5dOU6aDpgZOvmzSAdKRFcJp4BZYiZxUn/gE0Xhz9c7ZbFdnlQuol
oXk8Dn0I5EqSB/NVP0z+zNN6ijE+11m3CbqC1K20UZwhdQBX/OHAMzgaXdUaGHvH
inQwlMoAXCz3Ah5KwrprfiTGBOQsbmexJrKcgdYurNBFiLw964KxlRtu2+8jWcTm
k8SMW9cHDnUJkZ73WHJPZMTfCKZMfWMtARVBM0POIFOxHVnzMVmT9TWhhXtMCbJB
1ndVswqpmwLuCnBxM3M6HW76EzWCelOdiyflRcYiAge2hKoAhqMIPe7IW4eyR2xX
bxYi4kT2B7HB0UwUEH8Z8kFpeerWO7ReOjaOqmxLW5p121F8tMbOljm3OVafscLz
lJKmS/AtmqkMxyhi3fuxJI6KIjId5VrvX0S18Orn3Wi2CMpFTkECvKyBSyEiqZX5
rRgG81qxhy9xXMFIb2YMfyG7Z/HYCFMOgbU1Z7D2T10sYKPCMBOsFPPCsANsgajT
0kaea9YCtPMvGeA4KVWZJJLuikBGqr6QkVSKUcwepirBgpZZo30ruv6tLGPaJXLs
egZYiTb0ENpNIvcuu5IEST+fjfO3QKlVhFsEywFIgrcLFOnSA6IiowJbf+Gkorub
CtC3CBB7DSk9gngZO3B8llOsGt/vr9wAe5HSrREITC9rxU5XBb0lTFPBG7/7plQS
SFy+hpE3qszrq4zX2ab3VAHRn2eMJ4roHlUyVuJHCsKokxiV9kQ/ITk082cVOC3b
v6K1EpXlYLMbPEn91j95rL+IbmQNmUzeVpG48IGLI5q3NGMkLkE29OOxMbPNQB3w
bPuhxNU7hZiFTQvi7UBAxdky+cY78uQsmo3nZqyy/WLfRkOjE/GAy50UpnFc68Zm
tzBMAjtPgiYZ9UvuBmvrEXrLjScqrbD9DyN76l5aXdjK8gdP5z0r0CjTpmRsYnSM
DOAaMBP9zhSo3QhmgpJiupLYrxD3fIq4Bmsei2WtAqaiT3Rne0pDwKPjtfgoKLUz
DojBK2XQu1ywu9bhME++LJv88X3x/cPosFh4Q92lDnIg8KmT/h2/DcLNwoum2SPL
uW7HS3tUUBNVDKnhNpMY0T2joZ380xWnsYoQdZe4jrSUpADqfeJtTVOxVX7ANkEu
SVgPJoQgjyNZf6KRCvbaBVAV6JaEw3iX17pN3fOPBoWLwvE9A21n8HC50gXtFoaa
gcYOioauOEpGhWwUPJyQ6vryXQR/H1U7C9epFb3Qi6W9eFV02THHhn1DZ1GasCDk
mBM9PsJNlHvaNLM1PykmInV1FBwyGAhmW2V4372Jff2TDmuGafrxOuhiis8GO0qO
NY30/1lWHKgOC4yq/zuZV5FgjU6ZN4QwKJ2Wj3k1kyTAetjKez1EJDR5LNhQSPsB
vwcfcO/hKTD4w6xClvNyQU9KDzln7ZBN2nUnZSMJ8EzKU7STjGYL/9PInxRPKY9f
clYhp+RQeC9p9RwUO+W74pkpFQyc1Onq1eue9JTTqZRjv4zd8iUjXyMcNx1a96/N
iiDgNtZJvfJM5iHfZLWQmxPPaWqYYdVX1Kp4X0zYQOVsn9FQ2+Ene/YeUzUzGY13
3xituFmAcSz+P2WFfsG2fBG9N21U38WKlwi23cYhPaNmrN3A3Q5tZnEyLnxxBRAn
voUtmsuy8xEypxxytmUCpUaf8KqdooX5O/5zOSTwjooXWkmyDLoPjjWl84h+9Dv3
HlcShDU+GCps01TjzjcLAiLjaOx9Vcem72stzSnp4S383KG/ryTVYUiN9fSiUFvP
djJNhjCMJEr3wJYFywy3H1RTh5yvPHT1YqPxKr6gLf+Kwah6TUEXLPTpHzvk+RIV
GMOCPiB0zRm4fYqVrsR4yeApIOv7VIkLs2peKR2aAaa+FHuNfjvfm+MDl57oUlMa
gBv8g6s8xxsX2H8g+n/lOspJS004g7lNvSSCWbUrAMwscO+SrbyKFCC0jojqjl2t
UhkM1gVwMvsBADjU57lLB8F7qE1WVdpiRwZw6cAMjsL+lhvgZCtEfsgQzLe8Z5bt
o/eH0SdlZlcyIUgfGTUQQ+AuIHFGSG9NIvdpmx+41mMrKCdg2LDe69ryHCtps/BC
cGEN7Rvrce0W7dxaq8OFtbg9R/izP11Za2ASzC19mEck9HiCT2Bvfo1W/TccJiXP
x26a4Vi1Gm6dCShPqigD2HTWeZjTElcQ1Li1dsRdehm4F4+Tkrbg7VLq34DRMcTr
xJJZDCy5sMpk6hCyjRQ2OLVSHK8ebpsbbqGCxfWwZhUOVtdG/T8Ya3xLjqoIpn+P
D7if8d9+rdEOxa3p7hHU6PiIzQI8IhAXUGzlzpJkWI/PLIK9NqhrGHgeauCqImX7
0q9roVT7HPL7hBCFDL7qdXVGnnxR6UNsK2qdU1MhrrBkaxXZC4vNHP1ameJxw+4a
wDeDY109pkhNbjrsIoNWqOpgM5fJKTX+QWmXFl8dXawqOHvZWWWr6noUVGU+zIuC
dy5TVZuuptMRQ3bWKNPtfFLk+EEMa/XCkFkNpGO5Xcs1eS4kMCXwHydva9M4pExC
sV7h8np//JtB5413k3AioL4fo5GFjlR1cU0F3y/dK7lgfX0ACW16wC9OHaoQc2Wq
W0QpaOfYSpmXYb2hbCuYJiiS64I+JTpfr4R7Me6QxAbbNAowzvuJ9ASfmD6/+iXF
Ap+Js0QTIi96sDkjIUpFq7AUBZgScuK0OuSD8Y8HQQeqLkjM+OYmdJRysQJRZlQs
2oCC8A6yJxSgmcrW3iajvJbDumonmqFZPg8/ykKKwvl1MFkFk5Opymj/lLjVyhgt
BO19mmJspvaGtpJ8OLgD7VVViO9/AFGp7FTqhuWY5uZhgPGuC/so4YAICs0vrjcl
GscL42MpZ/xkIEePd3cV0uA0MqOrQSlvGShbxIIVt4Oy5jlyZnUDbHXhSm8KLW89
VQVqGtHDzAKAqM+XRuyZKHkPrj0AHvgKDbppjxq0K6GvJcgTk7NNvCbpXq6j9GMx
vUgiWLfrpG2Okw3wFrA9mCpJWKOhoXMKWmXb4rlKpmnNZxie6bJVUqzdWVqcMVtX
LNuhF2t6c7XWLYMQB87AV7JndogHpBcVfj6NTwAU6fbPD+RbSTkEZCo0EWAmDREL
ejfjgfUT/L6vShpADwEEOtNJMxRqnZGTRdqVkrfIlZjIm2O1p6BjKvgwx2wNce4V
+lizbzluuCPm3C1eMnbjAjAYr6IvMnMbIsSqtLq2F1gr0EqrsEjZS0JH81+oUErH
VGkTgSWxd/m8guvQwrk8HhzoEJclk+2gUlw2d9OhBhSdIsECW0iSa2kW32ReM4IE
SG1JJUIgoos0MEDLpQY+iSs/yGbkicp+H1w4Xg9Bv9qW1S/OYDIosPOthpSGwxNB
/dubRbTk/fklEo2TIvy9qoLMQBKIbX1BXKJX7CQYBDIkW2faOBNyszGJwDJARtOX
n49IDn5/uThr3cS++/3BrTlkHaQfT+ViFAzah/CsPk3M/1VEJ0HalmWkHAnXmLVd
JgM80FVcS4NP1KynRBxCD3MMqZANTqr53i+qzurXQ1eq3FJ9nV00Mp9/y8jTO3e6
jYVGuBKG8/wE+OPjUfbPo8FUTHfSIAOCaMtJuSXdK0S5rJ0qacrsD/zue5DFSTQG
JgPPZZ8LAjjbKYoARWBtczdVFO5lHwfGjaG7yJREphvJgXDoNkNgovi/g/ht+Y8N
lozwmZJfJRL3MQzJ5d/yhtO9OhF9gblThUH9rh7s6uiv/ytiUvUBifrOOZsiCnac
WLlORmFAkrMmlGOQ37wG5iIbwOF6qcKqG2/svur37rn5jf1xeeUQ8SWrhXiw9kUp
S8GS6Elmp0rO0NmsiiOmjvY43oOtYMmkzMs2Tv7Gftg2F37I3Qb6xlN2gBr9btki
W9S+CnHnwLLLS149q2ILKOdiDlbC4mn6pN2gZ4bKDoTddS1f5a4J3wSOmBKothYe
jtjdw4w5Hk76K7GI7mJtOVyR00kDlr1p0yAH90exEuNVtz+d9lcB73SNUKVDDUyl
iqc61IcXQu536lTUqrSDETJJsb2LsL80MzZvGehkY+u5VKWp/RECu45gbOAoWQSK
uTZUCkLJe/SZgvpCUGRxp5gSigMhQbEXYkCIn3lwCj6Gm6ApJCvzz0/t3v2TU1t0
aheXEoWVMQscJkMGVMoG+J4griKUDi5thTjYdmeVezeqPcX6uE9JU1NDZoeLKw47
iEF0a4+jciRkQLItqOxSwhc+OxJUuN9KakTX2I9ipaiHnwCIF7GXbVMQzSX/KhxN
qLIEfCIzm9lL1aavFv4RdANtDTNMUS/99l/uctWsmIdzzpMjs9kAXuvKzSnSmvIq
udlgYaAYm+TzbfENf2ulAzXCUPItnfsFSssfUo2myVZeFgzks+xaFFsQmExvNfjY
EvlCcrC4luxt8DPm+CPIKYhuSgmMK2mMSqksJlY7hoqqkaRHTVje4GyJQeoDjd5H
ZYUPTTSGYGpKVfnwUGQ5Bzp18BxImGoq87JwjUcbjTRK9PkJhB/WxjPbCE+IOh9J
Ia957RemOo6WDqLzUsBCUA7VwvZh3/VqFleoK7kkxUsxCQIaTdGAtcDLpY87yEq+
3m/XZ5V9cOZHfNmaovmdLaSIWJUJWj0iKK6pSskYdYJDHns0Rcw2tWd/REstZVQ3
iXlVR7AxuMmy0TOczZ0TDpoq/fJ1ff1FkiDsoln4QhydIvnWF0siySfd7R/kZE+P
I1UzfaI7VaFYeAsjGllnO4QjD2lDwlCjt8X+cMso8GGzfCufA537WtvmuwHaENBe
H0/Ro3PAyh0aBS3vfuXv0JEoA2LPpN9u3HwHpKZHfQPmFBZaBh3CHmt6wZI2aL3T
2p2ro9BOz9Vdk61qEXnnmQEfH3JNw1Ni81Rrrc7570HhufZetWbp5zHMXrFYWWOv
k4nAcpV344kCrvk3unIur9NoYHmsOOAW6q28S3QcIWT9f36zVRwGdWoeX1/EOreN
YwVz0vKEaPd+c1J8/ZCzvUBdnJOzp7StHDFoJNMMvOtQS7oz3czYPVQriA0gp7MT
f3DZCwBKlpS+sq7DbzN7ufcK7jPajqYZzKGasduMj9RUuY1HFPURohb1zyN+28/f
+HQeg/VV1wArlcSVc/frqhX3zeC1sVsfUR2Zuhu7TOYuY9nKFMbKW8nwQkK3qqOw
4ciUjr/xgEmtcU8f67u8IO6P8I+mf//f0v2vfUZpKjehdvb5lz0CbuYrX5z+oZ9c
p+728vTchN8gCFu2PS+nstBYPweYZO+dW8ISbsNn1vEKDupqe/BSHvM2Es2zFjgd
/Dp8EDXFtoWdJxFOjE3yAQcttktdDLB5o6uUgXMorUXPTPloW6/T0FLjiVk8ZxoH
gZZ9/KRCs/fFRaE02mxjp7WH6q2NUMfiutz97cSCKrbZITJJdGiUyVE5rQs5Qsek
5zFP4gnFY6gDtqa6GeP06hHXRjWgFq6BlqblTvXDB6imLtHNXBjndY/nvG0/uYGR
MKDbvoUKyNFstnSObdpqkGB+dt2G0seQvreljDvYzp7Pnqovf3r7FdpvmpbbUjsa
rReHBOuaC8zWSw7A//8cT21e8nfEOFOVIh5rM8YBtoXuZY4IRJxC2KMZe8ldyeUS
MmKYSmnDk7sxn64QEf1DfJlARkMxrBXuY8kKX+23UY60IssLaQp1F9PluoI58/FJ
L+J8EIQNCIN2bIBtcLvnyiWSPLCp/f//qPGThtOfy60YkLFuaWslPvQSvXHJg6lf
riursMvjS6N068hgxiWALzP8YqPL70IMud5WbNLRNeSGlXAQ2aDVKdb1B3gqc31N
f0/rqrF53wjC1Qo6A4MFzW3CNsddeiOqkVgTUOixsAfgnDLol0u4fDF+PAHMGZMn
1XyTpy2i7Hx5/+DMJB4nFeRa/TLl5zqZwKOg4UqFZhWv08u5PvLfZngpurw1tIMW
8ojRmIu4otM3EH4vAKycDIWvJJxG0krw2gKghPLbrD5K6u+0fzx/Igw84t6tIwTw
qRuI6ht4n3+F/DlqnvwqpLTsUxmfbSBB+nT8vl7Q7e+ogDPxfPvedK5zkntyP2e7
HOuiFbEJmhIBes1yFCy5MOqs+VCRL3wGpWG7TWLPMC0W03YLeh29/+JEW2optsUz
RBf4KwFRI8IbsnWoRQ5Ef3oGvHGLqOVJOm+aiXWYoVyA0PHja42MHOX1yRNoqbHr
3W83/OFRY0oQKpoP5UyBrXnGB4z40brTwNj5tXdA3LtmYsm9ZjtbhfXV01yfSAvz
OtV6k1KMLOTfuxNA26C6XkqY/WMsuCsDqvXZ1RU4y8mTxGaNSYVAg7hle+XNU45Q
etHYTmuC8+u98UXM0CVTTIoi6V5OUrudrMYW1jxPacblcDgI0B/MlJscd8N7WJ7J
nLuq1j7M93VUrKGnUpTFY1WmDmzOs5yRzulsN/G8X0bi2sJcLsaiHoBrsicAOhVR
3H6lWBxrKkQe4WPazyQStUGrkLTe9+CJvUtlfeZP5TMajlcZ+Ylb+m5S7TeYqQjp
OXoxk19WPMmZKMY6IMH6XxBUt2/DYDwLl9E8FS5/vI0GozY3Pl3M7TdTYqSBrMvB
sYNVtozCNz354V3NVVyDp/a6daLDu6XO+YTcqMatXCXIxB580DAVEP8/L1wM4u3v
0G6YQQw8GrFNIIvddg2T9z54DwlqfZFAGQczK+ar0rOf+7UNX2ybym97wgwss03s
WSYMr0sf+CFCPNPuVfpQBDKrOxgdLriK5guk2oRuvzUYnyKZ6iCdO6ntj0a728UK
yiU945r6PmLEfQQGfYovCxpG4CZsosSi2ZWm9P1Wbi5fFV1QCqEPNfhbF8gNaqsO
15x+adGmKXyIYkY5gQmW3f24okUA/+tJPiIYw8eyqJYxOVISssy6U3H2N9rjLOTe
yL1AbpCV/BZygQFBt9DRi5yNBBxQUsincjPvYvjL4YBi2nxC0JV9/j+0pCPCt+M4
OMP2zahv9EgjldkUURRifT2sA964Kf7WGxLtXUyvIslMpKJdakwUt5arEQ+5meNz
9GUWEzTROvn9pSjjhJTCxYQctU2+6YhRxnKh/w5svfCbd3WucSqJZuyTe8imbbdU
Fj697ww+nA/bq6UAOv5l10g+VgYkjwep3Fw7yyaSMikshto80RtEguM6TM+HAQUj
UnyawlCAscqdWmwU7E2rFGYGu4SrDq38GjIdL+saNim274/i+tYxc9s9BR/cBmab
JPhKSxD4uagkCSSlo8AEyJHE15E6k11Kc6wz9FslqO2GhUQssw2/Wc2Y6+vPL6Dn
adYnwmFzIj0LBYVzb7i2HKTqwVJt/dOuB3FmEfMIyt+WXJBdS3mUxXdvi6PnvH1J
GPfvHfNnSfecLntPcM+whDbttp/IeQQW1MWgKaOwEn1pDw7fkIbi876NCmqPVST9
2qREqLUo3Gz+5Z0+doPfLivebZKZK00+YvGNrS1oXGG6vltUgJhOz4AypSW97MnA
6KCizG0KJ/5Kt4NfUK/dGux1eXDZTxj/nQOCtpBZom88HUwvpvC8cSNPFOTOX4aF
rvizZXEJtK4CrVkGaY3yAvuFbEoC5u0scsVtYRbRLIBlIFWn0nr3VZjEOgB6p5e7
P58OaJtPVUVBmuC984ORqqYcZzRe+rx+C2UZSTHHMwBybNqqb2cJ6+XSizu9OgfI
X7QCg6EkQxui6bptZQVwrq9+WNGj6NStaa52i/NETgazYJZREsSJRKi7SMcpvkhG
sbvIPxpd2hppoSzJhBzXuPBaEzEeIK0sN3gi/U41m3z0ir28XsN9JCbsUBtqwko3
+8QiyZUka+YkOoFrPX9iikjUUETw5lcNGRGPf2AULwsE472G1od0rWXMpeh3de2o
dfRoFaoe8wTCodz09hKMLsHOGX6i9lTzG0+kcwp373a0fijO3OykT4e9hOkguI99
ta33M5LCJWN6LwzQoLd+LdSuI9hquqbzUwskoaRgQ3gc/MNRhe83lcOycZ7EHTjL
fVDTZIsoqXkF3A0nw4LSQN/jni+eXqR6KW6HS424t9c8NHQYRdH8XE1Y67iCFmya
uQpHlgirVWnnn0wpOjInx6axuqsYwdeiXQtq+et4XDNpBH/HWSlLQP69f9m7tGBu
324PWE9E5Z5nrqu/fSKmbDrJpmRKOUyN/1t4HBjdE5IF+0J6Ph7wHrGigM1oT4in
Ny2bwdGQK/wwX/afSP2yDXwZ4ja2BbX4VOtuxm7WYFwBuXTJoYqXOFIilvyldwYt
e+3EvXgIMySppttOOYYfnqll/Vl0v1haGI4ZYvnBNwypDG0Cnh/CmbUDs8K//G2A
g2SKd6fIeObNrTtt3TStC7pdEqsRs+DPkC/KWrRWu7whPpmFJUrlbQxmv3EVdmkT
2tKRYh7WOKTTK4tFUAUk5JchxexUZzrsdlX/31aFXIskdlWtn0xoxUFwDGJuB3/y
2m9usffnfP8RYka8dLCUF0RsoHYhC2VeWZHpWPK++8GOEKreZGeIo6FEmbYQMmNJ
jv2eoG5eEF4jwIs+3iDq2Lzg1K+nyIhjymo9Nlby5fkgQarcAvISljN2bNnlk0VU
2mL54Tow+fmJC6sPIYpqVzTkKTQJZr9KHNVgsDdUTxN6R1IxajscK0gTBiQWBdfh
1q6b5HImrhiT9LiQ4kHzXW+7cPidMGorsrn7rEfPSd/4HfTq7H4PNgBI9KMKczl/
V8tRbwX/BHi+nLNG6Kwykfay6B9PjtVeHqKnxxD15qjlfHv9bp+h1Mdpw4mr8v93
m8lOmxXSqFid8WXWD/2snzywHhqWRGM8q83fblm821djR1M7h1/pG3b34Ts6NJ9e
In7QOmaErnRKqq/UK3T45hA0nuO6/DcdcfrllNfMZKKWOhruGUiIeYm5dfmGy5uq
oL737aTxcYAJgRibq+K1UdGvUo0WhWdOejI5zjiw6jLn0Udfiati+Q9TuNYVgMIv
BjCbtQ9XFLEjsnOaJSHgPfPUVc+gaQV7mH034zGxWajbr6Ntol8rs9L4YYXLg3St
5KlY/nV4TiercaxPEwbRxBqbzcbVJlePbup8Qwv/li7wg7bvH15PDd9wcrJlQa4w
gIedu1F5pDAh8yMCS51rVN6TWpK5dJXjDw6XEYGYawyTri48HUGwzhsr1PD5nHJY
RKrashPnooZSIHrNtOVN8E8swQ8wlueV10owKruCpeXVBB0QCB6I3UFLWhBTRvSK
8m7BYzf6AaCUAFBArlgD8mfJ0jd9rseo3baJviH4+B3SaRggvnsw6Ad9/DqIEsr9
n7df+JqYyl2Wfbr6A0l0n6hjuH/HiIw4FUw5KEdrlf9Nrh/gK1ebSKAvxx+a/nqM
6tiTIagaxylI013zTsJNYGbKLVEi4d3xg5++ViOjaNpvJesuHzxKPVwA8GjudZhE
eyAJaluHaFxWAkPUWUmH2d4BDQdGfRpf26X+eWAWcJ0y12eNs5bLsjaSX+eycBJA
342fLRSbn3dCvG/KxpUpwnJ5wQHjI+3iBt5/zOXx66qotcSqFcVsjqAIKqksDI03
E6r1uCE5JCWIw+4QTrQnqnhXzCsV7RU+umy/aaOtJ2xxi0hyr6pbdSDQ9Lke3bsS
5t0x2g9/zHvjpRh5lUkQnx4bT1M0Dyu9AbaqAZiSdl+7t0UwEgdpGxvKPXcuV4Dz
CJSpUD+XhSZ6BRtOeY0y5/hjaLIhs12zf/doleLSMJv6VWUGfO3zf7/rynXaKWJx
KdqjI9NCN/zgbp0ZAHUJP8ENxwZTHI3swuxm5W+TK5md+qOu+8HgB77LqCAsNECY
9kaFy6B7fV4GT7Vr48193gCerT/FrOcQ/7urrmmK/mw78OVHEZ4d6t2tLTn/fSIm
oAH/ymacpcdC2HyC+xQyIMyKuJSiIizPF2b5vFaflnOVQPrICfYGcLaS0i/U91hM
5YCIe/sSvEX3lqql5lN+fA+ckso3kZ91/5w7HKEIFB0gTDB5wRmTBKn5jgLbt1OZ
krFUaVu0ncQk5k/gOw/UhVsxf7Gtx4ikewnDwaooFVCYC0d1DPXahCN4D7/kahA0
3KHQ2yI148op2TUs8ZhqoL06B9iFVr+SmPpCgwAwpx6yob2UrhTPzZVGLI8H66QC
hh3C/pwvc/ht7DNB4oH49naQrocXEEC+2dUPqFZtFtnWtQCsc0DD2dinxvS3f8gJ
MLLLE9IS9a8NgZIz4hfnu/rQEzs4zbbKG7j9wMgrICLH856+jnLzPtZpUQcdzo4/
E3O3W/nEHFTMzZitpBhdISPqArx+LZAcS2q8MHLuyQTubH24yLDbJIa6hzdI8Ubs
OMRn5oP/qHOqrWwYkWCeT65AG9XjlSU9/XFcPJWqrPvxRos2bHBoquw1xA5ZtUaF
pZ1VNlnHum+DW+Iv4bKBXCJyWP86i3rkgR11iblgYG3U89CTpNNAxyJ1qks161qm
s040rortAODkeM+FxLnhptyCRYY/z5/VNQXg09qPJx7FJIfV73hfQKV12ld0IZdt
/67shG+cTqdh8Go31TpeX1shbjDWIyjFUStu2r+2JkRAlBt26IJGmDZOwmw5CjoB
jhbLlVhWm8zsr+ZQqrmnMyX7Crl7N621V6ldZcoWBBRAQJUGxh7GpGF66j3fwd3D
jCDNwOcvm5rZ/T0NQ+HGsNmHyxMOG0l2XXcFKddB7k+Jukia2fx0R5c1QuukZP2f
Iy0YqGl25+MRezaoO/3UucV3jPcWPelzM5htbwYAJzeoK+oYxlMHTEO5b7netQEf
TkRBrdl9Uo5l7QZYwQZNgrA5IYQ4CJuZ4l1c3N8OxgQxp5DdjnOeBay1ai82Jh9T
wq4oZLzDMZ2iJgo+1CPXHBOsMX8A/nn6N/TK7gWFLAxi5UmKHpFEcz53sM/CczG3
mtkk1uWO0laGdE0sYhtjhiVQVDPWJaTNhl3N+dKdIVrVujCe/OT1OtfizQqiwS23
KERla7tdHHwqmDtP1BV4psv6e1ek6TP4bQ7Jf/A2VTZKaAOn9hVYBBzI159Fq4Pf
bbQBgpSPBWZMwrp7ulyhQHlw7bdr7Y/dpMROIE/VJREWlj87Hlfn5ahyp7zAFh57
Q6efwEksi3yUBF2h5+mbYEkMUKiD6+GDATsQd/92HbfMFAZmbjkZIbJeHWDynBkV
TSh3gbbNQZ8G5rFeSF0m+vfGSnefFoYdhxZyzlXiPnTSzWXyh9BoW38Gtv4rZHJP
e4ni0QRtDtmXcaxv1xNQSVX+x7m9w751IAsHHYgQcnmQjT1N1oD+iZR8B3Vi1rJS
mgMFU2AQa/l/RhN+bpWzXF/h55e7z42ULHKfL47Twx9aBg7m6gusD9deJO5nWb6g
/Uc7qhq7AG5CO5IxhfpdPJTGPVlT/Gx/BhdjgCF2ghABqbJ1vS2tY+E/D9zFZECR
OXXBdEi5lrnKuJ4Xo0d3+gvGqIc2vIMS7dkxH8OaBxsfaL2f7iDgvof1qNw9xZhe
V1nNSMGXxek0Q/LS835Dkq8c0a+U9WnnoB1ZZ0C6zPfqHKO7uGGdtlpuJimS6SL/
qerotn6dvqQNDa7Q3dlEBESFBitcLjteumwf/TFP+x4GSr6kKJV/zZThfCivmRUM
bxQDE2dZ9nsq9UQ9WrActkq3Dt0esLUBf859eaOWj8LVDKfX1O3U2/MkN2x8WwZe
3IeSAJeWn9WNYyz5P2QonPxqKJNIePXyJolpLT8ZE8+BMZabhfVvcrsrVQPijfGr
7RkMti4Qgfyji0taW3gDo4LmK6agvwP/G3+aBqlS4yzf58roDmUEtGhmpzwCrVzI
Zc30SIz7aYT1aixkqlfJjXkO9WUKOhu0VsGmeyTnRgAt5NytasxGBgBJ45pkte2C
G5GvNQkVBaNbdqL+qJ03gKn+FgrezT63ZKbZhutwOBwn/d9pv0Oz8+RYtLe9OMzz
lxyWg3fPkCPOJ9YPu66OWSbaQaiPlNBA/Ks+VslZfjrvbuQRFvd0VA2d0X89dmN3
ErQ/jVhI7Iez2hAwAePTuGvDz8flRNrR/ggnSJzeaF0D/1THS6XIJH1+c1WXemdF
hbPmyUgWlmvlBP9ZXADHxdK3J76rYur9OUofgS0Q0PBaYlVS5bXzuox7g1JTnGHO
6lLSCg4+0CyxK/l5fETfA9U9ACwd44guNvpbSL0GP57FniYAy2uQIP59jo26ROVv
Afw70FhukYuIoCFBTyYxnn6HWOT+Nfr2HQJyH9U7cUvfSRpsUUdMNj+26XNHDu2E
u4gNigERiYIIMB805Ao92Vzg+QGXJ0MlZIuCSMAsSjnsz05DZUSpSfqme8rvvVGc
ADsJ87mXeS2vMPbGJQnmmeTe05E3eXASPccbHYzANU8NmnXx584jF+rchuM5mKyf
NyH3dGbLQvxooAdp9C+DjkxYgOhoNYn3o++9FAOzevCQSTxtE0hZRUjlY8VLovZQ
6dQRr1Cp0OSjrKsgqb4B0cUPzpOKRgi96s6EMcpupBTJk62Em0sJx1s6ZbdkQOKs
Rsp23Lj1QdF7eXqWsm5Go00J2+gYxswZpT8I1lnlrL/8ip1jk4qSquQ9AgRtq1OI
dwTfg7e1lvp56w86GV7E4tkZs3VwQYKkwD+i5cvaZRaUZshpJ0DVFgnVTuFCz61A
pz4H+6ayiBZt1gPUVfyi3R87Dvbk1S8jHxH0O8LBo12y3C2xrthzaEW8t2VlIhoE
rF5tVsY6g+laHGq7FgMa+w3D5bnernLUakEBTg9k8qxDx7oMPdf9my/e848fhLFw
EnpBZaqpfP1uoojw9lmQOcNjK1vFjM9xy58mB8aw3Bfre5eMnrbatPe15iZjFZC4
tOG5JZCGWCEUuQk+NrGdUQbs6BjMY2KDIKloiHquezPk5CY5Z6ifeUJVkIf2dcmM
873h/QSByBxKdXzM62ykWHZ1/yEuTIqJaN6SPGW77REzrEk7DxTvyBR6CBZaieJC
/RdcxYn2A2DhjPRRenzcDaLMAaHg6OESxX3L4KP2OHahLQODGysdj2W7yAlwMi3s
W/k5bkNTok6MaeOp3lsVErrpTDAdLGB+ojvwytRXMJ5kYAVFkH6StBA8aEP+mkNJ
foWDZ8o08jdbojisgwWtt6IH2JIbihOkSeeL3A2uSDs6yRUnPYuhs5xtoKCanrIo
UzAW+j4zIPYZrhE1Ar/d5hQToBhaz4z+yK+M23prYWctvLyJoPHc145/EuwvUPuc
OAnEX/lZip8tg9QDlmGJYKJn11Wl8MnjWDN9f6B/RTcTT+2l8HpOjIiYroAm5e0G
JGUlowDOTO+mfa/fiG8cCM3+K1bYE4ACRSfcGbBLC1V580xykuovv6bwfIWUdDKs
mPuXfztvht2I51v98FXs0PanYsFWXvlTxmMiirjXvHvM601F2U5WiPj6/7kDw4JU
C6qJkYysbjdrRK+ZJgrkHO6uBNxlziEBsRJ/wRSAfb9sSN94OhXF3dX1o1NGhKyg
kieYWK5CwtfNy8PMJnY5iPrlldYJz4C8WHpcBvcC530M02kbd1LZDbm9HApvO29+
Hj8p99YUUP5Hp/2AEOisDxxYu1HJ9TA0+owAPIxqFpFIC2VIIvXHxzmfiDZlRLkX
73Fu0A6b24sFcDn2fJrSR5nzyHtzp7r0+2lZrOJ6GnuS7lMRyER+ZHSEaKKJp4uU
a3aqegR+mc3S/thPhDifRqtx+n94bRIfypVhEltyjN6dCuS3nyVDgLKaCqzKzJ6p
8XTtwqPOb0hs+q2WnAc/d7eU1Kk26s8J2BNdn6dBByFpDaI7dFmjKNoUwQLeFh3c
UsLwrwByIyI3MQKq14d1KcXX/2yOEhUVObRPCDaKMmX2Q1IVxONvy7pESrABhaHK
N4bVzKYOI5LK9F2g1SHthPVAQfXuNeJ/0SlS0lY5mq6jAxqaiCdcdIkMxTbA6Dyh
itM8tmpy1WQjASX38z8WLVdVEaWAtmCJ4gDFEuTp31ecvwaa9XidRKHjLclm1Q4A
X+k6JPNt5anlsKAB/ATZwaU6C+WeUT/zV5TTxYDmTb48g8aO8LHDYxohI9OfI1gY
+clYpSzL1vIw6vpLY3vZIqk6T/vFV1Ez5bFytJ3r9QZ3P6zu1DazBV81FuF06EO/
VJaWl0/RDajyIAAWMQWBNDuPhHobyX62sIqkdtoYY0K+TbBqUzLuxt0vLMRpQkMK
U8ypRsDwVicKoCfZU/GjEHFsVAMTkiJNoi9yyrWvrIcKcuG2Q7qqjJSj3lOuR+aX
8m9ONLwixxnSf8gtXgx/j5K6oe/Q6IPdgjfS99G53/8UeykxoerpWiV60DxVG5iz
wtoKFdBAV/XUZwJbsOCFVCs2cX8tHgDWUThT0fDf5wmkS9xWIvlrFQ5WS9B8Ufhw
+m1ZXwaDA9ravFfU7e92MtUUfdFqzEF6SE6bvWcrj7W+sObbY6OtS543xDn447M8
kvZxYrINcH5EPdxHMNlNGHVlQoINpBI4We+gcu28g1FwGFD7JCxAusZjMCcpq4BB
GVF5T4yyu9B9SKffLdDg2z+OgF5ehv+RLE56fTLdH9LPt1VJ17BShrEbgsdurREt
IHGZRQEmIUVbsW2Ra/qAUraYFstdP6jz2QDYor8nJDgZOiDmoHE2IJaMbTuynGL4
otAN1dXbGYJB/7RyRKYg86PHTEgtnME17f0ao8I5QYWehSjYBHHOCmjrARtG4iAI
nWPscznaW0lreTMbdASI7qdpgs1gPAtSUfqquPkx/stewu2Ck2HaRL3tXPO6O9gl
QEDX2CiF5AO9xdsEPhuc2/0293TrYuAgqGnJpyPZFrsQAM6KpnPThDdGKxPjBgRx
aXnjCbayJ/z1qZd9NE/HKNKR8YZIhgGrGmGXEwaNSUFvlOjwSf8IdwZct5i8XwVR
VWvQ7I8FefguWBJVDtKfvly7ygIfrbFZsFPbz/FGnM9rHwhmGVvaYMPpR98dImTI
2GL9FqJJA0jzCsyc/YBAC1v2oce8JurNnJXrUIAxbyY+g7Z1KSwA9tliFRb3ctI2
qEOzGsII50UHX7UWD/P/Ab5M/RJj5K4C2G//nIGIKKO/nTIK+Wi7h+SudydML8XC
kSfaVksWNkFrMiRrkgokV74gQ3F68JJn9rGzUuUegpMWGR+u8IfFEx6xffHPEUtL
bUTEIgANUJmHfFkE9amzffPjhBaoB1nTofzbUXB0MneYlT3Kg009O1XNIiC+sZvn
UrbD2VdyqOEln6O8qafvbJ0NhbCO2SsSQZioH15t46YdAhZMcyc9txITJ7RFBCpm
F9vSdYi/5ua2B83f0BdVfhCtH54KABgMDmVtMLY7Hi5UiFKBFDDUyBXnAAYOmml5
p8u9+X285wpnu1lfAwjiN5Zt0GE5DKkUc9vRINb8JYmg+HF1u/0RpIo6mSe7C/zL
reOLq8nCflebYzu7CClyJfi8wXUmSVs8h4Ej8fUs10oTfTqkoWVmus+afCOxd9wz
Nas18bUkOEwdIM+pJDDUklV2vlm4hoGcJVZ6HzOmbUGuKkrtyX97s7WozsTFRG8+
VY/em3ERsWBagV8J1e2lOQZIB6vkRYsDxFjixtqSRnw/uE56KhiB5pJfQ/G+BhjF
b6pwvj3WeBd2xJ+X/2YWAisak8MozcxaWznTMsE7LzJ1yF5NKmhQ+7jVA7baWefC
MVIHh+1njShZifgxQWGDc1aMS2t+eKXendu5PL+2ZK2yM7G4+xemMq8kh8wuR6b6
GJk+EehhFDXCOnMDQC5zZ+YjSIXzUZiBIyTKgnl16KK5pm0lFFVdjH+odqTPSKYz
94f5AReso8RL9FP66eORxAWSpagNb1OCXRDOb/goq6hUL/CV7b+d/YV8pNcLs0t/
wPcb9TnKVRR9xI35aTHpSVPPcWdUEU7FDYAD/n530jNcurxAgpHmOlkG6+Qnd3gn
ahZNWy1RQ4spTokM/U19AJjg13QyAPXPOEyM4DKZfgD88RXSpbGZ2lDihKeZC5j6
xxMy/HVINgDO8qxAWvMxWsp+EvR/BDJ5YmfrpTAG91X+HnbACRp2QQvwqOX/y09K
OzdLAjJWKo3p6q4zV5M5oZBnOTa2dFqKHbZooc4KjRyEuAUFTnAPp1GILVgPf6JD
3sUjd4MfWCOCYNPXbXLt5epFcPyJaJzC6khjNf0eq5mbNqDbiRSz5/3kHjZOXKxf
sOOWUZCrJ29YceBo0RL5Lhf+8+jMVGv8tGMxwATOe2py3v5VQ4iUPpWh6yo5xRBA
aS9jea4uuYX4oNGR68RYtWrwi9fcbOAYPeyHemJ55AU3PN7dvluq4zdCoqUcLhDS
UfhEtIs65uIPiqIl81KfJhYOw4W4mZjVMZNZtIUFOFni9auPx9Dnw8/31ePP/J9j
4XZtUb4ItWmVu4QImb2CH3/gkrsvC1n8e0zw7S6pKgab2DHIHNb3PCaJZCjKJj0L
8gqC+usq/9xcGcTXrcQ2mboHm+ruqL+hcZpoPoYPr4bS+8lOxFEln2Itae3XQf0C
Qjo3kSTGkfGhDfg/eOTGY37ieERS9iVY6Rri+kQdNTJ0RibD+eyeoc2YMrtScK2w
n05bNuGE/QQtSQGMfZ5lg9f3IvuPbePR1MVSSAo5GJzl4Tb55sfsz0DgXFwtxZYb
wx88P9aeU0BXjLhyj5KYVBFXTxIvFJFqFz1GhOSygZ4LG7S6Z5iRlLUok7Qq0Vzc
yG+baK7g7DKdiGyHvZl500KMkSoaV7jx3cOYO/juRwoBswZFGs/6uNEinEL3EHY6
TO4y7w2ecIEK/FRhzdHIUbSH+C24Z4q7PbOcCJu5kWda5oYUzDptZcLsDztJc0G9
j4UajZs0spRWPeZ/zfkHWeUqLOt24P+wc1ZsTcrna5Cr4rrGjLoZhot1IKS9AuTm
P6r4/Ev7V57OboieCMHFX6CFVNLcZlDIVw/bOKIK5e9MPRMWf6r9azJfzKpe8/63
eCrGL5qPdQH27Twf5l7x+OyfoqJteu16ClJJH7yekOEADVl/MYhMG0ef6yoHUiEi
dPziVWaMStJAX+MaToVTil/pb3JBxICaNyHa4DSbb4tSihMKMaw5pVMyyDrvOvKU
FHzWosggslicZx2YF7Hn1OMlKcToB6jlK0bYYkkCX+a66B2/CWDz1B4jx3X3bRie
xWQvMa3xX2Hj8Vn5tn+fdclBUTcGMkzOi6yk4qiUZRiCrtL98XMDv2jXpHvR6/H1
8bqOo97tQ+svSlH5RS3HKsidePPi0bCYkUNV065yQiGJOnsKbhnw07/5ZDiI+8IL
GL0l4XAL4pEZxg8B8OTerWkalIaeeUOzLm/zz/Axlc/YfTVa9lLaioj2secdkoHV
VWV5w84ju5v2ItmkPJgZQg7S+UoB/H5srk6JMlquKughWUFotoQ75Qdv1Nm5xwIf
fOkO2wMv5Xufd5NJPxSI4SJxvoDJDSkJXDUXK6IIL4DwZZlZQje75GIh93WkWs6z
sDZdcVq3Y9VYh+bveNcTiQLKTHABc3WnkrckCEffBPOuhq0JKp/w1ljuWRXYnGho
019DF0nFPsQ/I77ZLG0sqIScPsj9B6WpeL0yOc+YGoopOEkGmIzW/JaxXXHAATNG
8sNHBDQIyGWC4atM5UbhmNdNE7l9qoDupRyyvGJblIt9IKUrRIOpD5FFgyxxoy2Z
bRcGMZB4djtgUY1CTo8z9irShKMhRjhobA8KH7iIY7y7VtHkInnGCaD/+zoL/OQ5
PZjg11h8A6qXMiZliXjEaeyyYe6ahmxcTlcTqBem/bG2SB4cMiT7LCXAgJTbq72p
ISgdyVQYG/sJbZJaYu/oGvhuRw0O2gXd63UHeCSXfay6ADfK28JvKiMbGhKWjTtl
oBB/VqucCdRID6FGOBmddm6HgruGA3bcquVSskd96iBWJniDwcf9mb31zfI8YyqZ
o2snDfdTtqcFt8VEeaxZiAYheQbtsI5f7ULq3CitNS/+hClx3xOgm2yktTkMoH/+
ciI90nOgrEMJEuRiLpLGXDXkjQpL+VTSOVZd2uCVuGGLKGhAwI6PM49GxPbaV8AS
VH6UvXUwvSR14GhvzzBnhViHjUVBR9bHiD5Y9kNxqPq1bDgDDqx7IPxLAHttXyVN
opQG6RXJuU/r3HK5mJU2x3GlsJgDrQnOK27DLdHmnKrcL9kSnQAaeFa2eW8rQVQk
leZFdGoxkL1jSZ+8YhBUh32jbn98ytUdfmTfmAIarZKRbnbnVElgcYVrAvRGdP44
X6VspKbibJroa+ktmsFf2eW9PK8xcTKuL9DJgXgu8sjPTWdzjG/o54sMPFIJgJwi
ucKoz8egRSClvC4VlY3q9GsxeSeLPIL8bQO6xI7Qt0OAXScAWceroxVBo+FI5kW1
u1sxVYMGuWOa0WWZ7qTD8TOvtKrBRDrZYLJnnxvH/czsetMjipoiCLs9wDVQ1+SP
qed00e66DWp5mTxRh2/WdjWnKrtMy4p40a9BZfJV8HNKSRQVc3kUQmqoClImiHDf
4KWkufSQEFfEqb3x+KTrWyJn+YGyP0jVXJ8tpeKXLVf31w32Tf91hjkKPr5U4TxQ
KrBpfTdnksGcRZrdr71bqdlSOeLN1ykBwBK3skpZ0aG/aMck76i2yJ2MjTzG09CC
mJJVa/l+VsLVJQWB/l0m2rrrmX2qhtZaLn2pnzdT+leKzd4XqqH9MlLX6cIifrs7
NUbo4hbEQMFI16Diiqd+ZawjEnGnqyciwweRXSxPuXJT/NEw244nEDj3nYh/vwCd
PGjeZeP+yuKMYeGe/kfUpoQtgTacDW/Q4YLln74RHANrQhL5zQPSHOQzKkJ1ouoR
Kn6p6/qMunnQE1c/8TxM8QnkwR9zAN3A7tm5y00ClMvouCu9Wwza6ohXH/NKAcxZ
QgzZ3dnH1Pyz8sU/NM3V+NZ4sJ7PkUVHLmdpywIoQagKeshxhcUai+QIvXXNNu7y
JJGlPOL5fV6uDFBkfZZz4uLcHGC3iGKIvyKc4seVfd9At4vBzlfKYLrJ6+8Isuef
a510RZvTTAMQXx4MnCsjrF7q9adf+DDyURYpccMUGaQSb5VvfVXsL8tk4L22JDIB
GuDRAkB/cpGluYSD0wegY1KS7Zhv5TXsJXP+H+AFBXXXVbS7ChQHYIEpDIfH6DLr
MnT5RBXWCkxiLrH305c7J5kzE0KRfxtS6WPCOq3IHcAbv7vjsvWx8Dx/QLxrxCBW
7lgZ03UbaSDPqIoabSeWXNZNjPK3fvD99FuzNDmZJDdUgmzd5rF/SePRMqV0EY3B
yNkYaofl1lPD+smo5ZwsoijIN/DzTypJxR8EPJgQBm3QPDGc2YPX5UF8H71ZI5rV
uCKxMhIcoA6mNv2782AfPmSSB9RHDkmlPtzIgwQbtWQn5OGTssCZjaLVRaTCaXu7
qKmsIjIGQhNnJfRbLIpDIhG7Cl1xCgCFsoHENhxYeoRFiM+tuG7lROywwTELONz9
cRqf/Rgu9b0exx4PMiellIsCsRJTe0P4Zil+5ZJZ/qceGkf/jE0xGyby1iyp+fgJ
ywXoJbBcFqE7TLLx+7voYk+qk1EgyDNMFs9zbsgduWgbx/NdZhq1S8OPzSB0/rxc
tqqKdsqPQD25b7wZJMykgJQlp+8zEEqahy+JmKO8UvWfsgRv/nvyjsrXfw4dDcyR
NJ4aF9zcUkO6NnfeTq+HS+xn/eLcjb1TKmmN/ZRBehkQjig5q3cl8TA5gQ3J7741
04HhWq9UEzEpdFOxKh8Vk1jmOEMPqUZkpZSAPvf3/NR8wolAztMz5uueuzEvX7PZ
ezOErtITX4BYLLTi1Rd0+DcgLM3wC3ImNARWSosxyGvGRjuXcm3fjl+xBNmWIfsP
3y/mrXwaxmkgzp3+wLzAWVIgO2DQlFh4e+N1WrSfrgOcN3L8OZ0D7NspQ4LgIOP9
Y9ty1Jd5i1C+79MXuYabNwav0wZzd8hwgZYtt3A0TPlTCY4Kgrkdcg+3BQ84NpTc
Z18KSROED73NhH8J56MS5jwWGJNiWWEraOvDHoVXuduETvzD7C44rzOgg+vwhGAB
wB7LRoH0Y54DlKY8dacZoXrt5c3/oQ+q1UYmIiTR65rEjB1QKUMxB9L/xV5SwUbl
H+i/IQncjCoA2Uai0EWWfoR2oTELY010rKCDcVIe64XB7qd0pebfG5dOBop23Wrk
1D9/ywnEGcFig9HR1wBERm3F/8i+W5i9u9i60JPKW8Gu7RYNo6h4DUg9RB4lsOZU
Ytan5u/G4ubvyUjPOOfcoHqW7HxpDJP2SQJGI4y7swu8pts9p+p87C6Bj3wSBWq2
pD9TQyCky29sRR2KTn7Pn9RgiWO9nRp+en9qaGegIn5T7+IkKc9zZd6NI+GqlD2Y
0hmXP6CNlkYK+r4SDsTPFCoirbaG7XeheVRdBPlyez/fUlpZpwiAjOwPgZsQ+3jV
s/cFwt8p+7lpNQITWHeYcPkNRFHjsolEFZTcdpxTJ0TBBrkGdCLWrcb/jOsG+yun
uSY6S32SW1tCKZTdKj6oJUVu1TrHF7B/ohqLbCPkhcZenuKFUUQz1oUqR5ciaEAE
BQLhUOKuy0JI4irM1eBzYtlRHzmFLtCPOunqAebfIOi2p2BgWhq6m989o9NQlRsM
WRLjAZJZF/SQDcrXCzoEpQy8B0nz/Y8xrT3+qtmBpkq4dVpA8C/onrtGNHxuMoIk
02Gk2sH6LSJZV1LnYR4bn5r9GaJ/+CB6smT50NINKXEzwm8TsALFqtLJzCjYctLg
SKFCZZze10HtCSoFHjDAbsPC9xOX0NmgCfJe6DEGrfxZrCxEYbdsS/x2ges4Ocjz
ibWBApsYDtpxBV3sztMmTMsCYaElXIv2Bs84UeAXf5kFINDZf/SmEFQFN61bqZr2
3WBY/Xu/0PYUAOWH8Am9ozyBMW+sYFr5xaQYA4pQRv/RmFweLkFIcn19PYwjY5WE
DUxXeHgmOEfwnaMan7mizH4vGf0yJzPbMY2RGjQh0x9yIhAcb3Vm+gfl9vyNf0YD
5aaEdDxwQYRkGh+3KeE+zGAAlWA8bvnG8NllauwVVZQBcOdRuzBnWAbRcM4obkaO
dgyNnWPtf9uP0kSpYzgKlptcIjhZShzqDUVkTcwpzBPDyqFr51sTftkwR+2p+THi
p94K8Pxj7MRpQSvrqvFWFrHnSthIv6OuDr4mZR8EIADVs6MGJn3nop3aA6chIkV7
7m2bqTV5xRXUHLiwlrMcAvmoB5Yy2eO1U9RPuJFsy75IeKvQE5C99xBWqTszwMxQ
/WKQiaTn4rvMNncDFAzf6qhU/Mllvwef8uEqKYLy7uOxcUMUGki2uWw0F87i6z6+
5PF84E4BMXqSGLdcDJADj0QT7tL1AenUIOF62a0nmnbMTpH17f5uqp9qkFmYn/gn
3cFlXPz54xN3GNvLlW7sw+VvXphDzb2NcXE6nCbX/qcFMIkPWK1xBxl7e5ci01+B
o+sNu8chVday1klIKUOFxQs0pZksjvppHEiu8hisuxPrO6Pj7dXEGj2DM41sU2oO
Aks+FFawjhd2lbPmF5DCsEHvHyN613Uaqb8OpTqt2VkS6qKzsufvvyeNhbYvyyvK
FYYOKid5/tzlQSb0ragxs5IVyLwB3PqeLh3xY9mi+U7Z92y6xsA7r1wtlEisxxMm
hSAgsPqHTE8H9GLdN9rmherX88wXMHlidS8uOGVl+LfmycfizYeWztT0J4wu8doj
G0RBcOFC0P7+oZL4WnZnit69U3hHYLDLFVjzQcVRtkPnd/ETwY4nxajDPWKb+sFS
iA/I7B0LIJaZ6tDrbAyqs6Mis85D2BaiTP0OfkpY4VQbsd6hFfQZ0BEiGr2rvzHY
FQo/VgEPRawdN3Hx/Ui0zpm5a7mpDGxmIaG48n49qKTTzFjvuG51uKyNC0zqjtwo
fTmD0ubM2tkRYfMBDF7RXPns5oJJu6cJir1kjqkWe/zwd7mBQOc4uYHxkVzhuR4A
8wMUDIFDbkJfNPHtK+RhN+kyN02Y6KiSPXC8wkKeilBV6menKzWmtVtVFsR8bx2h
PMTHX5uoV7sZH+9FN/G0eNPzYU0sQ5LBlBb6ARXAoylBUsPCQExBTj7g8gqkE9if
aZMif2j1zE4N6ZLcotlfLWGfGmaGdYNL2Llsi38V8uH+oM0tCFSrR7L2mS4QSrjE
b73DXEnI4Ikhj98onniCmEFmeXaoouu8SencVNueLiqcDctPa/RjaKO9B/oiXjJk
Qa5gX1YSAVJSuRmii9sFHHKSXcOxqBCteJXSB6OlLLfLorST/2foJohLCzlqmwZR
4baQXFGhse/bTPmFnidJU8eKLJyW1FwV86NUj9+TgscRJcSgi5cGprM53R/j7zfg
uYHpuPbGHDsmxKyShNFisL0ANfjilGS8eoVYRPZOBRKSU+eEqTX3cgNi52fxynOK
OiyIwtu/Nv/1LCHGrcJjZ2SXWBdpinv2+g6AfwmjfDN8UwClIGEdatHzoPyi3G+r
W/tKROTv090o7BgU9CZkLKzkRRyOe7MFYj34Jrcwp6rIIHDiQl+m8p5XBw5C/4d5
+SHhi9XvxOwIg+ibnJ5Zt4ICcWb9tVzJ7nbrOasUy7B/cqUb7TY/LWq1YjdLzaGd
r+WoSBr/pHyYZFg1XSlwYHFF5qbd65/bP6t5rtM85sxfECWsQUy3KkNq3g/46JmQ
9VUNlGea8IutFRWoi8IBybkL1qj++2zHXPGVJJRlOAI5kapdLPto8gfhBTZFamtG
QY+TomvbE9fItHdnpq3YPURPf8Ff2WLzOBBz/uMXk1dlxlfObPl0VJ0Ewm2lqa/Z
enudCeGNYY+4IdJiBogqwcswsp6X6YHz0fMI7B4pEhFnvbhm0kJJL2lqFnzwBSMa
lLxUqxHAJDkh7T6cI5WWX7mk1WcxrvwbPsJmgXVMBf9fyFcRt0E1qTxMzQ3igS+6
PwTpj7MRTzZf/orkEUvcdxjh2D8yWsAbjwZp9bxZl4wbPD2aTAGllQ6EVM6WdzaG
93yg+f80Vthy//SdKcun6/LjaOzfatRqoDqHbV8E5R94cnTr/o++/6d3D9IHUTi3
wStBSQ00nEZH9cFGFuK38pmsJAF1NcYErDR+HzJbjuRI8gi/cd6u9YiN2MlXA2Gr
SsDMwV+Y6jSb5icTZm+efan+e6LgkofiG++FSBpsfj4aPOnn3UcfYRuBJSs/sEl6
+A0J1OstFBHO/5PkotPr+sNyzr5/IWRhulW8BGmoersUWyqCJXDyhc26a/BzWiuj
AV05WJeoP3ZABeEl8T4zLeaVdrff95Lv1/aP6xdtaDsZb8fAtcKCYeXHAzsSpWXi
aATingEiQpdwEWDwHj8yjQJV02DTsGplcfiYMRb+Gk5ucSWXyrRwFfjasvlqW7qs
AOzNqFAj5QRDKiJDjNlOKjh1vYCU7M4DtUSHQcl4Yv6fHrMU4yqhtzkVqyB5uvKK
mdLh3PArPr8goBkI/9Y8DtSByIlRwb8HiwTyarICgr3CxAqQ3A1NlmiFrHvkKPn9
CkPb3qXN1+RLZBjAZ4Acjaoc7VCvRm0FW+AB57WucNiO+niWsQ5JLOP5paxDGh49
YKqUtQtwI9RnPKGSIOiFZ5UO1NfU3qV2kMDbz+y4SFKgZqeUmAK39727eaKQzD1m
0n98xVdSQHthakeW1/wSVnkGcu6e7mRBaawmRdqFbFRKhfMkMhPq8zcxJEdi2swT
X97FOKx+QuSiXzxjqq5nx6QDYsDtl/J7F2803yrvyp9dCJb2bcoOnds8qlrn9Eet
guWYJ/07/a3W/pZOcWsMCNCPgZ6j5oT+SWrjLoUwkoYDhn6fiikzxlFFWgqhuEzQ
qzIwv+dMbCtxUJUOLX1gc7fOPsmDEnNNElWQ4lUzPyAOmyH+KTHL8GBPmpKRnDDV
IIpSMemnubrlan/iQrlD21E7WDFqbBHjsebuNVlj/5cW5F7h/KvtqWZx88FEoBfE
xMa+MLnSTbHcXolUAGrmotMu309f9djG9IforvEOVabD9OiDBHlBsHziswRPw8nb
tZOnXf/J2RkeLK3XC0fBOat+orPoQgB7VYzoGm3c16KdtwkBMnRe0QXFE7m3OGgS
LSdFLkC8jD4ULFqwVVnI1B4whL5rKkbF7Ll2ka6v4IuB/dv25FWe1ZOoj9po0twX
FoyBDUwpx9/km8LaTTLShKhx0jAALecM4yyEMctLBNj73eoONDtZNrViflIOZbVo
On1K4cgUfIPwUT97zCCuj16fQS/vxI2l908Emi3VgLNl5mR1wdYE+u+RnzkA9B4h
Z02jkWHPSewvLctNCckuuWTxalkK5O+YQX8VUGgHpDPKRCzZeYRsOYqy0fGoEvWY
NCjO2DoWkv7A5eLsAaPaFo++Ap3TztY+oFvnZI11cv4h7kQyodb1woPZbGoXYZJ8
8qSEO0iaZIP1fXm4V9OSGEJreJ7Z58rNr1S+Alrurjjew4Vzhx+imURrNM3kWGl5
lCVplfPszfvucNyiEn2WtHFQ7YsADLtu/gigctCsKLpziNM1sC2r0XCQoCIbCwDL
3XHit3tAmwUErJm6p+sp/HFXxZW2WX/hhzLbP3MPY3819HayXAhNLlXmoa8s3ZsQ
gDgcwjx6RRC9yJpsNXrMWvKUm07sD9bv42i4HppkYWZRzFG1F3Ti3JFcGAnkHukQ
qx4NjizdLRyhUk/QRk20iBh048FJLs21oC8/IJqDPqdqV82F3MsyooHXK9YhzGwO
QKOYkeEHmE3UvXttiFZv6j/D84mLSNMLazUZHFlOMUlZf8cG264k4aNhwHtGBfZM
u0PbvMwhoiN8qGr+Ed81k9tVEjf6LTw9xfkZUvKWwWsr7O7fUbXkvqX2IGf+oML3
Ir6Q9LYnukbLd5LMLQ8adz7y02bShQwEMCYA7GPzjZOuqmLKJxg8nUdnUPfA0iZH
8EUOFBSqamhQjCdBUxs97R1dhueNlK3y2N5SIqpJD4daqS2cs4YaUBa6/8M9JL4L
yf4iZfrqA6Zf0uILN2r0ZR5Nma2bNwxbcxifwyON6fA6W8XN5SR9RxeBGMMn7a4x
M3MrL6s2+fFTUWV+m9meBtbQBBLsXJh3uDHvs0gp6hsGnJAuwUnrshRW7kucFOtO
kQc+BgvqGsidlTGXW176sdSPwroazMu3FKuGTScXpKi2TDAEUMWHYoX+I9fEcC4V
XAEhz2cgMh8rJbD1ysMlA6UzWGniLD1Pb6g+7VTKilJR2jpvD0qPHoujuyq29BX1
KmoZDcr1izIZb+0iCe8mTaYGuJS4BaCMAastqJnYeL3xy03l4Iw92pWQPGDFH/4K
DVXlkh8SnjKXqjQh0wLuTzvACW+inYw85iNHGhT1bzeV3ZLn45WPt1cOUjPXDze0
WE77AljLbIknBXJm0JChMfL44XfDgZycYzoRdbHuQ6+FZO6P1EoTChNPz51QSaFY
qIGN7OKO+1uI6j/fQc9OR9bkb1NzMWMfsQMjZrYjAk+O2akyA2+6xAjYWwGknoYY
m7e5n8pLnmW094n9j1dWzApWGNUO8PK2tOEA2Rn+AARHMwSRqP8ARsuAUgqVXTBn
Db/yn6QvlakW2zY9EYz/5oOE85xX0cn/MCNkKAcru4iAEN3ouhZHuvxZX96/bUuV
vCPuErgO2ggLRmZTXWsVjMSQhRldp22kw/j03HJndiJjRTupYLYobVpAqGa613+m
w4wlYQl9fOw2uWYuyBr1cp95DfHyjPY+W0DQgXGtTfuPluSCkJ2bqd5/nAjd4pNt
wThQyh3rHDDbStxfNOkuLnuQuv37O2SeutvardEZyC2BcgK9iV07mQBit50xYGDC
fgqT718XIBUE+A8ZzEF27pzRCECOHHWkWg/8w83F6JnWx93ccEjkZdXe/VLOj2VP
ug6pabp7ieSXClVcVMHbQjpmH0hOvGzhU6+Wg9nGDaf9FxuXzWooCP31DvlDJUJT
0/7GwF9lrYNG6CXAIoFFFmihsr2909JJh7zAy+V6X8KInqXaNnzlA9ikORmpB3oC
J/RDZyxdODapXck+cKnazfxrthhLxz7ZpC06K2ipN1pfxf8GszJidH4gESOzRArk
TLp5FBZw7ByXjbuZFt78OrYR4en7Q4BwvBAeNxX/8auddcrKW8Sot/lRj/LjGsSR
xdpfJSo1fMYxKSN+q1Q+N56e/PkK+oWZHZRsbD1qY27rBjcdbfVCygujkXvyE6HP
PpdM5enP1cd/NM0EEN1NF8gjZq3eKTntyq7nAS33szMoc3T/SbW0x6nq971wyhw3
9Mhr/Rjj3Qfc5aEwfCn7HHmey+UbUtL6Ce1tEeOwhFrFHBRl7GXcViIrqabK6r2x
PeesqpLGs+8fdTgNMAU6qkAtVC/9KgNZ30tgj+Z0IJc32sNojfVG+zyJj71XXepj
jpNC3oJYWnvRYZ24ygT1e7oVHC4GTPHhCF2XGFpZ0kMx7M/nEOzk7jfOqDJge12Z
674PB9X4PMGC28Fx/aAOV0LyREINgaIvEOnZ9todSsCo4VDwG20Ht4MflPbajGXH
aZsYED1Ve55MVVF+FvnTBp4AudZtMr5a4zDJeyBZVV5a2Ih4LDPQImR+lQPVslnt
ABbAykLdh9+KnDuHcNn6gUZhTCZe2563w/apO2wTPpVUVrtiw39D7Bynt9cVJ073
sxXPjrgvKIKw+xTp6hehYOmxSYuyNBMYIXKQ9ZlbbEq6cWknoubf5LetW2ZSwbGj
dtrXi0syOplxuVOvNYqV1cDuIWjf1YsGta2FnM0DX/wRSrIMaDJcVjzVdmkpXSs4
GJ0A4gBxgBbnjqUa/OUUqGi3jiO5rCTTuybUQ0tyG/q8kYCZh244jox+ZPBo5J7t
0ZRTJBMfYEm+Btg9CoubB/D0DMHIpOU5ic6UzYNvRNq3JpBilYg214xnzuaQFyAR
U44Y+yGa2TgueCe/ClWjVHpTd/1Uc5K0KvUwEd8ha079HjdQ/8z8T520a7+UxhxQ
K3mZ6LZ93/jIfMCe3kkh6EVIUNyLyjhelzvT0DeD7rIH1iNHxlKT/mFMXAhJ1Exj
y29y8RQHxWbZCuxWxCWtoreSGKwFtqAUDOOgA4pYsMvKhov3IGNPvEW16SLkFHIQ
UdthaqhYeFbSDCoRvcik0EleAxVAAt7uf+qvI9hkvIiXLCQBMP09uzooxOC7dCAs
Pq16yE4/ffz4UBNjX5x/xstEtvon6tHVklF+nZHeSSr6xwFYfDjvnNcJYDEmKPEs
l6nJ03wi4YMfmK0ic/VcTBqYtxqOf2OPjgPEbUK0AerzEUwrryv4Xbjv/Sk5SOXo
kwd7aVWOU3el9GUBJSKNSQD6ORJpZtjqrsju2Ld7F3ttgz/pnlRNCWF6U+V5Wp2W
RqlaG+gSViW0nDB9Qc9QfePs2yJcwbADRqHdEXWz2BdZ7xeexR2M5SQsUNNwCSOz
hSjGG1gadMIt4i7E0cZEb2uUnrSA9gmo+m9FDJy7DQNmccDoCsMKI7YU8EfdlrR4
Dku8i9xCJ/vZ3Bn+wIupOnuLxqIddfEowW+e1qLou4zyyrePjCOtofrfZgZpd1DS
G6weUS3SWY0K4jro1/dmTIlQYTp72kALwI/36ZL9V5iyJl/q0FL83iEDECvharfh
Xav2O6VvKUAHg9rOZkV4Mg8eeOgZYWCon5SJUHFJmkCrPbyAEvDl1SFqjhvzuX7H
bBFaUZphflaoczXRGq3BCFFpC36ueiD7eJ9f2wthaDy2CLUK4alkFR2Fkhmc+blW
GaL4dwNXJYwNEgWFKa35aCk4pDYvyNMfhSBgP47DlBbjHRW/+YcgBe91E/FOPO8M
2wOhbDN+lqx4miE8e9mPtQhki2t6Tp2+9qdnZHXpiuisLlVgOe06FmHF2D5SMV4X
036dJerDr7QjWvWiK4MI3mhu7oheiFPQ37QeUgZO34vixdWWCmHKzQiOFdXg4VYO
BJxDCwAkNN6ZoX2E2/RbMJcF7IGlHkjkrxn7W9O2Gdu34U+ODugIj5aeUcrePcmN
Hnp54h8rFbQQvotqS6kphHWMqQQ5uH7IjYVFuxeHO3rsd1Z8FfFZDkMjLK0d58+G
EmDUUUb+UwPD9BYB4q2aagJz6HiXPY475XsFE6T5d3Am5oz87wKj+WcFPT3Mbxwa
jIhhhKemsk/WHOBQujLwd3/H4V7pVj84e6/CuHL8o81zk977lH8dDQmEHVh7IDLI
e0FIqT50n4iGYfLS1hJc0YS0ICGzDTZr6xSxRX/PklSwX83bXdCjdKkudLyc8XyY
AJqN7Vv58+pdrN3FYmNlbi/aVdu/3vwoXhrWmAxGpMNQS5lV+/ns5wqAttRzkD5X
TSpY67xfBi0dKrLKL7mc6pv84N+7xV0geD/Gn5+m8qvBVBCtBlb+NoScIwum1kW+
2Wg0qcUXsAdGBY20Bu9HhABCwQMvLFdf80V6vYweU82mQMcscYLEYPWW4YpgK6e8
T0niuVOvBrbQOX7hYau0hjqHNC6Bk3IET36EUNAHgiIPheamAxACLT4qlexx5+8g
mmYez/NW8Dc9LfMJ1FspbEv2n7/TlE8GM5e2ni3YiNbghnc4+5DhPFVdECHI4Bli
ty6pL8gU1uk1juWUSe2XhPozr4N6mhK/qHSEaHWZilOg3bDNBJWat8SijcgtapDt
a/VjSuz7s2wQ5y1W9EbG7Ctk2QmtKfamRvukAqeDvs3Ab2StkmsOmoQPgwJZuMGJ
xFJ1Hq4qiD7xp33791jlxZzJ0pDsP2sgXNGjriTgZV77aDZT6kQsyp31lfSWDtZH
H17vxlkxbV96SpMueDBrSe74DObX8MhX2Z9B5MUAPUUIAhapOdaRIxfwClT+DZ00
ckop1dJA13reixe6UpleO4rjwOnGIBUiSRUYMdwc/lZR+UitOlOjlMBBosI9mWhJ
KE4ArtMBtkmnR0yPAeYC8lV2Q0C5iZdg50IpkxU2y8iNxvoyTvODchJJHD+kuXUJ
TFAUhiRMNfU9tzN5gW4XOB1CkENZHTnhSe454ZNODMN2o7eNhE+UlKP77f3qJbQ0
so8XrQ645OkP9Dw9KoFWfLy0xeIr69DF1rK+83JFPdjWaAx6ZP5h8we4zB4JP/Td
KTb5w7DCGIXwh9MHRpFxBOSwceS1XRnN8zf3vorW/lCJi0W/b2JywiIy3RT6711U
3NyuLPcVmJFYSLFzi77zlmvT+2uukKk3AXgh18mO8u1Sgdb9t/nj5bDmPZTKjr5K
mXfUCv9dNWeRFK1IWnMSSHTPCI0AS6PY05IBhaa6rLK47n6aGxXiycP3dgGKqOG3
ezIsWNCGwhnHvBHkY73sUpIyZIltFlOrRhWBT1jytSBSG4B7TJJMW2gjrARRde4o
6lVwTvcv6EnRgZjKLerR33RsUePAEIMfnnRQO+Ap0GcIjzqGCrvoPLZuAh0hFiJP
nj1ymamTGCap5z26DxCIubV8h9nUp4g2h0AxJTofGneYH9OhD4Lfb3+kU+iZT510
R7+PQermTjyfQ+uacHP0NofxP+a//8bY0KTZKsoSg9jgV+dEko3+8UhhXu6Du+Rj
wOMIyQhks8VvoKCMFNX9KEnHy1aM6J1lwUVPUJirZbwJIsTc8R7krDFmc+bjHBvM
JZabDZmTauXSu/5CvtRbKAcO5mJSEBjLHsqP65DEJuGvDfIB2pjCnkVdKssUgOSP
+UGPbeN+Pfo726/UVV5gVutoF9BUfyh+1E3HbLI3LOcbLdnh3rQrta+uURzhHBrz
AaJFy3DUZRwfKDaW0dU4ngiXqwWgCUeaK91njPsz9OZM8TlHJ5qwxYizRu45m5n/
TCShHu0FeKEMdi4Heow5gxmec9sXyqHEopVS+PsUBceUjIGAjhd91wXsGN9JEtyO
yFSua8eMpYF0CM//W+sZxa3tTi4+mSinaiNeqYk0FgVyvarDD57N67V8DmI8FkWF
O9653QxMpz8VNKjA25bEjPo3ZZx+16REzHzAbIVIVbiV7RmJBZ20/q0RPRb3/iZf
XuLX/fJyphFE+IYLcSNkXcR97P9nWaN1YHWzk/kdzdtlJEUtnlx+KjiBlPXnufW1
+eHjXDISUUJZdJEsPTgPO4VB0RUJ+SfzYPYjGeq+25zReMjtauAAwp7ySi+l2wF3
rpJf3s4dmAtStdH9NclHtNr+/sJwx/DRooi3Pw9jbelaiY7fd6Y0mHRxbrdpqp3O
qy6Y89ROGXFmet5TBmthf9hZgWttuoYBZ4jsaD2u7xenqHCf6T8GaukSicenkGmh
kT8c/8M3ZHFno6pyMrpsACmyUapm99+yMkQcPmHP2+wcbLpxGp43Ows+ckWPb9OP
bvSzRSHfbaj4aYZlpbeqcNsWm2YGq7pI3NkBq4J+6aGrZ0F7O1Dq8NRNHHxgbxmK
5Y6DJoyV4/JwLcMv9p0yKHTL1GBUmBrTgRCWSH85X/kHMKe1uHOUCEOB/HtQBW7Q
btDUma6TKTIb82BjV4kILkTY3hmnZAe10gJoDreB4/plfdlAhcascD+DcLc+K1mt
FfjgDkkum0Vzpl2GXl+xng4Xa3B4fmaij8K+PWFyeMgqNS6VXZNMsiwHqkGQyPTu
Fq13RcyUQ38vH9kRh5nLVFXYmxYlqSmip1dXMlTjm783S5gwpr6Wuk4cAI+WEiwP
gWUlz+xk5lx7ZMoPt/sLvEdxLDt/rDZZJ90uU98FM9Gr97lAM3OTGGj+qbNxoRGr
2cyMkhkpIRU4nVZHwyjcTr3fhhEtOSC1gAaSNJM8bvFJLdYiYoQn7zmoydQKbIta
tvuCaIVe6bcgQXTtOl2EqkRmsJ96Y5nRmf6qRo3fDZVbx4dHLYSpvHQaYaNu7YoN
73VYWOQujzRAZ5dFcHP/RJZdwU2q7G4Mg9OflbfhWlZGQU4lz/l3I3Q1oFUMm3KH
P12UUxEz86c6XZ5IVjK7S/0VHYCKj/13TTnHgUOivx+Nxy1DqvPOIRiuaQhgL6PM
i9doXItuYOYg7HaHGFWvrel2mhy8OoAGnoJtxiVDXjkMrmwpB6jfa7gd4CCsYd5d
joZ8WolJneEagaKBbP4FlwdGdi9i05at1aeUld9vM9eLlozwynVotzZBPrukBSyn
eyM8NXT9p+tpD3Pl27onranLMm1KcQNl7GGV5505iXZMsX5syNwmnRvAG5eNl1zu
MMvRly3N4/GYWXzrke660YY/YvkKIzk49OUcR1uQbEONGGc16XzyZhdtdOrh7FRN
hO+SNJMW6Mk0qu6fsO+wXSckbgDQazRTjyZ9gSFxYM1dHMmXLu0vu8WG1Fbs3Px6
yD+XD0aX1X0exHE+/Nm0o18n7N5lPpqWsI2i5EANmDTezW36moDg6dvd4fpSpG1f
6Lyu4SgOTBbmQAj4GyBnxK5bcLqS9FlNT3CyLpUIwDomUtLJYvlUN0C3yPuz1x1l
NQRzKcZ1qrUvOgStX2WE9tkkDOUcxkOHaAHTTCZGZLnmWp+vqmaAGmoMX5F9H42n
Xl6AUYIUBWlhstPVySAGsfGuq+pHe6a60yQ8FJBu93TxeSWj13e8nbuXnUWmtgHe
BodsVPD9KwKijcivQN6qUntUAfM+vnu2hSYn0EhBluqmsF2QIRkfyG5K5KcC2et6
jRGQ7gPiYxCwG3DsxOCgdRu06nSvntUAnGYOIyuMx/Ld5qhBa/dmWkpmp1Gtp4VJ
QJs+GAKX6K1EEYUOrbaSntpjqz+26Q8dmR324i5lRoclOFcIlB9Olf8uOcCOg8+H
kUwkEHXJ/OGgEqSf/bb7GBM6W4lpKriB+fHXF+w3cTtfQvlHFtwNwV4+uTVarU00
VuE1RPcTnnZNLN2SYsHi5g5sj1bo3s9WAaU+Cyp7xWtBPr60CdJoDdwl7HhW7rj8
MpT0RvbucN4ocQhzyHjvqcKpG/yuck1k6/qsl9Y8BcZ9rx0uso9PS8uYX0kIc61P
+Jcaqy4sDTvDmVF8N5beWfqOZN32q7EGKGrOSSgi0xjeovRtaett+Qy0FwU88Q5H
upNZigbk9o9FiqXmdGJWtEaOE6emiNIQnYUUeIQhgXBpUo28JPS1ZVj96v+GTbSQ
GV4O6hXB3e/4gbRGEIKqUmwtQHLwdDMDPoQkWi50v4UmP5pyzHt1MUqyQmbui8No
V6gai8oVfzqJUbMkusl5aNOlFwZBs7wWNx7+mBeQFBxYJwl8ZXtxyP5y0eT2S3Hj
eURrksFJZvnoXNjFbrsC2UxsarwClzggWYhpQP0zR2FdXbfdiwPoqZQYRi/hskKs
coo00DimcU51NdWenMXBf6ILsaP3/F66lh7IlDdXOP4RzF5GspMuvOoN02RhdBO9
79F+Hv++eN5qj2XH/FsKHaqArln6RkjPM98h1bO/wsDkkQI/C+KkeDfNTKcB4A65
XmOEAJsOerLdsm50Yjj14zZRJczE6wDqu202/4Lq3DMEunrPSeF3L3b0ZNNtGRUA
5gl5LPRxJeloSmgiLKvR7VfryKX46wjnfDRUxMYI0c0syY8oRMw3i9pG0nbJPCVX
snFOcIAjbxM4h0k5LTEo45Gj3bhjb5HWC7lFm97pquDJm+E+GNLPGgetjR+G2zO8
+Lk4rTud6zsrlAePLsQfgmUVDoL+IJHZBSEb1HSepMBNnEh0YvQNcc+zwWT4drP/
ZTH8Fbfn6IaAwPY8flHGf8EtPu/sV8/cgfpD/B1Ap+Hf0v6HKxGHWL5LKP2h2CzD
xq2rhzpbliGiEXd3+o2biHgQAYixn7gr3TPfgkaeFsfutkyx+Ncl1vXjlGYfRI02
g3kM8LFqp3gpR1N22tqqEgNppb+vGIUUgmIBkKLaQuv9udnVXUSChsklIw0mvJBF
phpfmO1Zelv2Y23KF+O3e4+BjFmNaXpKngFT7YZpz3YLQDtpOHWqt2CV07GLeTUP
fk/lNX4Moh2ti7noxcXaCuztk+KZlPFDZr4NYmMBMeyIUqrEQPZydXxLyX+hKEKl
wm7JV7tjyzErNw7SqTLE/2fQHeN2bDmWzO+YEHqb+qSc9ZUukQuPq0PXiAr58owf
2XswxPBiJyla7QN5eGSUqA87rYCcRC4f18jRYOe6sm5Qo845HCP4goY9yKBQb26r
Hjd5SMN79YDO4bYx+KSWxMKVbcWrG7y8QstmRc3Tg4jBQYfyD76HZjEBwJ0qJlcD
xgPhHrJo0ulrNBToTNwtPYb8CElZdEpDooAhJIUzwDEQ5p9qpnvpGUs2t68CZ2CW
xFSfqgpPe3deiylImK9tQKvEAv5c+wdXjEgkpIIwJRwPkqPqqMtKanDTvu76jv4V
fvhtHwmYp/e/Vz63EDgk0YbkHLQIFdVzRhK3d6dx97xXWNHHPmJxNt51uyirOx5z
AAqmPuZ8sFR/HL4vhohHelUN5yBSpFCuh1GFpM+M9ZXjV6hYicpo8bkOZ4LntgCk
CeSAML0tuvXn/A5iYcLcAA6IldfByTzeGRrgeoFkBQ1A/T82qNtaGtbvk3BJ174v
gch2CwdDeAVuCrWPZVCrPy+jhzCJvIieQPaxnrjKgMphgvkpI9RmApbt6yT/BwhZ
+9lCSTh+M8zhipIDHjOYvg9KcbfjyfNpxKeSrhl7NyM8dS9b5sZ9F/Z6IcW3AQkd
ZH6hQFn9IIRY0aPzIg+2eZTVdAMMat7zULfCMsZpnz0PY9mVKpWZhnIb1iyBNOEa
ytNMHxbQKtIWc37qrWeceBozm0P0pcAHG8yILYcdxDn/cv4tFBcd7L+p/tbnGC7Z
y8t3gsjb9ngkNho5AVcDjea14nXdNgAWbfUdpXMSv+rLgtrMfA79Annyyeli0YNk
u/S/jU8q4uv5AZcJAeUkX62YvRBlLTdP49wRxVk89FfdrEiqJhTVjPrfe0c0i4Yn
W2+hOU9K9UK9DTcWz1E0Rm4UDMOl4cEpsttnLDe+ZcdGx7RgTvY3fZnfSzvZF3kE
Gj6v5qhJ0/TOwiIILztgrd8ymIsZ3QDhoyFgSFxk5vmDXsDhLrM0x1QO6GnZAbcV
GvCpePczQVFgesNTKZZfreYQVNN1rYOUv/Kcbfbi1CcLkCwZ6BkVzuIekIY25Vcm
Kn14NL7h6WtGwlCFYkmfL1+/R7NXDsDUB5RgBCcgroma+7sL88McbrF0XTsl+s66
7X0Gc8tCQw6eWfCD09mF2dmNQsD0GD8hSNGd2mbiuYs8/jBWLSir6+raGvccycrQ
561sWi/ZzNTjZdqydRC++xeNq1glskcGVVvPd8cu1OdAf+T/aNx2TRKl9pei1Gar
/8EuL2V16eHcthGFr9NuC83B8hlAC590+2d2OMMBZgrJHc6e+T2rf0GY5KSzxR+D
kBIMTqXYBm2Udpi/fyrIqlaDtGAJO70MFf1oUO2mPW/Z1KQ5zxZWJgx19zeWXVlZ
FP/qG9xwrPcir689jT5CVzz/+i8CBSvM8NnLKkhfuG+0mCx9oF8UUOha3AithnJY
o0f/Y+25bnz1Mr77yACDLOd9izpbzwalJb0K0q0Wr0e90ze7XD+dMQHdes//LMpi
sefNWo8X41fcUDEW05qKxXE6cX/Dx3podldUTLINrnrsMPzINdl0SsT/ksCneu0z
2zNHjWRqixbL121HKmHGIMmAElI+jhcGh52By+hQ1Uw1MozpJgkBlkmkIEyPmKss
NMkk13A/JFj/kWSgxcrSJhq5JK+AvzCuTl26GmV2//xZqtvJWQ1Aod3rFbXDwjpr
HRHaulSvHOjrglTOE3H2GEX5IzB6cfCbzIUbVsEpkUBAcDTCpmMQSD1PHB6+fJaj
rONJKL2wC0jBSaYkwyWEHoZ+C8TJt1aiQ19BaFVHyF5wIZjGAN2fhKlpWUvtuvF1
uTz1CTwGn64FtBULmISv+XpMHRvtTdtYP4IfplAbIsCPEJtwiTXFJ64oH28hPldY
TNU9KWcbii9r8qwlQCrK6GffHZvskEk2X2dGYGqo6gLmXoxxLHn2upaWBbiZFyma
rvW1jl06HS9azJobiDeOq7wMDhPqlRW7ffnQsXVFECWAz2aVszWIwIS4PMOm67K1
h61iLITxTJ+hM4WB68TfFjWMnBrleZNXXxkbRFbgydZ/9BqP0pUL69OX92/E8CPY
dd6sqxKknkbx83Ru0AdbtdhqoU6iZMYLJJKabCHi2bi/JRACbtJzXgyl6Tj6O+6k
2ywj4vGivTT3Hq9UQF7YG6BxaOSZNbtAU/lXoSEcnN/OY0KZ8efceHiNXAGj9oZb
yu/e1ZWnwP3SKGLOdD7XSuWtY7JGAS9TAbayICrO49DEoias2dEsZ8o9F66zile2
+NWwbjgguvCkjz+SkN1lynYzefyfHKBN602fK/RLrCMcbbUBvA+ZYEl/O0+baIrn
m7pR0dd9WzI1R4HNF5jXgmnvcSRAC/SMubejvY//SvceLTNgPR9vUW2VBh58H2kY
abtFw0RFscbrjY/J6mPG5tycJaE9wHto2sFpVGo7/swyN9eycy8hwi2PTyOHihtB
qDGCWGmHAZFMPSDDfFb+yugnGUcrO04c4+s0m2SIdNCoAoVg9F2llFS8g/tVN0aM
Of1dDke+3e1C69ZmN60ug9vkskQ69iGhB7lbOUw2cwrOcn35tn0KEyXOhL0rI1hj
hm4BPCieKs+BG98IifldgcJrz7zqRbo6/nOoxu0m8l2XTOhFmcPNCxLBsosTSvuH
Acn4JeFCEaBSAHA380a7dgzTIG7LSUF06RReY+HOXeWKzsiiC1KMjSZ8ibkVNdpa
WZv3vLw/4+WzRagvrCSLFgUjKnkmeLKMZ2CHAy6jrSKl7XWHBCXiZLEVgctBjNmF
zms1lV/FL9vdGu0HisQIniZYwihzsk+wRZaN9TApo3FXudb4XxbdBLWq154JSsEa
WsR8+XzhL6jqwpR3ODA97xhASX7IViQAfeuEaASnf+XguEfpRY8hbNENfcWrL5Fz
WCR7B+EthXkczVams2Ed4nsmvkzbtapA25P1flNTwdta3sRngZbJf30ny+mu/wPQ
Z3iiDQNiZp2VVXQVq0NtIJz6U4RhX0noB9XFu6rZOJwwqMGOePAtLSdch8cCgJCP
i7WKMkslhH0BSjFaxrtNNVmIWSwTREjHatyKgzhblBW6wztPRE2O7nurTvZ+DYVS
LhIXzLI1O74O0c9Ld5mnOXST4FfBO2gk88xsDocCtfeump2Hu5/5ogRKX8gsXTWo
5vQw7t71o67jg6nC1LUUOauS0qcblYTAK4FcgUwHzecifbd/F6Vek+CvJ9jkINAE
Fa1iXUhB2FwgEarjacLwzVoyWiNBaZrYZcS1qGjI6uSbaLYWQL0ZtHlxB5epNgiW
8R+A+HxEq6AuEi0AYYblw+5lkSMmqHAtJlcfGqfEKahnE9w/GupzyQN8hPfba0mj
TNkd5aPfPBughjZf2EbC3IJbprqPZulMG1ZJyoTX/xQWKYUElhwnqyTsWcpynSHA
ME+D2cgyvu3FR146/zh1VEoLIkywGGDDxyQ+6nycw6s332mjjPJAdZuzZFdIDWTF
Ui0/vXoTLyAcycHM8CT+aI5wShJl9jetOu32VuaTVyZpw0uOWxuEmnlyl8fqFeqo
1sDPnbO37oUDA8f1qYoRoCUhyeTGCubrSRrEBRu87Pcqt/fqgly8c42I6ZCe4AXK
2xKcEz0pa9KJTuIytZDxN58U0FLmh2TpSI33Y5Jpm6Ud6/ogs9rb3MJUa1ZNlFAR
Hfr9LHkFXyVPyJ0R8+kcz4we1onSOQsMMU8NtRqkSJL9ftovGPhUoGnw9I90B5f3
eGqXna915Wyt/S2j7X6slzsfBbfuT5O36vaQz0EG3yRMSml61bcQcyWyNwPO4jet
iJ14ja3hwgyDYeJStJz90zqoHIV0lvexgUoal01qDnhw33OnKXYm6rPp1Ahsi+3P
QNk0fDX5EsjB2qQSVNr4n/VE6YubEIi5bts78uxu0r6bmzWOyjSqR6YgeBZ0yxPs
Xs92XfhKHjb6Nr9m7waq0z0j7wwscRdXypC7XxeWNy521p+OikpvoRmy9BftM0vr
FqmdBfkl2MZZlfvI63yI6EDpzjdadMOrKlhA4np2Pg81amjYg1lV6Z09aTQv8csH
Un+xFR0vQv2+UwDdKw4p9mNrJXYkiXArWfy1kYLpskjoHBJiW+LqqUTGu4hOmvs0
xE9+pZK9axw0/Nm3NzYH+ajZPolwPvR2L2R25tfPbgH1kolUwNx3f/Bci3ViTZ1Y
IAmKSVmIb435NyzQx2kzgR9jYpSKd66Oo482vk8NoHWTHRL8hB9/47WkJhiJDyIf
3+AAGcWU24aKkwmkPYkWcSXq1+gRvrGEHdJX6McGCY+1seKGyReHJm/VDuLC08GV
+AF7SQU6P8kQ5iyoLuyJ4Q0FHr98ETvsJAPYZy2j0D4rGg55NBP7qxYKSQsUuXZg
ZUcLVnw4Bq6AuDw17U0tCFUyISrP8O4mTaTq/oQt/Qscff6KxD3Y0i8zAl0aM81H
MLBPaRhhIJUFqjutb0S0e5KNi+DrI0PX+ZkPr9jQud+WTxrmQDGkM9ca5YLCPRPJ
v08Zz5ThDQYD3q8fSdidB63Zw3G4gJFkhP3oe3Soi6RhSFruLk5M9IRllJG2XIr3
uSrgxgETRQP57QHbCPALr1l6Ijy5VCKJ5j81ystaSPuFuyWsWt47eVZ7QwqZTpGY
g27FmJ2VkdDtB6gVPyqdqcI5uQZTJkkIj+k9YskjQv5PJSkTgAAsLW8F4NKoVIZi
CCRCiKyXICRg63bhPjktWg3Qws/LRfJEyUEHs3aea+wWYyuD0ARUO2jMdYo8qQJB
g6w0VUFmbzGOU4nvSMPFBLhccDVilx2fzc0vLaxxuhKUWg/nM/WMuSfdAFLQ8AL9
09yItT/gABNGn3ux5iWWj0MGX1rHtg16wj7O3RT2gXp1srOEyn/K1bLRkp88u+QD
tUKdxfM14VM4nP2cFxYqUqSWlQW01F9xN4d17AnF594nvMuX8CKZAvqz4rQRbvyn
MaEj4e7IMjwL5JbzlwjVxr2hy74/CMH7K+29asjQXV1n3rie522waVL4pC5ItwIR
hslnYJ2TCofEJa4JNOw2A30jZFu6fa1X63ExI3HGKQhm1iSzOkv7GcY2hXTskdnV
qK6OMPn+n7TWgNK3qP28aCPLtsHBhosle3NWpK/tAmyxwOvsqiYdjGdBi3FPubUi
++PNroVlrOuvrCcBwftRKSgNztl19XKq7Bt+q5XsIbMbzbg23W0w4BfeMeg3wsTJ
IdmAtkJ0rG4sKi8f0mawuFTOCpZGduDdWHGmH2TKbyWF2G8ardWCJOLnEBxh7LJX
66Vja/Lr/Kps5Kg42Yi3yCV9dvMu92aIiGv/QMnjWv4yTiZWUymKi3xjCRbYkbK2
BQduyR9yrb3Hc2kipAG0MiXKfscrmAoea+TIA9a12rb+7HFu45afb2k3efzILLBt
OkK+NbmuKqrXXjLXCTfBo3om8XEAg77QPYeImcDd84NwQN3OKQ/El0Wb8MpPWouA
lkeZ2T/RJjezsmDU7/vsdg4/qjm4S7+Pk+NiansJVZKnZBf8sYm6iD1RT+nJS50/
MXgY2UAbLWkDIdrH/4VnPGT1x9mGzCv5hMKzu2SvZhknEkEIo2RrIWjglI+obhYv
qblsW5Z6fAJkR5o2e187BiGkPsyoGTJrnCQu6EdoY/AYurIP/emBhxB7Z2hNjAiC
l9GfscLWUONJJS35FSRC4Jfwl4d5GgnVlAKaBHWWowXZHEgydq/orZcZwJEiAWro
RXy1NZby9GBOyN+3QKKbT7ec0/hNtQJZMZKYsTvvPYz9v5+pQPAknF9YbOxBKuYw
5hrt48Fc4Ko0FKlukv4U2ZNkCSCAYo7BuHDWZ0jssF8NHKTmx5F95/1LeGxW6Gud
Osdwb/idvuyqeiBM90oAM9Ik1llC+IJZwBoGl4EgG5dlvdRnSd9QoSkDe9fExGLe
PR8BVGwfywXpUtmDG3zVZF3tMbl6rtkMmulNo7cfBqRpSnnb/JFmYFJeBQmQZhu1
BBe7+Fp0vY7w+PTY0xZ1za4KYe1XC1/SQdgE04a+FwPFvwLM7f2w+XbL81C9/D71
ouRUFXENfMXGeN54CB8q4H1AeC/SpYLX5ovtHCCFGt2ssaP8dNlP0zvcffZ40VWl
V0SvNvU4dr0eUY+nsItPM+LABUo2JQz3YmNBA5C8VU601F6FbvU6VdurFL6l9dxz
4EgzR/Kv2wbdt7UfJo6FD8WZPBI5XVx66ofqyzImMI/viDyjTkaUj3JeBOeES587
gAGcObon2D7++5K3gCfTqk7xGsfJHYrA2Uu/KC3lRWJc5C1tl1kwsiA0DhocOVrz
kG3zpr3ITPu6PzTGnrSvloVt3wLwKl8qun13tls0Kdwx/Wg2avT8zHPDT6IvUYP9
RXJnhtY8ee4P+wxfcd+/Y+INJHb7yMj1OW/oxGa0TYWsGRafy1tsNfqelQOqS6P1
1Fm7MYLipiN5I/WEVwifvbLePD1bPlDyqz9UswFQ5l//MZOp9TaY3jjE11zVO/uQ
ZG8bivNxCR9SgJ+QtLSD2U3J15KW4ekdNDfXp2djZex97AY13KgJM+cMvnYj66OM
2XHFTemqctgdu7nhqaH7OmIeHTkWfCJufNcta4jgmiLlm5r4gTKtGKmHZFt9EGO2
3acZy/RjKnEjD4qxBlsHg8K3bxLLEbQbxyvGHjcFTnuKHblFNYcmQaiDb0bNIvAp
FbGZK344Fb5ojINC+nz2ACIhz1g3TDf9DlXoJF/vj5gS/IgHqquyl/O6cTALuLps
/3+/LOTHvBwCNw8Fyz6PzvsffKfqukPGn5/q0WZZuUYYKq5VmmYT+fS/GAj8Ribj
Sm5qDVXiHn9XeALPgC9t83qL6/BAn/hH8vpiwMqHmkADiMWB7EGigOdnQcCR3urj
QhwgDBWjaOnBRKPFRdNKbSTD+rFg/iJpjphS7vuMQwiqjei+LPwGDLE0Qc1ChzbU
4vx4wYTrVHxXlcMGDBrL+YqF2hIuBti4WoTrFUeHeFEv3OUgQMAdRyoVDvteZbY/
BqvIxkr1I0sc6W5wu98NRWkNolK5pBR3K6yU6QYBfwR4DVkjIK9scjxuCGkCGKtr
kXxXKpBiQAA4szFIKr/2Ir9dwOc9jl19wIxA6C6oIvv8Yqm1aoQ3umMH98t9Y1WV
DYDzrGOVWMbV9rRVfgTRG+p315Jm+yrOfsXuzvOQqrHpl6TyUETsvfi0HuaWQvvh
eapXQGOZwu/xo2jDOJ+OxI7FTg0CfAclJGl9WxUg8wo=
`pragma protect end_protected
