// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
atzEn67JZcUI5srYZXsmBix533Nr4gGPuRyXu/tAjM/EBh1doFPEm77KRicx/1ebEAz6SgZtzdEV
w+K5dvsT6amStm6iy8ylJ9i1q/njfjhfBw0F2HWPtgNpVjBbvC3QMnXdTI2KB7zJnHVCQiAL1WhB
SYEhAlZlASUx+84Cdj9qu7p/FTnH/sd8Q1RpIwvGuogMpcMda0zVk2lnA29YjrNBvPyXGMZMBZJ/
0No1TDsI9JSmakFWpWdxEcbsxGBSm44N8Vy95+2RRy4X5hAx2yzrnoHhB68hwrvGjZBdGsGiSvzL
teoPYctL6KfWLLDtUcIkLXxDOnnMnORGmpRHfQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 50016)
3OdwvesahCVDqmhN5kc+4EWimwAgcP+yIzf1lB00MkzA+H9TZNln7hkeb3JDh+//BD0JaZcuPOnI
oFj18Wf+Jpa14q1MZtyCQhvTDiP16KLgMOR6g7vtxkQSX6SamaLxX5oF5LhCd6lvhtCTfDbM/lM9
fZ6d22ZhFzs2OWNILmsoQ/d5tiXc/TmCYaENltFz5MYHbn9iuTWr2juYNu3LlrtM4E0OMemjIfJG
RgysrXHv7KQw3t4yMgnfNcOm9pigxjXQO3I8WFmWmF8DAN5Ykb/mOr5CzhhuhN3QwlY1xi5fs8Ix
ZSKWuuUtNwAY6ikzDYAtOsbaRRhaMpAbsk24pLpxugDqzXb2dBAi9IKGBrsue+fCjQCxfMWXe4+6
w76U9IDpsfRSJH6nhpBWWzkyuE8VZtGR89XErF/v3HYoBMohkCkzbYWQhvb1KdiLIvaYX2HItKnj
7D0TXZ+yGZ0HsKul4R/6rCbTV+oUSSPGjBxJ9xb6qCYVcGyYL3UfktBDH8XJlQcBbb7/+7GsxNhD
fPyR7Nm+LMPU1JjftXpwMMvEEQHHSEVCxSZI7SMS1raGtOZBfSD5vFGKLy2hBFGFLZARSGfu5OB8
NE9EtMNGuxGiiVBtWPKw+h4NSbOPgF7o4qWV0OwiUuQPTrW3+kGj2aEdlPftgg5+2Ww7npJd8Vbe
B+trTD5nfrd61AsbbCuXN14wgXPmElZZjKtWZ5huxEZmnKHKOmD8r7kXt/HOS9GfJkNUmj1heO2J
0tBjVBDlmXXbPYUOIGfRUWTOHdk1rD+tISvs9K3OtXY3WQjgTQCLg+PGfk5GgpT68WQQof+v4Shg
fxJJ6V09qleQfzN60JGrc8vewENkPFsnMLl8IEhBayH4XsH4l9rRacFygLVBO2dcLcAUcNNrZdNJ
enrjG1ZS6JPn7A3t8TVV5sb1n+c2bs6KREmWL2GqCrbHoMxQzTJL+gBxGjFUNU0YMjAVLge04SsG
M3QjjJLUWfz7n4MSG+pqVnPE6XCw0QZbCazCspqYTsf9yvAV0g4Wu7OeDJK+ingSaiRwrw9t/uzE
geSb2i1IrxLCFDka3MM+GtKXoJHfAAin4GPTg7zimLUpG8GGcBS5Ro9c3iUGYrGNVm8N6r6PDHyT
0CgJCx4PVZ4menzG5eW2zowHkPCHI5HQeS+FLV40FplrNvbrVVr+EXkSyHz6A5z+wjIHasoMUl2U
AZondOAT+z4XzknY7AW6RzzHN8duVommo09oh9HVztVjhslTXYEj35ItopcWqZX6K3nlTBUBzmgy
br8Mnmu26E0qsSaDvyHuR0ti+67PkmgbKxFYeHfWLu3WOYsTYztxL/Bh85mU6Re5x34pQAd0FCnI
6nVDMylrxh/cGHmID5dU+2EeJnEOOBaJsOxHbIOssXon8l/CwxttTQdwtGm6gYOCwFhKYowpCTLY
JQT+MMTfd/1r9Di797td4sh/5W15ZyWzLhepDwNvlyRP/os0ozWMve+1JYOs7IYHICeRnx5xgWx4
VA0zFmzfWBnqEismpkyX3p/cb26hc0R3mUHH0d75TDTHJG1eU/VCR0Y3r8QeZv/xVES7yh17RhhC
54gnCjFn+RTGtxwl8Qk8RUBDRZvzDY8oD4NECzIrIPL5EfQQiAYdrcOJt/7jfHsm/RrOF+geBpMf
g8Zr1JIdoJ6xNDFdquZd35E8IlL7Xo91DuVUys7m8KRGE56XbEgOc24/uJMOgvZMxKK/WhdSyhQF
hHr1MLHf7FIwc9LF7KjBibWYeJIY8YuowPpYbZrl4MwDHRFu8TgFExC8Xklngdm5l0eXwJTMn5kx
xjJjSwOFvAy4Wf7AGisPnb15Oz5XvEIP0sUf5mI14aNb+HQYm1kaNnSl4NvJ66b3yk3CjUgxwi5s
1IjdXPKLSS7lguZe3yz5EKCcY2tQtP/D4xwJaOI+iRnrUuQz903ZTZ8Zm+JFUO0KNxN0mhqvYKyC
6Ez7DPbpyNuwc9Cf9csiDyLez7vd41XF77+EBla7b3ZneOtOa2AtyJzfMJ5qnO3E5vy83TgUz9z2
kpN2eqOlzLi+rMTahLB6xD8ttgpbkvrjR3Jz01Z4ZhK7xyMjrAhO0NcPW5oOInOS3YxE49TXUVZP
1SgkUrhG1OrjAYzE4oxbJBg+d5ZoZaYQ2T7Isg5BVXTsaEQHA/Jiw7yt1Eh3iLiPpczeEjendf/9
8vK7DrFA7wAmzLdZuX48z11FFY9/Aap9lbojXL5MmRIRHxR312woVPg4cl2qqWDrsq62TWxKQIZk
/xx4Pi1Xe5xNtnkhmbGoaZae4cC4t5k/aN1Raj6oFHpsiwLxKPUF5MFjIICI57P5mM3QSm+TDXJX
bSY9drD0JZ4CN1BrhJMmJVwTrRQitNc90rkBkiCfFXJq8TdGL4ybyBXyEfEGw6Ybl3/CEJlM1Fi/
7B2PoJhOa+g4LOCUG9TS7mLEvripDSTltCiYirvudOwOX33Y+loRyZEQwdcX5OIgDYty24ReKFR+
lEf2+lyQfvip3EG38h5LwAslQN3seEefRmJwdrRhKx8mEMke2u2lyfWyCT43eVKpn/bQeOdcEXp8
SBUqNVZiTmCxSgPAD93grlVwvqKeKNIxZDPgEt8odYp8i/dF4DCuhBPmymco7/FnzqeLlfHbT9Zl
ShkfKD3iev1oB4yFHvTgTNQzH7bVAwIGe5aynVxWEnF7CZ40HhmuS3ImR7X6+QdYhqZE5me6ST5X
fVIsgiJUAE+4OYAeCkWHR62snAXGxtnVbq3/pC9BAmGetDWJ0S8cDSuSGrLmJJu7uDy40Dp//ye5
nSQT21dVdGVCt0k0TxxrX6SNQjHebgXO1mhFtwF/MZB7V1quFAK4I1fKW54UOY7nm5UXvxgI4gMz
3+GSITaBzVvBDRMQl39ezdmRkzBWCLFvyoarVPl1J18UeT75GpufPSDL62NoNtr6rqpXkze4/y9P
NgSObxPEUe18sXrCshoxKtQvZVFgzMvRA/6MiZd/BHX15sNdVS3h+h+25867QJ3QxLDgCmFl75SO
NcLUomKZaKhJ4y7FUiNlxfePP4ZvI8a6p0gvJmvdjW6FTbJB6KKOhhCw2yN0Ka3xepP6aCmyLWQ1
1P3X2JUcu8v6XeKaVMZ8u3u/5U9XZlKSsYIjLegI1BXZo/RnrdoCAy94s1ij0C+SP7Mhuu4Nvz2i
I8CM84B0mBdJungDEXqYJqOjA7KG9Qaud6UN0DcfhjKCD6FvwUjBsINvat66BrnSopLrgJlJrqsZ
HoFxRe1uf6ceqXfyxOxsg1Q3o+2zGSRB7IUa/leo1C7KEToO0auJV8SVw1VUNPPwWVNpUMqIxyyE
/QYTglhOk83JbtLdaJIu6dz255fLpfB48Akp0ygQiE2KFoKwUbLmwwMdBT4yEKtE6nHQjlDWIRCZ
pTw9fRoSR+FZ+d5+EezMeuWkrYf1DKW892Li3QXFkF/ylpXmCL8K0tXAi5qMuGhwh52EzxgH655K
DSLk8XEh8gMybGJoitNDTll15hXn2JEUhbrYdcWOEimzhoHkno5y4AS3MiBFQaEQovF15bx2ocrl
caNsbia8130pmHaZ8Mq+H7Yyzcb11nttGWmvXbwXGQgsBH8Po4o+rYZqFm5xQCq3KxtJw/oDc9tJ
MKuwXXip7LIGIqz+GmqVX0FduZcyozgGPZLvDUhuPe7fLVu+1ClUUVIUNX6N5aJ0SbWUOdp5EmTh
lqss74pDJ03sNB+gEswtQmYwGb35wlM1BNlEHP2EUFLjvWe1Ao6OFMdzMD+dNqCKl7yLPKcH7vwD
p1wZ3ufliKsa44y19oufpCz+dg2KqHKJumrXvY50DMDgQI8xUL4HUSH+cKFqy09H7Wtu4SChvAiX
yZQJ1/A+XlRZ6cXiMTwkcLnjQL2xjnx5DQrql7TwVl/GHxp6oQyQoetWn9y8Y4u7D4GL1HegdPNZ
yV94ch+6ON4CbnKcCBiZVou4feXW8impE0aCbysoJIe/+xFFtfuv3BPQZV2qJKrRjBVBzcYUyYDv
4ZFUznBZL+5SRXVzMQ8YsUDDQnK1U8/RLr/tN4uCXXISltiWrhCtx38djT5jp2uzaghb3wghf1vf
G/prSyo0x271uhNnleBCFHBH/WEh/z1x/RAarOtT9Rux6aChz/YUrVvBOBinPRztpLUnWp9NDfgv
FRICOKAGSOeHQeVBgM5fghgD7x/FvucBwu+HuTQKSIF4XWNSoQohv8iIEpYyBqhLjFQT+o8LksK4
fBKpTh3HKNfxuiVzKuX+rVdTERCsWebTHlr3obC1JiLBLtSg1BUUOiwpVbcS+q6I+dX3afj8UQOp
8movJ1d/dc9m+Rz4Nsr8hlzcSWaZsr3hXMHq+uZytXUdanyAKc/Bsbew28epAm1CL4ohgpuZnVmQ
o4bL04vyuRaz3JcZ91RZs4rf552N9NGbUPkkURAyGuPbCNlqGU7N28P5ilB8+dvLpjSWhjsT+Y5b
LeowZ0k5e++l6dqiNDexK0DXq0wN+PapXwuoZMq9ggLov1vTAv76hVtxXE7/vCyFmbszBedcowNj
9C4fz9flZM25QxpzXJws3dn9M7Kze/wg/3k1tifjhFoWJxxsLVrt0JqKaPwUM8fw2qt96IouSaKw
zIZSFeSehUb7Mgl2yq8QdX8/uoz7urjSQtNiorCfSuRZDYRzV1x6BQDmObwR/FU6s+Ll99c3T8Ja
9zM3HQX0LXVMOUpb7rUc8ZFUKUsitSrOCD3kNw8v2OsTR21IlS+MAyGDOCv1LQvON6uDYtrmtE8T
MXOcSSAr1ixMYcnsPO8HChoj5O8DkCxkBFFhBSKcIT/IgxyzuPtV9mKXduvknwaCSipKxqy3ow5s
YAXQRXeM/d3HOzvvRGke2RCFvQ57nmyRyFtCYcUqH/FoMZC5rXS/qlbAUY6+SF98Ip5oagE11j78
RFHGTd+rJX5qtoZq56jX9bQDKjn1Js97DJvLa4TH5Rz7n6SwbvfSXh77UuCkzB5DI6ClU2amQ9Ta
JL4VzzB4FdN+jLKvnOk+E+FIGzL1so6YfjEJsDSWj+k4MwmgTb10rPHBbGTk46S1veNv4xxFyeCt
Ixb1jbZX2iVxSig3/cIuEq9086KFdrcJC8EW64vOEYPpuaA34TG3R9NcRC9+QEhmgXjMT4zP154C
ET5WtLdQ+vF+1W3VbGphQHbtBqU6IPLcQX8xFoirNeKJ48GAuaRLzkLGLmnYevYaTSklQXkaqzI4
q8I7+0F3+YSOXju7V79YxbX8Dpbs65M6aKIoUAdaCOM/uEfsPQtqpOhIJbd+jLTOcvy5QIQQ6LL8
ajKeUtwxATNgdzB3L/L41AbFy+x9Y8PZl8KNhv/YsF9hATHiThR2qKofX7wKVcfh1orpt8PDqSw8
D5AwvwUUPK3SY1cgwpDtMpDKo4XNgqgoHnuNM49A5JtmyLpb0+4f9lOIQVB9JH+fcQ7iS9+YSaKb
pyUaxgjMobVLW3xOdMv5EuAIr6APyuvndkZuYh3R9/ctANOLyShpJ2jwEoIvKzfbJMXThR8cpO0J
7OpntJayw4XULPuXtT6/wSqWZJ/1UuwOBxrNT9tXP38mc0jaWBKveDvyRNHYNzF96HJ3OCwt1ty4
ZOO/iwguyN/4KJjsIsilAr6SIInxD4dZW+HlHv2y7fqgT8MEVxP+in6Oou+VFvUAHkg2x5UFVV+g
t89xSFe3UPqb0D7HREmsp0ppKJezt52ZGhldjIAhfmehqQ5dg3zad7I1cNhff3Z+HID9rBbeOasj
XdMipk/ze7cl23jimSnHToU7fYhWrlOukNxacMeJ1ZTbuCzbFlyIcG16fsaiXA+cw8sQe+DoJoBZ
x/zPr40fWW+8bCyhJ+Ookg5L40LejW+WeXmFKhaMVbSZwbjbU+S+j7CCrWDOfZvsA8wRSD6v1u2R
NaETge8R1h7uCZTCpkXwnk9BGB/rcTOOVznztXxOCPjvi19C4Y7fEj4B4/hNgAW073Yo6GM3wa51
vz1Shm+29ffLu4DE+iJqjVUrdgjoDnQ92v4atyGnuUB785yVGi7ACIZtV1fW+Asos2Tkm4qBRwjQ
4LXs0Ae0AZtUWuq47r5iL7arzP36jYJ7XYexuJVxCwV808KKOCQt1Kzxq+0Zsmh1mYZDCI3Mdp4K
1aNmV6c0rHRwjTDkmVgnsf5A/29ZIOfBklFGdNtiXOg0K1y50u3J0jvPgzfPI3LB2EQ643xKtL+A
sICR6QyxcphxU5oiH8lJpctiXYkYKYeNg8vtHRO5enPeioG41NOFI2k2w8Tt1OxP4lWvSj9Spyge
MsUCdu2+D+0MFDgujBK0IJRGVJT25BXC6BrPi7p9ELQoa5olZjZR5gQFtse240fuzF1pDoUX/7Sn
8SPN7QUflkeU29Jh4FYi6EjWeC34cmB/kgeHQhoPkf1GTri6gqb5tVg9SfYJyyFnXczHGK8XSFvV
vhIZ3nnw2oRfTt+XFCokNbyEXjRth2aLgChHrL10JWNv4ZIAemQaAuY2TjkMzo0f43gyWT7KPzLt
k/989eABhk4aC5KHIE6i7/Hnv7HfDVHrryeId+HwI9CQsSXNBjayH+azAbP/cyvHzNvf/ilJOaTI
CMLYWB2x7h6x8obpV1AUy0Si0+YMVuny6nwU4ZM+bIaauCZdIGzyZTDw0Vu4a9GKtNFnCoXMyfOs
Yxvu/6ByO7kGSsDdIWiZ3CQUtJCdp+AnmLDzypAz2fpJ43kbM7PyFS7y9IVBwO1LLDtCrLBIgJCj
PmrRRTkzH8t3nP+rmipxt3ynTXVq5THFnhNkKm806tsm01Pj4Rz+Z2fNSq60VoVUx09sNCBVb+2G
mfIuryZ3D3h2fUfCywxt8AfEvr18l+TcrZvNwQlbS76xQMvygMCVWOTG6rg67Z6GAj93IKdZFjpR
hp7yHJdvKkyhUHtqY4ohLp/yrphb/fXzzwWfoM7VA+TiPbZXjCw3RofE0eu+ecI3Pf17vlikWaN4
V+l/ONo3sIUOV1ZtAFFJfv+q08GmrvsqC77MX3QEjzKpM+WZif6dZRm7q5jbbgjWmsfAiR3TQBnS
m/8FGBucPgX8h8m039ynV0YkH6TO0Mu3NZmxgaikdsYgUtAFZUzZTl/bKR6aLY7ewoZ0TPpe6j4H
t/hfuior/0BjiMJGDLyJ1hchH+ho7h+AwocFOp+QSRhp/QzjQWn0019XKwXgew3lp48GyLWKrPv0
AamBc+QmZDslkZggGzgiNzCRSLXLBz2YCBhaef2U0cuLYisqGyGf/le6Yvv3P9/o8JsxRRsnWyK5
Kyl+Mjf01UUxRm/TlSwF+jegtO2VNJHRjyVmHluYkL030eURjOURFD1LlvTCjdE+CZs01j6D0KvA
N6CJVCCFOX7q9AaxiGkjxkvUtMGI4l31XatnOJPrP7RGqGifjnYxkHE9uvgK7UdWce/qi1uExuMh
os4EGSRc22lj3tODZzllHtaeoKSh909GhqxGwGiprN5HyV/BF3rwqtLdLIp22aK2bKcDCM0BD3oj
4C+9/w5FBrHIgwC7G1mOCtXzTZmfCbGYeS+sRzEQ4ufg/zl7XW204CKjNXgjOJdVi1fzxQEzyuL7
r1QkI01MKxsjvayiBYBgJRHNOPYK+gyu1tHdQSg+m8h7eih673Fa3LO7GgatzfhOC4yt7MbLqRuq
0AwVjhTouOtNDtouSg1BEkgfUEQCg3W3q3z2YMXbSVROjEixyJBf0WwN0+JB1EFA0FONDu7UnlNk
7tlYBSXS3Zh2prB3qrK4gehvgeIPkjVChtb5/CWZwVHSt9JGrRH9mNQkBAgj2/dnvqamNBEksVJx
ty8nof43jIz3kReNu/ZYXSBUDpB/QAuRYrjGE4Qy69hKpfvayo2q1AimKE7K5D/vHrHn2PbgDrDF
l+xqWAA/eSFW2xEtZlHzPnzhzSGB3sySON+SuzDC3iHnUJ+oT/43Lp1azd1Q8mxujKPi5GcqIqr9
C4CLiuEKtyD7XDYg0CFpPC8qMpb8KlCKq3K+5JD3AxCZcvAkUBjgInIqF9BOP3U5NOYuM+/6LcOi
teC/HbpPyQvA3Coqcin+rmXrfAoZSiwpGB4JLfm6pI3cPMZn2bhgnFOT/cSM0cIkggQlSSNVk9Xc
0mrwOCsAMY/PkFbK2pXPKSRHSREu8yjwZm57oAPVtJt9EnLPuEP3qaxzbkdPThug04cdxrX20+2f
515jqr/0OP8Km4a1XWzbHIhmcofzHW2/g7WmsUSCc+ISMEiwL57P4LjOJ/JcnLOKC+xiIti9uAGu
fbbtmmhGy93HtyQdeHHh98xLUoycZR+a5S54qExGis0oNu8RcDQkj56XBZ7WCOFP+mGoss3klk91
Dwqyu44NjLZeouteNAb9mcR8Zb2aeyOx0AyTrZ7OQmGk04DPR6Kc4ps8DuT6FlJDIYscYAwmJtyc
9HiBQVbmn29JyiVzRraVHWLRIZ8wei6mpMG7rIAptArIEB4CoBzUQeI0Cly3MF3EwhgZF7d35z6x
uR3GSZxRJ+rcX5xh9+MnxZ+fld5AWQOr2IAdBQAFUxfMoJHDwDpIdKmxafuIENYjibY4Kjj1ugJQ
8Bd989lzQ47q8W8eKTK2a/TtU1bf6U6R4Rk/E2lujdhK2kegdNPEFvLEwZJnKq9b+ZqBhYK0hkJ0
byq2yb6es2e+AdIL6YC71Ih1ht8NH3gGNBxYwo6etm/sXu9MIuzCYzVujEWlTxjEikvX7uG7+RLr
TKEokgbUVKw4+xxmc0DqK3nlBLgb4xMN9xyP+vC+EnRmXEMaJkLgCY3ayY1fJTkomER2RMV79i2P
Lp9Vjer40rqXigB9BD+gOMFj/Bx3ivhkJNys1IhZ6nocm0JLQxRtPY4mvBG/knfL4oiAemQsZ7/H
V6EAiszDoDM4q84TmfR5t5zllM++CJgHVykxCwnoSXRjGj1KJ/Ay7UZ7C4jYbLK2O0WJ8Y+PIbhP
barMY265h1+k4+p5dSly7pOiNa1FyRoxeVwrMyB52z1F5XM1hfqoXR5kO5tPRqx97qjFoq285Sj6
MO2GIut5oUcT2NN9RrQ2TUzxTHRyo6ORQDMw1VOtxuEPHv6ITyy1jDpPrfv8WQLEnQCDpYX7cUVD
46FiBI+0SsLaZhqUjnv2o2/UUZ2eQnCjzZDcQ2btDYwlJQOcdvsfBZq7mNpGzEjrIDHK9HOowxea
8cgpW/77XwnO9vvZ38xg7Wv+M+32W8O0q1VPwz1MMcOayhWi5HBg87nzCrGJ6uHvAXubdluZwXQP
W9OjMXGz+c4x8mHlM6BkGIrgN8s2Zca6KOIFCZZcqPJIaQGn8gJer8xIKgfQGsdMaaIFrJ1ekmJO
0WEp6WNJ2cjMKsq6767TTuepLE7UsKhVUDlyJLZrmQAOadITVqR1L6wD7NzuyAMjOnEZj4fMgtNb
7F6w2bYGUbBZXG3Rke7EMO0kdgaP2nUQWrgoMN3xlumOx+yP/MiyTEeeHQp2WfbNWVkfblJF0v/A
cVkEXN3tAs8mlSU20qvki7RPP8RF58HixJy7qbe3K87kkZEGBQC5Lvie+VK6ddx+Ngz9IwfdZel0
6TCoSsrzS/V9MjBNDo+X4QGDRl4vVoft8/peb63ZwxAE5CjK8oDVeNzvRqYSEc8RdaSDV8HV+BBH
Wz1g/jxCOHlqBYvzGoA9OQFp3t5s+N9/lGFRKXGohPC1gLXfMTjNBKwYn03B+Cc1wY7U9emamZc+
oF6J5AbRRdXtfTe8PLMK8gLV9ix3JZ9/Zo3jwOc+Gq9W3syTs4fIc5zzdhMtYAfjQnedExWc+Fa7
ejccW4RBCsEyy/8MLzS/vomH6vqwo+AZdT00Vb7SFPly4z8+QCPdt0rANHJJkR6J8xg5Q9AeVKOl
p8AWPNL0hWr6MYT7aCo3np/Uk7Oxc5LZewPl1nvoCz5gwVvpCFh6YNt22iH8Ly1sKQKi7JN0M8mM
OAnnDJBokGM3OW+7XDXyTGdyLJadTuB5Xx4rqxuG578SU3Y87yway1iuPvcTZwGnL152TAI18fMn
uwcIKFGq9SW6N/DQ24MHmb/0C61YbQkAzFUX4gPBrBxNhd/YNP/CqzpA7rRf43oGs+WyPoX7Da6P
bSMp2ioFZd58JCbaN/ndZ8r0Ibcq71a8739NwX7lJZZwATTdX362+9CV6HPYmPrFLV73F7zmPeJr
QFIgopkKX0psrXatBFykJXgoIaKMBcZPGKEXBf/Mhgw3cXA8LWK0N7eGROEcDnSkDYCc+pjHqW7J
kJzaoUKuAAnlsNz8yay3B31zf4hJf/ysJZEM5BqAJ7NoWE6ZESa7VyQyZKaoC1fw4/FOu3lsSCNw
ek/nOCJ3jXBYxaNS+00BqW56m3+n3lDnUszQtnaxkgSnUdIfQWM4wh7jysR4CUMs5KCUtnHa7O5h
PrGHvzpKpn35ZxcWdB+VINuERT5SCZasHfbazSQzvMAP7xL9ypPopY4eXXPIVYmmzEm1zNUFZTvj
Ucm2+fjjsyIt4w0QSVTx+D6QV8xU8kJRCx9uXi4AlhOo9KXov9HmdAcyZy7wxwwm7w3A+/V9BaRS
YHQobOZ8SsHuLBAVg88Jwj8x9Nnl2RajKaSk2dElzVuGd0MGB9JjFttE5/nl4tpLTp5K4Z7FN9qC
8GgBntgrcI/qvIUuKRdHOlE0TETyX1Mz5F58U1Ds+m2yd/aXlurOn1PPmDQi9zGtwopWRP1ApfeY
m4PnUYycYf9tSavp0usdwhWZUz20EI8O3sCN+loPfk59+GgCxx0UxPkPypInoeWgDph0cwfHvQDo
FW112dSyET69By9CT3kqXCOZjW4RpD9pllfniG+T7mYIwjjU3xfI+HnFsPk1pnyNauCgOqUNL9NG
X88Yrk1rqoYwGxMaNlg536WQ2f2E7nVH87kMtiQPkimvQS/q5c9Pat6E6LmQuZeq3INRtO+G3kFB
q61M0fKC0hFazgadBCXgP3XWrvnWtV2FNpgURJNWDJ0shdR5rt2ujtl9SrTNzE6eMdqWNJje4IBB
pc2uCiUKfrvdmZ+yS9eQ2YHxZfAxahs3K+Qr2HDo6FkZj0vNih/i8TYGsToZzGyB4caNkwfv9gfU
VftV8pjlIJtNg0deAXxam9E1+MoxtdAR1vvA3nKgbxNluNhGCYgOFVNQF133Zp3/ntQ3YTS5afGW
tYvlcSXEyjDo1reewCBRdvxYL9ffWHRI297wHiSO6kKIGLsMO02gz/3XlFQmLqt0lEEFs1BFdoPB
4rlkP8+nytKSHl9h1WfCVWfrJoc1u2vN7lUr22NrTTa6j+CLnS0IHTioTJOoWtLmtu4Z1BXhwrw4
OAFydXpfxvQPeRdCrZdD44YYRJOxxq1nPHEQcvr3o0yURZDw8bpu8ZejrbdnW15xo0nzGgQs46jT
ixErqOehaD21fhUPoydhgogx7y6cf3Oa+7zzfFnVkLMtxbjhS7rPTxNU91pGuLKLdnQimXfvUhlH
ypS4mbULArt/V9sA170tY4CawQWcc8tZH72O0cMgjQs10/FWaMBSWAvZ2JYmaG2Fzf2twfJ36uOO
2X9SL/+ehQeNyaT1e1JfNgfMd8tY3wLyJc1g3oimsSbUBcrTaThfh2dp3IQS6a0cVJQcYyVgPruw
yfc8D/N4vv+57ortIStUbMJ2hkhPdLb1o7BZscrzkXn/VsX0bMpwTJWkrR6WuUioEA1vyBaG82aO
1ofVC9jW0tcYcvZ9QCmHPZa0Rd8vGxO3dfUeSxoCvUrM39jq8t94G9XLD8g3Kwx8vMYSgOF7U5em
y1t9bNoP1S+aK9p0ENgfcw0YhVe6qmwXTEASPN2xPwQ9S8pSVn61v59R9HpFWhTCChFvrDaNH14V
zzoFKweWw5q1nr7CJ0MHCFLXtl9kzH7sWZXUx/PVzIBIkG1eiIsYkz4zzS/WmzMJfRcsEKS12byM
MDzP7zQFh2N0jQsZYFQVhrZB5havLyF/YamQTW5veujXwA2rZQTZU8UolVCUE2EPYDD3XcvMcITI
GC1qGYX014jeEsRusaNNSpIlBo5GaW3jLvJLqMTi+pL5kDXRSwZv7Ja05cxLhDeR+yUlqHLKwXeI
SWdWhtjqOw0HrTCDml6jF5J3f9gDM2KReoCb4BJyCEa1EG54JK/H0wJBc5SjTQwJi2Yc7gmLwp2S
or1bCQJoDt2Syq/pKxArfXOIkYLfClF0oaPlmlTTN8kvKICnEd5DZn7zoqgpPgwymw8kChQPGdBN
FtuaKN4P7MywCTNuXhc3mqjfMOcMbsXHAtjO7l0UUL959DqYh79eSB2yb4qoxyCBMNwlHF6+Z6lu
8hUCtudWrr+a0r3lvsb4y22FhE74f7dgntfLtojB3U/RZ85NeNQ22fddBU/QJAJ8QcUfNB+RXNUi
qIx/Bc6MmMDMVN+TcL8rTDrxu+eZOlJ9tVcxQ8sx38nnfujM+1pIVTRE7jgERPrYyXyl5HPwqa86
fgPucWn1Swz4BLTsXYS64lx6r9SlvyR+G6D4EmKETWrCuktpvNbo8lz4qt/dxQeuIggMZSNEXwjq
Rx2EXwR9f3I7F4CVxMnk5wexD969GPSoR2jSR/h0k/mN03d8HIpMf+a26t4Vk4a8y3rBHWiLra0I
G234wkaBNtRXSbVAO7eI6zIxyhhzEXSQ1n3siPGc3c28IxvJHYqozjj5Bg29jEp3VQSKJoy6ZsLI
bSU/xHZXnXxn1ZHumYiMxoPxfwDMMlf4DQLCWBM3DffbPmPzZ9BZScOmYmXsCy+2ejVSiTpmqPzn
K6f14abXwBPkO6DNzUsTGI2xuJSdo3oqcNl6CRZBztr/eCKUJbsULSJvxf6hALu9+Hg0weelRJbG
x4xS1oq6i3ldv+G8DtNkqHihYb3Nof0u5Q/t1oq3un+r1qnJsF02Rl735h2Fy+SXNXe2IKrrYOZE
BKQrEg96FlPPSrCP0iPAt/9OnlctU9dxQiA/EfLwN+PH4KaoK5pJZtEXCWPSxMpBBwvmnJwN8xcj
ebF+SuHnglp/R94QSeHTzso8yImHrUIB5oQMTUvAFjjbJL90uWqGatQNDxE0h5heuUsktckpyR4Y
enCmNdTvjvuLIhnd02dC1Uz5Wt6Mm0YSxXue1rD5GOTV+iffffLXY+pOXrWjUGtD1XLKj1mNgMVZ
RIfadAC+waqu5bE0e5aMaXWhXvOYIJ3x6/FyAR/EleqMPnYNa9MSaKvD8B8W2NKV2UMjO27ejqDP
32XBLxReBDT1bX3gzG3hS5pO3DLwiJTIU/2YHbwIWvS1Ru+h+yBstcncX3dmoWQ9lNZCRrsnGeW7
d+bPJ5hX8EK3sy2ppsyZKX/Qq2VNSSntwsQUXK7rkloRXIRQFf3D1sPJOolELdB4BpYabNXYUprv
FpZmbO6zZpS8yknymRYklsLTYhFnM/3s+936TsoDv4V62XLaNevOV6W99IqH0rgyRtnv4cKVdL2F
eWCLaVj6iJYaSSPPBLV/fDoOVv2q4FrCniBJo4RbINMzeyVrYlP/2BueY9FqtIjXlLStuoc03G1p
+T7lPKPeoUZwjT4Y6VVBJ5SOp3Dji4qnEnXNpFUGpuMx3PJHYxDgeXkEig/xvK2KQF/lUhW5JQlD
WAGZ4xBIL2yjb85pdVfmZIS/1077UlsNPltHlet6QhNS+FzLjZtGaFzQBbwkxaSK6+N2nlWHA++6
Z3JT/EMhXgeGt0EpqZdyVmfuba9JgmT0Y2RMeHWNiexdYG3iZ8Yh60Y5pTSSKYVHQsMXwzSi7djD
oHzwP66OTn15ne5RePSEdQC2d+2RUoi3XQHfhFLfVM595H45ToZtbsSrkjbFf/4PiPZQYEBQ5yYe
zeVtQ8a8xVncollSxG8nbsDLRTvPQwC7xXgj//sl04mr2lnFK0z7jbeOVDO+CmV2bIiAaacuO2y/
eeHX7SKuJLtb0DtOitsM9U0lpoyuTEDCn0Oq3A5xKNmxz87ZQFgOi4RQOB/I99kR1rmEUiYtd2R2
6UcXh5+wXtBzvw8NwBIpJcTht1iEz+Lv2jmXXwjZv4py5m9uFtuzGODB9CH/yclh41xuyf3ELvcX
GO9MTu09jRk08YVkiKYNLzUt5SisYWw7qv7lce55Jx542AnFt7J+bH8SlW5Bush6JJ5sExO7xYom
ec6i7XNQpQSNpTX8wuUsfwbMdM+LHRtN5TQDq4SrxpIOGF3DtqjpZqkBhuJg7diZ7d3D2O7Eink9
cF3zTHfWXqh2VEhk3o7jHyOkVY9Wmq3qhyerCmSoW97duu29VzeSx6TCn1hUfkcFf0MW4dHjaQM5
uQgzBLywhFkQgj13SeHuCEqK3iDR2Kp9gqvDKolHFhz3WpmXdwcxlDivAcG21ccBzr2rgB2jCzKZ
sMTpZbWFuDvTRmwyE8VGsXF7cGjPawMc5UWd0Lmtx2klJmi5JytZeDVdQjryaucVUrc89/jnj8Cq
qsd/cwgmRDEdj9Pa+O9xsimXIbi0PnWadcoTTGm6OVgIuJG8tvmus3rMlZthRBezpPufhxa0GSxE
McnHSEJtqkjDyY1KoF5wd6RT42Y3qT39co/wY0n7Vh6pektslGErJWTrBrg1qAfPoEeQyrr1khLO
Ny+QK2tqLQtqisP4L0Ony3oFKWKGD3cTH1FqMQWxlkMEMXHbYUgxkSYZKnb4XvTteURybI1/93mp
eSIhcxSNdG3kLIJttdCy5X1gKenwvi4c+/QT9oURjFe/UnrHK6yYTzUr1+rEiIb8pDxaEANVD2Li
xSVFagUt4oH6x8aDPytg9kgAVzosUo4T+bQrxl6XbVx2Yw6agAix6VJFmdHfqBOeXZVpfHBNi95U
T4YmRgBdkgCRzZB/xjjkFKtIfFM5DZpetUIu5ixJvdBIremh8MAQDOdUJFrGWqQNy9bZYmZ/F7XM
+Mi+FzA1IoVmtZMbHkMp1OI/Hz2XbzWt8NEUfcwaZAGbnkm0svIaCCniVSz3HxqPNDI3GGF3EyrY
c/aAvzBNIMFcaQzEl3S7DfseaRbISUA8cwbEewH2FsgIITODrmY5bLL+CuBndZHZVl/np5tYBq+4
uCBxKGwI/vQ/B3jw4BDLeL4BfYtdYMs7M2PddOrLX4QCCN/i8lftRKYl5WkxvfkndJBjvDDFCDo6
QqZ38ng6TV6Y6eXOqevs8uc1vY31uoEu+2hS+FgcYqDfZuM1oX0JSYuD1FZWEhUQPKDkUWVABvGy
4QxWyzEWtWUIjsQcdmG3dWmxs+8iNXhMrLMDgp3geEEP7PZXuGd4WKGzTr38qzRmcgfowGumNO8t
RB2oKsCCn7TbRVQcIRHEel1cPCMEzKIi2yqMLgm6C8TSp95vkiho4ca9f3u9f5uR3HcXLbIBw3fF
MEjo3uScOlJ1L9B7Iog5ld/AmvLNnNopvXIH1IxkoAH3nAXBBjYJ4zx3VgNwsMJeQu6ULbscHGFW
OUrIvthJBKv/tN54uONwhsn7dO7ocJ2r0M1vyjo2VhbrZTQscUsgIoOev2vWymntc/ShdTOf8aMp
xg6ODnfIc+GC2uERhCa3NwsLxphePp/0yQGtg6pCSdkYJvKV9SXfVntPQenegeDgOHtS5kubzqzY
YLd/t0HrHqxDVTems4EqtMnqjsb8zrQFoqhNL9w81OG2fJYk2M+u4WC3/tOpq4ooGrnyMBa1ugOm
3nkxA3GW/AxF1YJgiGdIYmUDddrQKmnc+OMkSxXbrR3Ni/3cywCbTmb+GxE3KyYGx7FwyHe99ZQW
1tzK8aVPdCp/DCqDytBsXziDQy3v/E7etndWL3XT+1MlSA/hmBSjqmSpGTSEuD4PyoHqXPXAEue3
f8It4o6fAYIFSj8Uauko0Y+OwiWzPO/phNNylNhWg1SwioClDeO3vYENVk7ElfdSbV+Vv7liShUz
8nQAnICJMgfJ+Qkzww31P++5xNPfvAU4xA2J8BMfKyXpmnBh28nlIQ8C/9eBy5gla5lNeyAt10+S
U0GO0lFshvMb6ZfW5G7+lHuV85ox+5c6WQWJQD/BLHMw77VAYysiXJGwbOJzbO3cO58hjBHxFDmn
roB5lYYP5pB3viEu3l8eSV8oP9B3/cFi3kK+jKoL8UBaKQxERDleSwvQFh+dZeEpMPHjkESX79aU
MWuVrQJ9G/aDSbFExQe5x8lrAfi0lJmwbaaQkTG5C7n1j+Li9dKqQzKRmbYBKg0ahhSAafmbqhkQ
Bb0mGG6KzCt+bZj1jTrfTRVE6fVHbFNsPRCmMeQmVbZxANxmtnBatRmQI4k+YzQLMa7wmVj6ZpVI
LN8gy4iSOoGEqRNdgw/YGeNtzRzRCQU8apkWvjNl0hHwG0t+1urehtLBOFpdhUw0MgOX+VnA9u7O
+dlJ5rWycH/fJlcVYNB3GAiDYP7Z+nx8X3fgTRA8O2RfK5guxBZX77Ccf41iJp+L6DK4nmrej2Hz
l7mQIprgetO+PgznLzS4RHyX1PC+IAqVfZ/sUE1Db3WFDnQcbDjsw4BkSx+VHyfsoCHN3Fkn3TYs
KKAl3pVx3iGmUCmOWO6bkw3OjwD7O9Sm6Dw21dPnoM/xa7ghsMw3ULQJTiZjvAI5gzIam8CeeOU9
13P+WUSkuejRFN78xFudwvSPaevj8e48V8xt8iu0J6WByH7f8SZigN7JOOa6UchUYEc5Rm+WHK0s
y2zOMHWv1iKG9ENomtfredKCl3HfGFJSaFvQZ8xF2kYbxZfDkBJqv3/bACkVgbzwF5VCnOcQLcFg
U3LmCkOWkrfXq0yQYvmO20aLrrcSTTK0/V8clVdsKnmGxWoFIVhl+TAw/KVICXJXpH93lYE7jzdf
fuOAX/a+caqdsRUN+IoG09Dhpu9WuyiV/UYJ+/oL7dizsBgD4UXBeAbC9UiCUEA4nbrA6ZdQxbmD
RW21FGR2o0z6J7vTAmg1QXvdrYkQZ2u/gzq1Sm+bYmD1nXO9rXmFzpxmLcUzbxP+31uteQc2jl1y
41cE7PBl/SYulOr3RX1r5nnZNurtv+ztiAeOWrYLJxkG8Haddsnr/wi4JYOxCWu8ArXkeiaw3TRm
VaU7tJFDG3Xiyd7dHgAh0MMmkCHuvr2hUS8nxNxOujvQ+iINRk7KPUUQcLx18mFKuLi7qicf6w12
CUFaTM0FsNRUY/ORIz7MQLQdh6tjYOqDB3FhK8xgf+KW1jrdC4zN1HoXPZ5z3CXVk/IpFYDW7wHS
VvavLTGWx9Sekn/Zf5JsSHeaoKrVhrMnkNBsfu74APoe40KeJS5bUYHO797VWLyIzR9llNzbqm83
vPopwcaVToIR1hMV/eFk5/xYN5XmzpRcGdxtTZhDvG3ngVExhm3fWEYCvkR1IQOtLvu+JVyi8FXe
18p4S5jDdPfMOmhR3aFveLDmPArU17VOu8OeT/HFJj+e5y1Vcx+WClkJRDJwKgFzMqqjC13fLLWo
FixHu5IrtjvsGQYxtuTmBqVprfTSgBQT62Pba8Y6QV6Baxb2XhCNxWDnj9xlRphJSv4eeP4aPLFW
cr2AtKjcKNF3N3HWlEwtdYG+wBt1da6JbnY2jR0mJh4TkaAbM0U3Ee05ChC/arIEzJC1jh3onVGK
cjtzQNWL1VxdYijlQwys7SueSr5VUOhtTL7uRDSrZOjy4QR7ffkMCIvn9dav/bSb6umm+esKx+vZ
i79xmsGeiRuI0aVQ4N4Q0/5RttcRHqXff0qVsxQIkqSezvN+5RXv+FTv4qnwH8Bb33c38KV/dKU9
EN35Wq0GFISXMnxguqx+YQglimHL5x2scobcPIW3uFjOfOFzbUU01jvvzl6/5qzJyztP2/tXOMiv
F6sr+V/OWYFaBbqY/3ItldbI8Kum5loNyjv4Lq4rCm6Mk1srnCSB1MDa/UWZKtKKAI1ZlsU+/Bm7
aaH8VH9v/9s0AJWpfDkrolgftPI05sIv2/SVgYDLmBFYntNGFJLHF0nmsXzSkIaAuIbhV2N/CUH2
6399eyFhy/BKnu7N875r4J9thkbV29F0iIDhOzy18Umk4+fSbtKbowrW4N420KXu+ahQ3iQYiExK
jAUvPy7pceozaTrnaJd+dbOCu7p3oQek+XdVIiGvFq877KHIP4nAdJSYDGb1QkLMcpqESV5y7aEn
5Kx1f49CUoyjgN5QPhdaff2xnvwL2Bzuz3OZpGFqGIXcIhkqXj5v7B/EQ5H5ic5HrGi03wdNPpNt
T2YJMn5ZddouXqDPKHDLkd8MCt59aDmL25AKrbBS69WCFDEioHASB1Bd9rHizjeNoX5NOnOwYQTV
X0jbv+6z89FGpoaQG8YBsJeyY6/WHzYLfsvljrSVgZavmHdEpVmNN6SMlCDDtgnn/3E8QoABut3h
LCs5JxiCOufbb9scsZcMmWy9y+FhBayHXhUYvb2b50+r3mZV3zWjnrjNS6MEnpBdo6jst/NZ77xt
FJvFr9ZUVoZZ4Q64H0BxhHRSVtgyB+uMLmdl5oEq3TBvSBVFBYezkK3smPfUYPzFr9Eu72GydXBN
jM/Em/vhlH5MrXjy9uZOKXB4uvQTcD+HzXiD0tdRCPeWz3/MitjEIXwvPjUp4w9RhDFsQsMTdV9G
CHlw+lHrCiCdtcjdNeYHgYoArOB7C/+uclE+U8ZX9xWVKt/w7A/1eFPCQeZYwj4cMUcxgFVZ8HS4
7/wc10hGEpbhiJpF9yg73n/1t+kuV6wqs/ElBPTus8v7idXkPrSI8qBNYpapKfSdQTKXk4NXZIwh
yINfX5Nw5LuZ/3ulyqSYxFV8tr6gzeeXtVOJEXsNg82HaB1vwifHoO+zdi0KulPjeXKKwfBR88gC
010e+U4eYgiZfFaTnFoD3dhf0XcfvboDhL9KEz6L/zKuwOaCu17Iz5GN6FvRmWSd9l85bC45aMLo
QIVdsZplZO6DkhruOT7Oa7me720Dlfpantr1FcIsqW9dXVY8uR9BfBP4FekdpGOZbRO0f9JJRpn7
x1WpHpBKnk8CqhlGIYGEbWK7YaCphgcapZ6+jIUvoEyzM/qQ1T5yFonXY3N8E5+XmFMubDrcdtVE
c10dagCg9G5qgTvcN2FHYdSUyB2ENK9KqPOTuqF6TULFaG4G6rniGOqbn6grmrNA10EemN1Q50++
UQBVrFm6tosHWOCLmLTrUmz9QdFfjvMSfmghyLDt12mvtuaQTXETIBMSNDW6vpOKK/pqE/L3Wz22
7gZI8l5fmXMS1PKpRLzCeMy5ReSL6/SynRLZpMnc3LJo1ZW3a++K1nhIQagMsC6R63wFx4UTOmMs
SvRWFnvkCzMbJ5f0jTdVLivCnh4mvyJTAzTA5UUePa5vxgNy7M7dMTDRCMXx5AO2Fjuhj6EVzlhw
cvi/Fp7j+89gNFCT9a20DLOOsO6HNvB6b8O3o3ypG1h+V04oRbWW/0oyZmbKfEj1ODIJMHGXmnPN
RVDT2RHoCzvN4bbEC+6E05nwaCBJRMT7MiBW7Yo5itVSNEof4hno+KY0P6PZ/eT3aNry5m8II1tc
ay8APAm8LnJ0XXfPUo22RTgItbuzBFZuFsydyAf3RT3WOAvxW/0tu89Z43mPyA00EVVRCDeEHaW5
Qzr95DsVN54nl80H4xiigb0Vk0JX57WddKrfTotYfF3q4qPJCvZ38pu7lvOe2iZY1qriACwun9cR
IYxVttSKMrX0A4CZzyV8Spbmg/LZz7TVooHBB4ol2gZxgCjwUPGDihPDFnicFCROoWHVQkV5Tf0X
SRbjv7x418r/HB0nQg/O6zI8Rm5Z5MxBVsQajAoT4QBpbbI5TRAkBOzuqMoENHrr1uuQusmFK6Na
f3WZHwHXStWbVYcLcnyv2HjUqdW1Kr/G3TcUlQHnooDlqP8LSAolJBSvm3QeLnrYhNfh0EwWIM0B
y3EusJks93dgoQIoFB1r/zS6zAyc7ECIkZcVfmIZsTvwckp16aYXSU5AnEWwQvPx43fqL8YSvQ3/
sve6HJPFE2mkSwqIqGKtJcWj7Dp8l5PWJhPEtrmTc2KbRdZey7++AbkTwDEL8drw+0J/9ZKoscoC
tECYco8qKIwXpa8V6H6ujjONYqCtlvX326QYIFFNJT3jLKYgFk6J+p8n2eyNJm4D2AS8dALRkNwZ
lHP4lNBpkDrHKLxIfYty0kXGG74EyuIiGpPs861zO12HNpNvxTK5/j8SifP423KLIYbceoISiDcY
gbKvF9AYSriPNgPWM1rJqicQVQ5ZqftCK0anILJXCPkIT2te0tTKHVWmp0QtkWsF5CFc/ACThppU
9z0n8JxvD0ubNiqYn2aHNNE4RrfhWS+hPKmc2ySQPYXeZTimAOm7YOHkGK28JC4bOHJ2Kzp+xzJL
WWQX4bWMt3KixBrqKhSg8Mn9v5A++EGzfZuu4+X366fkSKNnm+1GO0mSnA5Z2rFVqY3e6AqQESbQ
Kyub3FTqst5vk7RrssNmXEp6KXVz/GO7wTw5gr+/t3NHmvn7XFD1YWFhjXT3D4l5RdKcWZTowcZV
bzEUxKe9xjI/f2hoJL7vqaC2MBgh1XqoCXph7b1O+Z45wAgWynRgorv3WbdijGOOsIJF52l3TW7r
G8U/ILhAJy2UG5eJX+YjPy+78vWcZxyDozPKZMCBxnKOjAVQx3f6rB8KLvyOcVWBmwYF5NHvWBlI
Ua67lTP+PsNu326CMaFm47ic4bzRcbebp+VC129Aa6V8aGUZD3aWlDba+eWoR/o3XzwKqRF8NT7+
gMyEM8h2q98ypz/Kbu2cXJBOSKwNhjIRtfs3PTJ6xFdhaNDBdeScEXzF61ZNImCyt2JmM6Y03ujn
Z38Oy0SVHfSZdVz/fFnHLWQg8pLfBWo3Uli0BlQVNegzsN0yDndkTEnK9gKAx+TG5pDwbxAaW5bO
AOxwZ5CZamYgwypMIlbLZWnJrq6M3DSKzRmU50KRt9e3nBg4dCVllRR1hY7zbfyDiN0zlDuF1HGy
kSEl8n2Gfn5coV9XNfGW1wxVg6TAy5ZPophIUmqJ5tnCxbeduXVmLpQCBesgH8z2AVOFGu32ZUY9
YjKMu+PB94Wpz9RlZiiBGnz1UrrLg6eBGqXWQyuBRGuDl0QRsKAUeCNLPPpFyXLgew31H8ukmRY6
xgpuuDUb2WA44HbxZHkjnchGnUeqS+8aNd0luwaMIWEfHFOQLpVKPm66IMt5pJyDOcXvo+zX5CLd
jnl7FeSCkU0yhadxOG9QCTVX56NHEAV2BXM3krRz8E4wgzqCUKxo1wo0e19fj8GQm+1Mmk4t4EMI
zOlyz2jB8Rs9jUv6ojb7Wc9cExQ7oD8cBB7rbLSbtCvOsVZBQb4mz18css27zFqd1cBrTXFvo1SG
1inTlB6pptX+bpISSpTJmxJl4vlFQj1gV4K2AuoWppmgW31XZ9IocqKDvUD5wJ5xlkeLA3NSEW9N
XqgvXLYXqSCYORTTvPDAyq7Zs2n8+JjREwsozNmo0yrFTMfnsWaH8p8RgyrQyuSpej3Q3tnY9vvl
mSrjQyDGiaRi6CM9sgtD8HhSsKQgpDJH7P/5cGWhpc7LpP+EioTmCHnD3170DHL8+aEu3ZG6pgAA
LsZNbciP6U6ZsCCZEGzHrOSJ552YttOJW+AG2R70cbcOruLLmAprMiqPLyo2VmbYtotr1kwGamvD
eLcs5cS7uN5Mktp4vEayqtaZNCi9ByDgBpZjo7f8kK1HZAoGAjcP5DK26oCeboIgumWA6A0DjkZi
ZtLZROwFkXkLQApPPM3PDR3tqioxdaHrB3j0o8JQaMrUaYzlkL7cKYN8kTXsqPv3dJn/oMRkWkJu
IBaCGzqaWdxSy7OjzQkHhYwcl7vdOYbw99qyOsRo3ZoeoHN7NNSwf0QbAeWeNgvxul7kIjijlPLn
tsyWmo2eY5jtzlSGXvnC2SWl632RpHBpmCKbaBLUrcfWBzlgbc9yJHhLX66EdDM/dN+sn1eqtpzr
3xxUIPon4rtNRoXTVlEOTNOwlEsPn0Ap2us+/6+od9BD78OYptXqVL5avLLJvTtYUOtopkXwiQsC
GTLlQ1pt6eIN2ZIzEzKeOQclAu4eL6Kfd+C8R6T9t1Gl60Bs9XqPP5piN743FXzNhFGLkPCVaC3D
gRCN5bHZhrwT2wUROyGgVfurIgBRErbLr55pQGq3TMwPZUlDxdOfNBixiAd4kvuUPOZdcNF89vWg
e00meA5GYSREdH6Au//PX4fgHJnFUltVSuTqeH64EIjgUbuJv4ijevKW4N4Lr/kRWGOyats3hm8V
3F278BIQ3QLBfr6aSSa/IJCB/02TcsXbSGZFpmo2YlaOafrNFAWVE3+Az82hrqA1D/A4iSp0yqeL
AZAJtpZqD0pNdnW9cz+vnLg/y6LKXqZVZ2FOqMFPVoh8uJvCeEFYqMNnWLHTf6/19Fdf8/RPOWPj
C05meQWM4rSB8sMjjGxiDbXIcZJaSV/ksy+JPlSyohxSercGsZPhcx6wT5DcZs1FZBh+2AWMkRHl
wZVdCSbXW6uNAWy8M8Ab1n/NMzxUaLlXe6wTY8GGNQMZJ6mG7quxjIBeSDzw7abBL6urpuEatnJG
AZr/O3e8iXuMviuLabD2D5jvAyAkeFNWikzXzn1YkBeUOw0C3m1MEHyKUS6RfWVrdEd7M0AqCa2K
UqLlMghYQkOImT59QMz1+f+uWfZMRWr0iNgEIujOMxa307cbW+JS0oCM8GDblAQqd3LPn/sw9HZ7
pNViVOP+isX/c5qzgz8BKZn1pyv1thBGkhVXulQDble6JSlyqntLqJQuZWZUzONwRQvn2nGXbcsy
ZcHDIqgb+NoMi/BcU3bruu+pZJwXt4WFXnL4lRa6NZeDx6k9IlDipEGRxuA99tC194LW6ptbrzkg
2MdxNLkGVcK0NmpBEdDTQijmMoI2tuDJG1JUO1QEGxpdVMfhCndGkvPjDKcbBa6u3WVHc4sDlCpt
odpAwAbOROxrmeLYAn6oLhjtDKFqPQehi3Yft8YepAHkEuSYOtLUipcXPSFZrd9ODbuka6jH2dPC
qczkIU9t1S7F/DKNDCU43EOmsOOHklQq7J/XqLvQ/qa5engC3zqTpokIenMMhMb5bLKMxjNQljOy
7nXfffhicxxpq79EJz+8kGWOhpK6ueN6JL9vbU+O09cBen2aBw0LOTsfLxWlqZh83vDCO/FwMoEV
w335a9YgHVV9tKlCpRBSnzfAqwe3LZAm6vU9Jk315c2wfFLw1biBc4bvIUatwP5IS8l3wTsBC28d
cfeDEGeURqZYXi1RVmFaCgBOxkWgM4g/rnASwzU1tWRTFY8r2ydoTbjR9gMoVB5QXFWt2wM5U/3+
IcnBIXBZZLNvNpqQeNSBTCQPuEuH/pN0vjGSGbJRmPPCxmRL3VblYImljRrvCCXCtYB8Xb12S9un
zJX/mcShroi4ThLfbeqcbzM75MPIcjwksTnTJ0u3MCgQcrJH0hCCfWRPI5Bo/COjDgyKWE6XvDwR
CVGP+/34pPQ4b/tpjMv7CQxQSvIWRX7Kgq6l9igGHvMoyW1qCmT/CudycUect4IK7BLmditPhbz4
9XZkUkP2C5bGemRFzzwxCWQ1ucuBO7433LiXJ35GL1v6orOV52dQBsMy5TgwML0ZyGuGX3/XxOOZ
2Z+hY2zCkyIblk5BykBZQhZ/nXTxXE55vNJFnN/W61tT2fK3CxDwVUdh0cnadqzHoC5xHJnjG4Vv
5FVR14z2LYItCOEVH9pX1lTtHRSuOlb423i3HzqK2NVP5rWR5OaP85VEyYFGLmLbA++jia/bdhau
DYHbtoSAu147RBsGPffwoYcES3fiGTAE3ttzOlmpIvpgVUfHc/46Ecy9+aKcJZ805sWHm4q5yh+s
e49ipzO+ekJNC7Jw8EStnlb9ywZWQ6hi8YFVwiebQDgn88hsrP5yHHKAtWSJC5S6PtFVfkOYnfi9
Pgfrw1uHpdHperPRdAkRAI7cc5ttd/2HV41eu2/jdbwFfcHsMJmbEKK33+CYzavtGtK7Amaf8j6Z
ptVB/Kw2EBozNBBX4x3TTllJ0OU+TiqfgxCYUbGda4EMRv2u0/8IoJ48/xOB3kda57z43m5daAFS
2VRETmnarr2/6aiByWRS00FeiOK4WfD4yCg8KmzEnlt+iR/c8NokfvEc6Yzbx9GrWtgVw6O5ro0N
6G1jVFWf4TLZnYW8snI5OOfszpTZ6p4GdOCSkctEjQGlF+e5jqSJJZLHL9SSIkEFZkNMnu8K9KmY
tDBu7a1COPoMFleoPNDiAjV902V5EoDG7C6WDDOwMHQ1uByFHLxB6Jd/D+YZrVDFRydcMDEDUKol
sT8lIjkVh/YTuv0JiTX56AfnyTtNQ4IuZ//SMdSYeXLNhdKFPhLQ9iQYTpA2z6wCtPOsEbIqa55z
BonMRF6ZnX3eYKxTuR45Jzgp4doiAcW8cd3mvZmk+BR9mCxK8STW1LUDL/4wJE23WRy2IfckCeqp
+MUovjAbmmBjt+ayZT56dCnDj9sVbgQ5NDznvuaMBxpnANBBLW8jY5HDM8t8Tjzr02mO3ScPmqZB
ISHZsQUD1xJ7WBJQSlerToVi3kgY2vK1Cm0JHNVinSNb4OFWVsNn3JXWVcnpMkBAobZtOTUJ6OVd
F+trqUOWQfFXw6k85JthIaRc1GQLutt29UxemFoZwXkkMWRdecPBqGL6UwxC8HTL9cIE5oXMKYjh
/tVhmLKzGYns7D4iL4BIzg0TukovVy6WWCMyFIMHoOry7K9VFfXXYfG+suD+Vtu5sYE1te7EAA5c
M03KtbWbE4tS9GqG4Xar/ZIaRHc5zDMs5iPEJdURiv83DfanMlyD6fN1Vdvd0bVmsNNhRALgyrLR
8q41k+A4QZPZ4m/Klw1bmkkts5iqaNp9XptdHp9Z8nMEKhOfy1zjBABdVUXS4nHTsSeDSUz0bpw/
QwPjEWPIdqbGpmkaR7jEpXzOsiQxAxL6uI8HXq9N1DN7fXXnSxKfzm2HKuhHOelAXCl/y/Lv3mTl
RQtzrLxBicXCoUvd9s8Tyy+y2DRl4pfrM4bs233vaiKrNoC5t9V/Y6NzkFd8rwalPLtyJD5FBzpu
xdNb8TRAGwALRev8U+OPk433rDqhFD7ZaoPeAGlaRyHy2nELlZPMQSndEl216A4TxgO6/axAaU6A
GQL0A6bKugyirG8deFfbSeziZN3gBGVXok5PNMKvtKc9tF2QUD+J7TiLFUUZbMvTCumfbvjB1lIY
PhynCWVrySS8MdKNv/Aa6m8swKyebct3wOwUFIhv34tPaHyxVnz202vZVsNaZtDO8JOo+tzGDF95
vNSNYqdRZmHzK15hm8hS0c07SHdxE2q1Tn7syXMZLudPp7v/wXzC3a7OSct7aAn1Je+9mUq3UNdi
HR/r/EZL/ueiv2q6pJJ+OYUbeKIyABbooQeFgBkMU3rCJesPgyGq8mftxuRJVaebvPDa0qSfE+xh
sC6gMN0BMHcgZRF87CFzyrIS0AArt0ljRPTRI9osOfXlWUjIWMyk7loTVlzwwWyWKHkCbB5Iijjf
0uBS6c/VHmML/dhnvN87dNPG3Ap7KhVZGDOTDhWnpHG/eUCfqbDPuqkqVb+DTjR8YRxitv4qF/yy
4HtUU5aufzUex2dPiuOCxHeXIg1p3/8yOGwPGgrgfp3J0vkjMp8hEhY5BOrMmI3SO4RmfHRyuXG7
WcWA4q/nr7rskE/nrny+F74GxxE3sj0CK0Ea2jZ7zXX+yzZGSTkTZTJlySWLFHF1Iq0qVxH7XZ/O
+SbrtYzjADy4m1gfGBsnbcc6ygs9S5fPtOccV+zg8WYumK26+Yoxve8B1rKI3j1UxSwSkzy0gVyr
K8wduAtcVapFRiASnt0BZjyDUngarZnzJxX5n9llDcyVncbq9p51H5oV79USyxygP5S3Hgh3vOJ5
43xYHl+eTX8i8thj6ranxJp9yMmxjgqweoqEJQYzmU5Kge7m7FVdHJ13BjEVt3AxDlnZIpvZyji7
mj45FgAFpJt7PYm2o/vFrDGsZ0hRcAnoPsr6Cn03QI8fgEVGxkuIEi86N21Dyv4ZSvIP45YahCJ/
2odkMoZbMQ6r5KCAknkNarfrAFyK0YylAmOFEW7RvSHfDEGBCPnbwwhRAgGidb2Vf16FsyzPLD1g
n+dfUqY1jjyXTyJ9QuvdVyszYtzK3gJwSRquFKxZCHA42aI77VhJrlfws1i2r9n5lx+IrJEsFrRV
OCAQca9ES/Ijusa9Ag1Je8EkwWUIJ2LGKGfXIs0ynSKboTFILKqwyYJUXNM0t/tz0B5NDucp/0H1
OB08xHIETKySyOfVjA3VK5E6RQBiRPffcbOIxSM7CC0aYOWAYzAhXcEoey9BZYk2o1CEhszdDNVz
0JDZ/8Neu8TYv1QAdbobC08ItCRpo7zKxSfKbzyMJIJTiwt8p7MBUyrzHqg+6rbKk/CCQwJwaBAW
tbgRP2uG8pEr3JksA9SabL/wup6ppO5zPYF2weiM4uaLvOyiE5gDtLsZV8zdUH0Lw8TJSdYofhff
lcX1CZRU6Fsp1P+RLPEpG/ShZcjzVLK8YqV+uB4xw4lQZnTIK5wr8TokHUYVRGnX3kmKcXg1Hj+u
7ppQD0VJeK77PcIsFRBo6rUm5Hoew16pKjo4U4mhvE8ksNIBbUpaHtvX+HmyCJIZtCwl3wA/YvpK
++5bWUA20FDoYloY+EF2ZLJghPplu8YCW9WG7f4mk5tUmFPNR/Sjc504dEoszBSjWjLtWqp9fpT1
jfXsORJnxXd44oHc/EScEuox88dsc9p0awAbIpyHehNML4KDUrVEq1lmxYmD/BJgb63kxw3fC8t7
0jxZqzO6CYcXDdqy9Hcw02AGMeAVw5hWjK0ovjNBqwl2uhgQjm86uBrMC/ekor8neyudowqekqO+
fkdlJ/Ae2qFVrqVqKmUUG96IDodb3k+L+Ef8VVuTaD3YrsHbOZ66a6s3Xun2nrFoFFWxk4FEWIAW
uviYUxBuzEQEQzW+i86ix5ghwGm6UF/OTQ28CBmb4ONfpk+ToZVFVF0DMZNttAb3UXJCdxnqiAnu
vL0GyAnmSEcLh/JQr2rJ0vLbNc6cjLUQf9Qu6zr5MFo+lFXz7K5c0797bFBPCSI1Q0gNz/tFe/Eg
iauNfEzohJoYbzc5cHPdVsQbpfv1mr8KGa/JfQHfvnK3thqQRZTqSkiEp2a6Q2aYtddor1c3ZKNm
7R38x2bqshsv4H02WzEmIxZ0yASR8nuOA7IIJthWA2VuSDKO/zJ3s6y23d3EijefaEsjwWJizcd4
uCIsZPhZ+dQCtIoAIuKduMXbhTRTb/OfeDabiskI5Neqq3s6RbXDZwWtVgYLtFplw+TX8OAKPU5r
SRyCHihkvifp9ohUqfr8lHTACvmJrhxnewNLgq2GWAyykeIUqTZJv833bu/CWSLiOpLTiCVkaZ7U
WatAtyTuCiuFsWBJa3/oD5hErp45xwBRd/97MSYUF+GjWsIFnEx50a+kbkk4311dnSJ0mkPj/hgr
903eXLgZr+0ydZT3YrhPRvTcfXCep0/AvsuJOcORIcmfDwqu4CIg90DfSkbpqpcWSv3WZ6w0CAU4
HROHhVwFUoW2lLOetOTRqFK/Y+00U0vTZG+3Fj7kU5qhAee21SsppAKONV25Q8MjzF03HYIi6dhp
sVDm2b8n8E4xcXIzKHzYNgrcA5/h5ASlYfAKEISYs5in6EWIacaW/EXg+a9mbYaszygiJW9YQd3u
PSJWD6Yex012Xvm3w/I3+p6MA2KmnKfHaEfmYSRmeiHqBjoQhCYQy+l+Ot9ql5bsvs479o7An4JJ
vcqtn5KqtXIQckmESUMSbcd4KJLJa56dAcHXUGsYn7quh+BEklW35IdjCKPm/NjJZb1WZcZGol8S
t7aPYUwgHGm8DknqqBExzJsYMcYu/Em3ri0Qw+ryBDKDDQZeBXNGAWgecPkFUXqVyFjDkxu+2wdu
nqc/4PVIP5kaiYQEqgoN5vzAf42vynMEWKpNdTRNfEmLK2D15oRT5YFHyg1LQlxH99O+tbpdFehs
yGvXcsdDKXUvSnyXDI/xV0Ko3nWVezi9KyyNDYmfcUAE/h6OSdtUYV0Ecq16F0dK4QfmIrcaQDCv
XqPzEfQv3jdIZfEWGkvsD8W4SYlGXvKX2y6ccGSlUKjhvfXpvO15eCk6jZeuOyvd+xjVyQtZt81F
suIRjsSHT6TsOYqPHkNy+Eq5/+HJUmzBiNPVk0ZNiWLf7pyTC+DcyxvOBmmA+DORgZ7A7EKKJQEq
xAMV0c3lAaDeIWgAwi8M57zm2MGEmSpF7DXbCf0b3CnuZASN64QiOXqSCWGe8wbQBpHV5Iotm2po
pT2aVxJ8YCKsg96TfrpqVowPGeXSfz5s5TOSVhn08NqlZOaDIR1XNp8hPt44I4z5wIffPkAA/cho
XJlYgy9yPjwonuZKVxDDeCsUTc26Z/yOE4BOuD+VLJmp/LqYqeQXE+hNwNYKZFdB4fp7y+67V5H2
OJvmkD2iEmARGVpoOyhLsbk+9frkCYZkg6VMeui7SOatsVRtqfX6U9nQmYNATKv5J5KBwrsQC9I1
0QW59GCDmtjTGhNLzbxbzZL1pJsZKHkrGkh9YGY2oe02GgCA8IhmkrnLr3M7tlcfI8iVx7hl8Ya0
VeFpERWgcohYC2LLMbm7G2n8aDzDAWj3NLJlUJCRw5CFO0T2eCGuMFLB0vnbBNdEoPNuyBv3KbGL
Vr0F/iSaUFyGs4nR65rWzxP+95bDOuOtnUsYUi6R7PdqJ8ZGlP5ILzHK8GodBxtZqLRiXCUp/iyx
IzlJeTj7CPTE5O8jNJMzkAXflGOyjTK1ToE6GpoKEWMpPWgvrIGeyR2PPzah8Z7LlfzmfjMTnzVC
0f4QhcFSxiONTLsURq0Z0sepriPMlEGNZfWC5ut06uY2GEcVAjrqJqBUG7m2SZBKuxarqOP5ttxH
6sijmin73lrNMowX/2C8ynvrXZezda5ZrT/ea2Teg5Mj82X25OT5R/ELm1JaX5SPzTo+GJuydO4A
AwLFyHmXeF77OuQAd+ycNxrFqkgeQbGJ7TSJGP61FSsLDJFtTRyhVyad3jFYK6RnVbNj7PLUkUn0
P3idVymnO1aO4xn785EEDZku7O4wD7MtyRMZbas3gCzW0pqOk2o0CTrJ+Cf+8JU18l0c5S3nDTOK
xJGUUW3Px3vqEg62tjWv31N71QRCMSHZmxKz4LHynafgkuM1+vj+S+HyjxYhrMPQJLTPBdN0lw0I
1Gi/ge++HJqMaFHGacu67bvNqW98F6x8rzGst+RvkyS7+zOJcbq23JdTpQDD0oK2a7zHT3y/yCkf
yGzzFRpRW/7ZxrV0pmloNU2QT/Wmh6z5+z2J/hfRr4cL7yWDcS+8BfX+EnSDQGK29FdoyOPnzkIA
KCI4jlLFSs5KQXtuQ1IOgVcBOQ++zWFPCqTAKt5oBpeloOj16ecFU/DYPxAPNN1tUA3siVi0ck+f
+Azc3DzBrQ+U3YqD1JA0C3bsxs93XPXbOXrdxrg2Z/wY+1TWzAV87MoQiqJ3Mgb3og7zGnknOKzg
eg0ZwsioYzRgmF2b671oVLBLe34iMonvaeV9Meecvlm2A2UElI+8qq8aRXAS4P+FxGcOUTPM2GGp
ezjZEbn1DCMvwAArDNemR5y9Z8J4F+Ql9l1iVppl96usINZNkCC2NswLjUApm/SeU7Zn0Ib5Wlio
4S5w6YdnegciooacivT7HIstoh5K2tVlW8uOZOS7GQ+UKo/tbr2f/9HL4s9Yp4q6CkFbWnoq8RNO
Dw1nmY2Su721sSRgn4BWOomeFg78aWF9/AIRKiG5+ky+FIPYFq/z2zDXc9N3Lpkny5NAKU0HEPpf
BYT2ZVMGIuq3P7fjV0Pjd8uk4wdNH/SocQbfNtNpFpzehGNFd86l7qxcf96/sVqyp3/etFbW/cqE
wUmOE1nXJDsg9yEltmjQ5YVvwAFaYLLb4cIl7npHavPEb1wQjUrS5Gw7/vMuKljQFwO6R4Uqmivp
8kMkLM0YJwa2gLVYxaDhu52FlAYekcj7dlGkj3+mR1CLf/AxOe/5fTwhNQf8ZCFK8hAaoOODhi0Y
Myb3qjX5D9Phqs8t+ohJ0iWQP+WFpHkjaKCYS69LRGUv2x3uPLbkzrXjIfy8r33l8JyYPdNdqd3J
JJRPFQIIhPXIycmzQ0Dfqo9BzNFI3VRoCN8PNDrDo8CUM273sBbvkZ5LXnIaiSOlq6ZpGNSqoWCS
P2bS8DBZKhMcfSHEGszFVbEQ8FkjMWymmX67JHRjDFRcQLiwhZ6CuMyv9kvUTJ/jcIz/Smqt5FBU
s8LuOyYnKt83VxukviQ2QRcQ9venHInC6R192w0bbOOHQ7jd91DHYVXrcO8H46sbXKKPffW7Eidd
/P78GbZ2A4LtJfMxlFaEfzVaKHzGYBEHrjUmRZYhQt1NgwoMMadoye7DH6pXbaBKOCSiuiXtu+3W
aPkCMh65qw/mJy4Du/15o2KY7MRYDs0GcPuGvdb1kt7uQqh2ldYdXpJed/HT9hFONSOsXm4MQXiZ
8c6y6psKAbKFKZWuD98qzhlYek3XXKQ1dFnccSZKfR6djBGXcB/a/dn5/rWuh2pHXONDvaRXtM0b
TbiAi8wU58rh3Q4+6hzmTzCZ3ijP1ZnUj2PPfbujG2o8nPOBGNKei1gAcgqnGzku20S5narizbPM
jZDY+cPjkuxAcIru85MRPVPzhW6Z0IESB7UOKf2r03CDw2QcHX74yiOoJdwNbg4QlFyjFwohVesd
Ek1p1dAYZwD65j8jznntPVxFrgYzB7Qww9YqSOMgD/LUr9yZy9HjFGfuPtHBPLZVaFw5RF63ee7k
EEAoaIC2mJtoUi5SppueHQCl9tkpL3F6Cn69jFhG+8JsTMogVLqDK8BNUdUg8sA32eCacY6hBh2j
euw8rn4Q0c64ObUE0mTMNHkMpRdlWneczGy+NwT/glG5GdchJHaEN6Ta+G3TbJ6w+iPUmUu1WzfM
tg3pYqK7umUYu8WyMW7GhliL7qwayFOIhwOybfBJf7xilO+yt6701vH/fb7apktem2o1NZPEKeEV
wHgtV8dsUDgWtIzeTx8ElizIB3fMn/NHm2aMZ+mVS3WOAPppB49np1MGkOMTKppL4uVxlAls3IeS
Akdsvtqabe/jkxDbCuVy6ujAerLlqphLw/7gCPlMiwLk7SHm68AzKie0HIQHrCaq8EGQMcgjzSiM
K5gH52lbAvKq/QjUZ7lo/XGHxN3Squ4xrvw2Qp1KmAfgZGD2t1v5bSkxma7eGqv7DcKiqSysFd1g
EReGpOkiJCC4oEd34AdMF2pK6JSLzF/b2XsSIGyW0mgpuS4/c16mBd8YYH/3bWnc+eQkLV5JAI3c
EnotqIoSx1NcQ9GJte0cOrtmesXlGRHL3Vsdy6QQYoxIk3bBRiccJ7Ww4vyDNPyFk4BrMXkj9qh5
cAo87/inMGrLLdPrjAar2LYZki//lS20w9agZ5tqi1Cc68aOLPGYYi8kTc1l17Z2cqkfDase77z7
e+Rxol2/IgxAfozdAyeqNKlHMOVW6ThqZrBevlQACEQ58s8h5cOPsz33pdI+qt3UEOySn+slroox
RmcbFw1DWlTKRn/z+JhyaLjC4xyqerfth11oxxCQYCrZkLBPHizLbOVIwGo/ZoEZs2ZvSHDPhIz6
i5RGEg0NF1qNqw+0FQn3RS8xyEIP91ycj1m+ONi2gHw13SugrBdDsXtRRmR8x3B113i8J2r8GTjO
GtDj8v+cCA0y9b8gKlmUabBbUoswNqaGoHsS85lDbAewJIhErmtltWk/ZiLGHa7zZk00VtEm2TQH
fKspAIu+OkzYF0Fr4HvTXhhMn7uMKTaIob6pgxUlpX6aCC+N8aG976dhbwGe2iFIlcznlyua0M1F
tgih6/smcjIkDx4wm2yJBjgg1NxAhiv3zVR7KScBRKZNN6zsrUBiNuL39SpVUtGrqlh4QYSwyL+/
abumQozgTC1mTY+am/Of2stWN5FHkWyN+vbnPwCqY3F0VOmixPUNr+o5LpKtnZjqm/Ue3zVu/2ei
r+l0UzLm2TI3e2GSlC9GEZ5abmTMrTFq3myeyMF+YnJtGWyKa8L6nR3ai+cxXtkN7QtbxuedcdmO
dii08aCXlFuw5AAPa7QxhsXQT3sT3geKNUCL71fRZ+H1BF3tENt4V/KyexBdb/qBOKIjZDoU5zMb
ycWmsgkBwik/oDDhaJ12DwpEKosk8iYvyhkWmpTI5mh7WWz4cItZ88ZQCKllk6Jhkgt6AiF+Nenb
CkvZNNJ5SqRuKbjVixGBeEBB7zc/7tbq/Rasi/6w5TH5QpmdV7dgzezfRMGD+ncywU4Q6HkgMCHp
40oNm585xKL1LJC4fyG7ctZnzl0APIHVGwasoTtns2fKFYbJuJ1h+22UvYgfejwmsLdhcxBexUn9
F6e037GlWdDV8FwrwcWx1uN4onP7O2gbHUvYh+z+qSUOJyDIaQJKn124rGlkU+qas2rs6/vroOaT
S+nTI71ryU2T2ijxMH7CGrU3sVg2peh1864hGBM4YqEUD2j7+tYsSLyM9d8woMEmC/Bg695nnmTs
EQbtFqorKCzscUjqM1LspHGDKCLupzHp7YS9nuhvV+5OEw26zCD0iI9aHsAnqep7pUDl5PC+utK0
lLlwwHfhG7zvSkbmNxar2E8DuENweiiP3IuX/7X7W2ZlJLePNqEEDLNDeJhUcXHAG5P1amVDnZFe
VCmiSNijvBHLBQE196bRCjeIzSOqTJBWlEcIP19KFth7CXtlK7YiddA4+ccGta9hphkMngzp2/YJ
ccDn5RFn7wni5ww4JeWmHz/299yMW2v/Ds4RLdoi3i+cxk2wHbABK9b1ra40Cl8i2irtVqHZJW9d
t4GPJuBzcI/e+R/8xKdaSsv3TnINRYn2mjRX1j580vmlITg2rEZFSGyxPtpRp1ZJyShvnOYj65TQ
0voVvJ51oFBGhVeuS+hwmHoQuJ2kWlbx1Ck/kzzhb9OUDZBRxrtFwlB8CgvfjXFnm1B7KRudwh+I
z6lNriYFHuvZlqB19/cXgNEAhAJz715NQAVXop4Zl54/ZwTyRbxa4Reiye8yccq2ByNvIEtNOUB7
ydVTcuJAOV+5aRIutIuX0MrzmRmp7j1vhWrjgGspwnRBZdUkgbntLha/xMVldj0+j9ArRBeQdghV
5h6dXiM1yan9fH5Dw247lpue8tB5638OakIQQ5Ym+lihN8YTduSVXWto/atgJKU7zdiSA1/BOxMa
Sj81FXX9zBjU1ihegAtoSkmpBqSje4gHwb3eD+LvqfxKjuvyPOdu5iPQsFT2ICKJjazX39EJdmvM
I0UD/ilQOD0ztC+gDMtMlr7UvqTBIJxuSOaX7lQ5oGRX9BExOdBp6s/Z7Y3Zz4eGyK114Faov0xk
/s0TNm505s5FRYhRdT9efvDO6ooStuSPkFQErc5nLPFn5ctLmCRmeXy9AHJ+e9ZjQW04INSki6Yv
q/UuclUE/ru9RIptXXSdDtTHJVeo6LXW9VDTCYoTvOV/zGbdT+0aKSWoN4sHgmwhLMqj8Gtvxmvn
ig+xnfnUBl+aSUq5+h3FdlOpvvHzvbchZjUVPehJFvnAgqWSYitgq1TJp7s/enhrqhjN+Mf/2u8V
0skEWEt09pkEqrjwexcEhX71nWCFmrH63te3ZlfRtOAkD3ZbQKjvFLqI74lIvzbLK/p//SLGf0J+
6AEv9uFWBcs/nESORr/lDJB4B1NAJkJwy3PGvSo0eHHyAOWagOW0go4nC1KwVDK0qbx79FVx1UMc
xF4PYilsAn7gzLz/7pTGKQBD99alGC5i1X3VHxJyfiue1uEclwPI1MRQPicJMXsJuFhaX01uK+hR
3Kz0wgjI7QJgiTqPL7EZ15kwTayieQGFmivA8eQw5kLvmO9bPIVZ4c3Q9upCAtOba2/GLc/giAZO
jRzrym+UI4cdavDnX5ZML4GPejXJdXNc73SVuKT0wCe0//7q6RHDI4oh83xKQdKMvGX96f8rSplK
1HYShZU5v/ren481zTC4ab7t3g/1ty22gjYjqeWSp2BqXBfJptxM25LHAd1nI2yKNv4RAvoJU48+
vKfUHDTmCl2+zbwWjLkd1VKKxV34HSeb8CFrQUiC9Aoext3POI3Xa/Zhf8ae4270eSA6wTKvia7l
sJQXXqUAP1Tpyo6x6ZFLm6BBGA1ylDxxfPw5fxGEnkUh7M2cyLQ/LMpBhBBwM+ShzXDe0eB1SGp5
5Qk5W/5mNMYT4ljwJtSermla3/WeGrDmbsr3GFp8j0POlFy9tvp9OZQygODC+joY4ufLXLQITgTS
Ha22h2AmIuf9Tj4knpr9ayo4OdTPe+l3x/6BdkjoueyHBbv+dbdguKshwOuU9z8LJZYTrEE6B/Fe
dAQuBcKdwG+A/P7yhLrHpUktrS+8MuYWKfuoSM4nil0A5mgvif6sZ7pgntx5NwgLyLg9Ubvwm/ZG
f0Ct0B5/s7K4ZKP8kKxUded5xlEY01ynhTZcrgWJCBIvZup0UP0fYD+dtVZgTtDLXOK4gwTyGl23
sqNcWKhatmQLWv5bj4AkiWosN9VPjcGX6cNZotoYsCf3TDhBGw3DcgbMfl2hLpuHCuPj2Vj9AMmO
b+edeujN9B+1+Y6VPiAXvhYtZA8hla/bEls4ecZ2DBq6iwoIAwmJBBdR3o9/TFLD8KekHQZHYKB+
Knn0wVs1cOmToLfBqGCJm/kGA9f4h0mgr2rLxWDZ8crr334IeacRRiB2D6LrfmStD+lTO02FglFt
k0BeXExGptuUAy1GkHTbnxN64O63CXwZn7IpAUabqLImQcLLGYZ+ASLuw3KY2TTJECuFzANvu4dx
Kz/J3cgVB5Rqzp6qzF0tTSjOZeorVKGBBadFxgBplIfuUyZ/vSaTUP7c4Van9qYQtc3ftPzXaC0p
7e+sxSRMe2K+tQJXuwy4hiUJ1bKXr9iewFYORCGPovXYzYYNTperZrinEalTsTO6moMdpQOvm6e5
AICkO4ckyW3LRT52IBeV5Nnr25i+KxnZWgXy8fzq6M5Su7aX7X6001dicl3XhrqT4kw56B5Y2dHo
Jw3WwXxFgx+pQ1DNaScdTMTj8reTS30ab3JJthkja9HPU/lmg3exEhHcRB9of6O3NO01s03w0pkv
hZFceGuGPrwNMFxHixa0hsN3GI6xl+osRVdApEmZjG/9Um7Uk84vihLxujL4pE0PvIbg0yjWyC3M
Hy5bJQ4HNXFT0ViLd23YBvenXMzuKu5UisVefN2yVta5R/R25zfHzBZAYk3q7zL9gFMiedqGQlw4
pTjxejAsmOMAOznXZCiX5HP4odX/CTfPZo5ILdcZtjrtaeYZLUeCiEauVtRTyyUzUVv8qi9v5GZK
YPHLr383vpQ9/0YU0TL+508KhFy5Ycg9z0PGoEGcR/XDcPWbeDn2mkkiVHHLzpvf+tNNtwZ6NuRx
eeqKO+zy+YT9qx+eULtowyX/kZn3BHFMRKKT/vkgDIHXYCxox9LShe6gvPEE1WD3MKuwqotJSlvZ
HkgxdFr73svboKINw34TI+AzOBM1YnpVJd91bf1gYdlZYMim8YFDCeqowX/pLVdomhNb1n5GjbVE
KpmcKUcQS+DHVPww2Pi2MrdSZb5KpBAj1qwb6P9KPWJ3fOHTXQwEkFm/+CdzW6LyOPdIa/57q5MJ
qTg71zUOgpt5K51ItFWGDWHfzq8MKReOvn8SrZtvO6xuX2eFz1p72a+IB9M3+1qxOjNeKUKrK20S
lCrb8KeQrQD6BAKiYcDhcl13mg+d9+eeFyl4KGaz28p/tPxQvRCUvPh2OLB1rrewupAqoVzvgNQY
tpYdGodZKa3EAPqurRq5/Cic2/jbATrpvutePXcIquBZBR1q2FQZ+NXaqHcM463uSnf9AEcbRNtn
T5Ftmaws3U9uWqrJ4lcIrzMUrDy/aCvaTpbADit+qQo/nk4s6jIga/3xBh764Ktu4HUZ5d/xV37/
xDdeewEPhq64GjtQX86VwTtMdXaaW1lqYS2BLdE7lma4Vrsf1Ax8um2Ubk365fVVxExwZETo1sWm
3oM7w3kGketjfh3Yah0w3GxrBEUada8udfxMFicfllWEEDNT0EbG84tgeXDEUxXRxrYbtad222NG
PsssGDQo/fr5FX5UeQ9C+hr0cENlTc77I+se1wPjlbGHNiZBukI3oyQrWWYa/OkqBqUtlYC7nSjG
otf9XqysjVe1JySQCwBepzEjsxSpPXc+Mn3yuqNO0ayi4g8grfb20XlwPleVh96/NMLPZsa0/Ez/
uZNkBIHhIyJjjsYX8xDdMCtQQtLCq0/U5VZz+xITOOFwD8kuwC4NgBgTog0Lv2O5BIUrSFLi52vj
ER8RbeAgSLkh6fpc9uBqZT7axZjz18b4QqO4Z6YNZj7usNd7/xkSuSVLZkhb4Upe7cZ8Z72CtKrq
7Gb6bBKB9jio5eR7Fr5XK/HhCptoZZtzy1YWN7qM/KN62mfyudtcofJwqzbvtmTGGphefPeqorrJ
sev329QBfPYQ6kGn/bz6wpKzn0eTCdieIr9amDaIh7hfTnuP9jUg8w4CADkmjWftjhvP3FRFyiCB
84Q+qFb1kbuyRQra2yJv/y5zR1vf3vuu4ZnFEDtXv2tsTclzxtmrOmJbYQGgI244jbDtjq0tpfoj
WwXw7X/T28bwWSe4j3QQikRME9lSCoVr5YAH57DxcuvPKrS8olE76WQ00gN6cjZdhRXPMWrFapkR
J4pHmTosScow7uUoeRU+Bhg/pNVbwcn88/RnJgdzDDutWJbEVcOn4SPRxd9QP+VJJyVMjmkP9jOj
vrZqLxQkCpqRN4AMVtx/KI0ugSgC358nQygOhJpB8k6njO6Pyt7ibr2G/Qs67DsOOwP0/qGFdXKA
SkY7p0RCOVO8gnL0JoxNKmuFQBePJmBMCHh1YYEyX5zPCUfjlT3C2sq3+aYxQEKW8ElubwMIPHAt
l2M22JGp6hAyMIwn0lr+icYEMLBfQY3MLmq2sP5SmUzF5zCQ3GGG73zrNQdCkG5ghepsTKy+BqJh
BlvGCsuch5M+sa2gC3U2LqU/ZdmrYl+RNWuD/D+EZdpenWW4fpFAhpjHGYWm6HvRdCnqG+gjwuGz
SdT839gefDb4uaub03zfVZY8IxD7hur2d5bFObrjdSJyYBjyYO5K5Z7Sla8Ge05CoeuJlmwVUcQt
bLRgmhPPMksguqZk92TJxaOjLDjaFVr5Xu2/POHNmRpoVewmQllEK2x9mKGWs+ACdjOhcCH70VV6
3ZdFjROcwXu7YArer6hr+9xWlyUyqAOmoYv/tNM1AXM7hgm3/qUGaYWQF3ykjcWiP03V8YUBJfqw
vuJx9GQuNQClVX8Z2H8tM6HH0jdWb8JgI0wmuC/YCCGuaYlqzf4xpMS5PHzFcZlXpbjsufC1Q3sa
PahU6hO7Ld4ODPWfNgzhvYr2Auf/gcXAOSE/1p47tGYrJQAaDkFzJxGtuUenCWfo56xAEt1MBzsQ
s2tfxGL9i6QULyaVN6uX3XZryIj7HwqvfjoA+PjjB2Zj0I4pLgYJFA11MFz/hdOow7eOVzFPpDpR
4jzK7fiQQSmSGj9eMsR1a2SRGR6twMeX6dFWFHXnyP4MTRh7bfdZhxiyXAl/YrkDAGUEnMZFSBCV
AP8Byi1VPQ9WKdJVwpmYw4VLN+fiQ/fcTBAdE1Aq783QpEkdghKMZIVNVj3qEqlyauti3kx403zk
zIOgQ+OFdOhF2oy/mvsPbv/fsXKHNS+YmFycPMiFKEevxa1zkAHsx8zrZ39xNqqwboPX7bcdJOSz
qyzUfxzMcZZkcg9QpxJwYijOX5CsF4RQOPr1TB5AlAEcmURzJti/IgJ6BUEWxDFRmDrxQASGO+Wi
XqhGMbXgaS0zyIYvhHU4LAa2ZPwi7c9WnxJWyDQ6yaafL0JrQtVvpzNz9Jboga+D+Y/h/QjqvAf7
Tl+MUh5+ICx58DD6dQgJ+s2A/NarEl527PI9lq5D7re8oZLA48bFrXdEhxA/Nk8azybbU5n18Nm9
zgt9LJe9OKvqbaThJNZf8csM9yBvh/HammJgatae7MetLFrSDU5TXkqAgA52dimAY9gWmKeK53nm
/R3w0gPLX8kF/kuj90X6IaIQrbKBBu8YJBdyxE5EVyQLUHN/ciUgW/DRJDOnqvks0PJIFDBXyVqs
eT3AaFMIIY2xAHSHo/ELzG2affzocYIywQgVMTvFBMLmflYVul8WWAXi3YwydRfFFfD9n3Ext5XX
T0av9Ffxbbwnvb7Z7s8VbHXAnRxjxiEqL09j2zDDPhhkkCS/nBbn3pKJJbSulvCg3oQWF3BLm2gc
0ZyMxxGW2WvpAbXrjS5gvlXCPml2aI04+XbGaAhUyVlKHPVfUa0jdkvQiQH1lM8uhOl/R8Fck0Qw
9vZXt74obuXJxb0+DMYxDUohn8aGQe8WGnQ/BwIjmPPu6cehWakovyJAPj9zY8xelxzoAHKrzxFq
eXjPhyNDOdReA+17CgNPHI89vJ+BzPjN4UKAPR4NwuQSHzWpRamlZTbLEDyLGW4kDdaLiO0luoQ6
TbukcApEzTx+J98Vrw8bZXW9eEXMXGoq/B73JlILYxaLdG7DzQM0yGABrbr6cHruf1H/RTr2H0jC
SHjfVEVdfVU8NMF+lO+Fvpnc9BKS7QUJgGuR6m8Qp63OmxrHafx+Bp7de6RKZhUeWsbJuUuLqDEf
tn747PluNxeWxPyK2rQED6IL0Odfnmn8+TW3ta7BidNdDC8q1w+5hEPlDLR0eyhAGfznvsodFygB
NqRhMVqDqEG02jJUjDTaiEoRuJUjQ0Kebbr7YPbhjjoLHgmPuOPWR63M6fFZ/YrQF+IDlwA+Urec
Fq76+6zxKxB5MzMbTM6hRCfs/4M3n8DcuyhTioV8l9TqixFGoOtpIjJNelkt3Ig5NbJ7vAOdlSHi
KJOQXM7+YBcTDNIIZKsVvwxlHA4+iqktkufesNIPM/vv3/tRL4TFwUWkcxHoqLSU3aDSucOGrKvn
3uGvJIrKQhVfVcHIJZMxqQ8P/Mnc4Rv5fMONc/4n8Xo1Klb0WEZy9n9p3iQW46L5KXyzSeZtbh+p
4w1ub5F92XTz5AM4wtmgtLLqEJP24WiIXkTJaS8O2qUYvEC1wA5QZ0/CKdjSqUYQEi62ejJFcXtn
rp523S31//HIyZSTN9H6iNupmkfyD4VSbtQ/6ykxG8fshRE8b7MUqUGHgAcF/sQBNoiUzLZOEFg3
xFFTl8Sr3imj3I4srExGbHCLew/4HAZar5bTQO6DPY16O3mqqgIx67uZQB3jTn8XM7F/8tbL8ThY
x6sjwkyzuCCJx3t5LqZQToOsHdYzHlkoX6pA/wzG39+XAQTERhMgAX+zGUH4sRNwWiNuT7cCllKk
BbYJSeYxd6WIsnayWPaJnQYYpcQ3inMlBejCgR2EldjsXtpTUMNLLmeS710nNVp1/EPUFlaO3LS/
ApdDlu3H/pn7Fr/7pLZoXarZmasak6rR6r16VleH0YUIJJ9QRSJMX0/n3jkCvmmpHlXAoaHnHdTK
ZyClfHC6idm/epIFYrERMNH+TaMgAfjObylMJwsvrbkfgBAe2CKk/h4BFJiGtSo+hrQLEVFPnvS7
dpPw6zZrk8BalVPN/uL4nctr/kJtDNOtxAlu3M3lyIb5smud2LatTlHEYH7FoOb0cRy2BiqP1M12
LAGXSsaVV5Vk98b9/tqak8UMMmXoLqM4LKcJdb/BCdZDdbAUrXT3cXRK5exQta4LddySdQNHTWXN
ObEBNRX97lNTTyPq1Vix88hCpTYWd7OKHr1wCuFzhVDF3miCTDHTAxIa0LPKrudYZEUpcnNe22qR
5UKsLON6UFNLz7HQwEqymuYU0L8c/vkQz+Ll1k2VbnejXPtZVr2ipvbS7fcxgazYKaa1PoNb8l2j
bRKFkskpztojWGwT3X6KJibW56i1536sE0lP3svmLBPahj82J53QVqaDhDAd+JJB5agE5rc2G6pS
BFh/qtMvkyk8JzvSTv0XM73y5RJeKgylv1QjHjwl80G5wl1cgBaDa8fMccJemy7omH7qmJMeIP28
YynigHFyhjwPvPm4lqi31lEuWWYMYu9MNBTQ/ZAf6s0GPQPtpFTv7He0hzdJ+W3xya+7j18tmqNb
KzM53l/XmczRREjQBL3Xl4X0Ol2N9pbRn5O/a7PyhMGb/xDgl3rEx7Pde02fOC3Wt5pRFtXliGv8
2XzioWHtY2ruKkSSsu9HWV3tpq/TsuwkxocVOOXCHtUgB3pPe45uX6R+VKeN5DUcvJfmXjIc5+oq
cN4TxRcuMWL7qC8JKYraFxpljaEcGDBWoKbrNneYNXQo2SYMTieuRQrtHi99h/zqBWXl5IzP3tp5
vIAjhnrL5/o9NRi2GZsPUf/BmBD90g7JigNPLlRn0AWVEchowj/lR7repm9R//Jfu5QbNo26z2IZ
WyJ4mjctf+X+9kOMbTa71T1DgVJi6k4OncJAApWXmOrbIE/iLMp3zJ7q7MiCuSvGYkhOCVpZW8PS
8CL+D26UV6CEW8JqrcgNHms6AN0LWDpktZpbwnFN+Wvx66mT3xjBQbKtemVQQB83KcQ7Z4DJV5hn
MEYLHwpe4U9L24+uubuIqoK6bAEH32F1Ic2C1B5ttj+i+5YlotFN5rWjsSkUd1OxyAywIlkJRg61
2GumyLR3fCsitgsPt4kOhJhX0w7lW49Vg1E0NcIoLybWztmp6ue2WBnia0kBxsbXhw59EBq6HK7H
S1Yj3d9k056lNBuBmlJ/VMGQn3MZDFkvelBZl6mGhdmdBY21m3DJ36V8r/oniEkR2oQio5O8Y1vv
wdL2A/sJjthnjN0LzX4xMppUyzwH7j9cJKCqHKZSd4hhlMOKwyQjKnc8+ASwJrib7Jq1GZmkKvKD
qUrpcfC85/4JcJp9veu2CfmAJMyS6ZU8oqWbh55LRJeNrYGsnwiUGtuTdewPbJcS3ACh0rdGt7uE
L1+W60TsY2B7dALD9B6/x8pRYMECxAY2yH/TPaaipnkvZFDEsF2pCTlkeS7Ejqq/mk2DfHM1EjBi
KY8o8eMeU76HjX3Xz4o60lS1Fru9GIuetL4bvw237MQkTciYxRcyTGG3djCi638ovu3YRMzv61d8
TTpwsZnJ+VA6i5gUh4y3lr/2sLWwqeVhQRiLpA7H0ufrVZHIfW4uQAtI7LddJZGRDzToLwKTXJ8j
Z3bVfFzqc1GXmGJjDB2z8OAK8SaHdd4JnoYFDHjdssNoqYErR03CbjQZu17qAVP8kKj6dH8kluag
f5oHRhGSVaLj+kWy4WPoRQ2ZrIEVhVuF1Ol96AKVe+0R64uiSEnoYAF7frneuOuq+unAOkXybnV1
qz1zueM/VUAHbt7stC/7iHGxCXR5h75O28N0jYxmefNl58fH/v4j3E3ZTZNIlnLaEXSJypbaHDjv
++sx7eXwIkaYVLmg23/SfWEH0Nm2cD2Zlkfd5iiGuY8sVKkTYXAENMtVuRPk8XhZsd6Iqg/ghvBH
292btppWAUSb5W3L9HVPdWHlNLl2VE+envlUhhbkZuxxGnvpY8v2x3Bl9b3TZ7Nfuhjph5IxoYBz
lpJeZpNZnxOXWKT+dONHWA8islIuBlr4hu6Q7klaGDVSUg2HDfrgodfaW12EAoS0Rl0BRDNzqtbr
eqY0rAZw9/gutkrE70lebWtBMdUygv2N4/I99o0EK/YbovHaRhl/RrPIGjq5Ri0IfvPRXn/WMIuP
aze9rxkD0AbamBqIB9/WTnxHo8ME3kyO0216KT+WfmeONK3D8oM1wvKnzw5cZIy+pLcrQU02O06+
czEf+GYMH6PQN25kbvAC9ZBLnd/ZOvSsk6n07Uy7Unp88V2GvCIp4JhV1S6bm2ahK8l59ZYrw5Gw
4E9iu9aKavO0xq38Ye71uBG4vvQPqEJZXGHZ1S8wQOU1XasdpWJmpiqSPGlytnIbhVMyd/LGPbZL
Gi78kS84oPJCiq+gr5u8bI7b1icBFsZqYjebZ5xMNxOaxhxXarVSbbYpAchdY92cD86giZHlsqQG
TYFKUtsCbQpqehMhoZBpVsYRFOwlu0yMaWAAWncczGhyqgYeCFpnJHq2sByYTqn1AUmmj/VE+tQ+
j5yc1dNKMqvo+F4T4SMgw0v7X+eZnuY1/UTsrKU9RopGrYhqey4lMw3BJpZecSdujaYkRymV2ZZp
5WbTrciRiApVtBNXP7SxQRdcMgJDzX5owb2m5lFXU4TiIGmnCT15lYPt3i/YavUDPtWGRJkuAzTG
/gTRGvEjEC6KrLZG+2nl4acG8u6nXfC0MsbQBBGePRsjGf6pjGa17W1wuW56ZT6sthGBPHdK9cyf
+WZA8KNqYV4xubCsJ1WlrNoe1gf3PcVjBNogl45Uhtk6R+lOZmWV0058zay6oZLVtb5FVLQUXwz8
R26L/I3FYprODQ7jQuNm5NwT5nio6sJ4UbiFW3IC6YeKeoWG+lfNs/4WmvxaHzQ+Um4p6pRfvK1s
aIyknLXZ9Gh5c5KVtUlG1OsrktTjyn1WVHxqcv2OTXnW7Pv61AH8NtdLFYchsrra/oiUrvrs1v7/
cCuzsvtHjsL7a9se9PVHVDLKN3IBQ7tG2Q4wPTapk2TqJOG3I5uvloFdw069QofpjY+hqLGZVziH
4OLlsrr5Zds0fTcb1VJrVqgCJI0QUBB4qJIumR9IWB96Q8T46RllHuqJbK5VZt/BAD0YFgtrC7eI
cUAZTtcKAIxI1FihqHUuA873mvz/uRW5A38eGJLDUSibVnzsfQjwCdMLz137KPclfajZMoGX0+Mz
75sl0Qp2hwBQIxJOmEP0fc1JQk4paZpc02y87PPwP1obu7YxTNf6gUU0hiB+ad35bEyUgbWHhIuQ
y7AtKSKtE4sA4AOjWNlvly0OhF+2oPDBG39tnskdXot3vyn5iZbpkukBLb5gi+U7dff4Rg0u7FBT
L7xzi3B0MLGdZfugJ+ZEgGRcd2D/w2IoLCuoin8DpOIDRvJbD7sZIYcRgyFC0lMeEwiAlBiEYUyL
p8t68HBI6IKi77zZTWZbI40saEtNSznTgVoZHHiD8tKzo2E20rZzwrmLX4R7jPtfdWnjGlkpmjU1
tyGTBXVvmo/TQAtUBRB9FF6DQmLdm1kkS6PppFFqPhHLjBVhNhOnE92iMVpjp/IrqKZ0wyGVYQNp
Xinv0DmmAyH0DxFNYIw2V3FWaw6nMZhbjHHcqqn7eGuTQMqljbBNDmIko38frAWgWMfuUzE9PEIr
cqRE7TeTrK4g76tci+GqP16kXIv7uBQnDqAjRlzHuwShiLWns6bEYYnCvhjgNwxtnXFj3hjf0tqQ
vWId5Sj9Wyse9eeX1hT5iYUmlo5IXiX3O/a1s3NMggZvB5VdqVHdiPgYVcUXuVXzhx6ksssmpcx/
BL/K3PVG8uR5zS3C0CEFG/50nVWGpDZO4JDgYum4C2eMlEs/8dGpodPhGDAXwscUPb70vg5cmdHg
hIpegUnPOVEZzEReVZQ9Nz6I8B7Ro2sY4qUOqwH8cLj+63GmM/1AjxuJQvkU3lefGc2SSJTaPujL
202ArXYQ3JPf2GM0E9ZVHItYVqEQiuSA+n7leDVaYHbE5KZ23S5oRSFi9h7mBlj6vhnE59cvMaky
+ycrUdPkoYAFJP5/2bLvHvsf8ZNEgM+zNxxM0TuKw6H1MwBFLqfB0mEyK5hibMzybLgJoXqksh+L
ql6ivMbOg9WfoP2oGkbWTfNXrbRgpMHL1YdfLWvyhaJ00pKEKkRJqxuO24oTm8oaLxXpzRUtE2F0
MmN1Ni0OqNWcLx5Dy9EpgcwAc3WYPyzBTI0pXVurbtkJLfH06md+ojnIcP0hZ6BzMeq0fzniDBdh
cH8wJwFhtImMBpr/S7iAGTKtFKkV/1jJvCg6MkFjBnxqGRt48ZNHBnzjLMW6leowVp0t/BOGCAP7
WMKlHz4ojfdFIfLr7yisyIZQW398qylmq6B35hLQmv4DEovxP36aSMCQ7WowUegEWcpQgHZOg+Zh
8umgTaUQbo7ETuQf/CjS7bMIN6mrHAPPpLyfuHlrdO4uzUXUri6NpQt3AqFpFLXIg1d44eFDfMql
P5hmh9OnEdaEkRbKqdRtV55pSwRN3ntuRMyJxHXIC4oaVOrs3Vz/f5+qhzVGQvX5GbM0ly9suwMI
pPKvnI+ZfPXN8GBRY9ZjzDmf9eQ2E9Xm/NwtrIMoRWr0iNw8M5ZNxI7VlBawLscoyHXc+7NLpPH7
s3EWG00OOkNwhrciE4qhhVZ/0ryyDTnbsyigIVydfpDNRAgnBExD8SXIUqQTxtiMpnLviaNHu89A
D57smTu/eJf5agZ4slb6gBe4PVO5NdllCpKBQRweLUIbH4WIA0dKldLwVp8LybmHi6YzkKjnqKP6
3RAphC6/FgHzDJFrBY3ZOzyDheKv937oLJaSp3cqw6v1xC20ai+gYUdku4hXXfoKTK4GQGKAV8Uf
n6gczFv0QHkhQCTB6zev68NzLkUMYoc+IsuAhXHTxFujT1kb75hbvDLYIe7alcEJUUA1vy/ECd/j
vt6eE4bQ68g2Ph0BHw65c8Z6PQTzP9fLWmWkg/dmi5BmhaPi1kz4gO9WKMDAhkZ+SsDhLffaxlJO
pegzIPzJXuiutTHo0iZ+8ZZd+9rkGar17Ok5iJyq0UDDm0l5wuzH0AmTCk1uUJrGTcBHWWV3JMNb
mg6hZ3HHLKleWkrbn6IeGNYoF8jbePeeXDVJMv142kEuPAtukbDg8d9xk/5Tth/Wr6KEdNpFXReS
29lj12ZV0ckRniYV0ioeNK6a+pQSzRR3vpUHq+TQMzfwssVYJGETMSdXey3RPHaGggKEedzW9jTs
UjbcHsdrlqpG1EJUYuST4pyFkai84drERMpH8cPqJ20UaFplro7FIw3GP5LTrQKRP77idiud16og
vKredR1sKgmSKtmYoTsHa3iu1aYUONqFBq2lRlKg6U/sAa4EIWvUsEWS/8kHTU6TkeRH/zTGRb1r
o2TSecPTMClkgThi2PfBs0IqBRDUmvQ/Z0yTYWU4t+jR698grclnwZTKHWbfb8fwvfjoOWNZ8QWv
Np1qFbsBT3iN6sAMw4CJyP0yURHEnYZAsJO3BGxE6+7AfOJmJb8o6GgbROTLxkoLLA3qHlQCzx8E
MxFTNhgfovvNya9maEO6H/Sl3KD0ygxLplK0ww5iTs6De4tDbH3kzM4gLotPTcmWfTwJHJ/x+fPR
mgndKde7H/8lKvW7KVpTdltN+LL8GZo+l5XXNUhIYGp3P4pOkRd/JPHgKZbWn4nds9BcvJ0wpgiS
tRjNoPcdJZ/ijGNufX5ctCLKw9BTpwI4oNjHDw8nERms0SI+f1fh0NbXhg7FpOWeYS9DGRCktha1
yR4dNsJgdGvPMOgY36Ut+ENEeQ25buORyUAMorTn68dt33WxEejP8YhwmsnfPnhqOP0qfDdYGKr0
z9wMKf4oHrvDzAUXCkKRh5nK7+ajpvEwgIz6x0HW0qqdxzNO5WSZR3qi+XzkK8iqVVWp3qFSvUzV
xyATAdjLTBCH7B87KV7RipW1d9XOpkCjR6Mmf1j/5q3GCrnAfrDQmFMeoowOlsNvQxOpfy9QF5rc
at7B+vxV8ahpp4f2z1DCYg6UApGRPKHExIG767LbxVX7qNYk2RWGkxEClyt6uj/2G8BSWU6CNzah
/Rx7lZPYr1gqlCSCZ78O2eTRIYUlIweyM+yNGxY1jLYOGpBcdRkllwa0bE+crB/peuvFQX/UrHYS
w8VA1nPNHakgtP7AG/eGU3XZc3wb7ow4WPrvTHlIv4K9WwVw/IRDi0ks5+splJ/Rj41nAkmGfUCU
uonQk3qs/XilVHdrJHuW6JS8QjjqIc3msmxorRQWiq116by2TK4LUnkCNF966lF+mDPJR+EMn1r+
aStJ//D8fRJkuWmOi2MuvRPg8/1dtuYq4wMdpH6EyYfbvpoovIg6obu9NtXYTO/j6b80XcMT6fOd
kxH+flUdkrzdnY1spZc+CvbR19Th1wG0GiVc31NiiIirQmCDYpL6GnjmyEW6EkfyWB2VnYL7BuIr
bsNKnOJN6gNPzNaW+8nUJFJAozLtJo7/5cXB0/o353V9KftnovX47Tw4fjgzzY2/6HEHs5wkN7vp
dkh/BM6O6QET4+z9PGQbjWKLM22mJulrHY4iDFz9LKZ9Lkjy5SWE6KQXPz9+dcqS7B6FLjkGDXEA
nJBnb0g9cpoUAo6p4odylymprEJt0I3u8a86utRO4GJld8K0fm0o+g35S5GS6sYRkT1MA0MIw1zp
YhjQ6FGwLQUXWuPPf3bLgvcpIwqy0NcEkqwW9SbRGVkcm7QrfEKeKswLPobkhhwopqMgWhDpe4+h
/hyQU0SyMMqI82lLm7qBYwbhY/Ljzh9P7ZKbHGR/uUagDqvXSISMqKVsNIeAYe5XSl0VP3ojISuk
ZSChvpdLnLgcKKeoxNtD7GsR6jTgxvYMOuGw2OsBsKJfaaXTOZua4Q7L/U730WeFUW8mgutleJCb
1a9yqwC0qa6YsITq7EyzqQ3cuoW/1TPOrykxLiScty0TOgCygycNbXjb87rtzTmwCIr5lknx0v3L
mNzwBZ9HpPKPvXMm0U5KQrK11SIGvCydg/G16KPg07INTyWUN4SZ+i6I/yZNsIE5qGzrJwF9K6uQ
ZukCX4WANU0uOaHrZrb4f+q9QfKF1SiVo67h2249yQDOWzl2SgbJj7CMPND22tNtdkxbT5e5Pbls
2n7LtAGD0wMrLdoioOWh3VMaJigvdgXRv3jd1vgUlAO1OTdUWmCsdJJ1KklxYLb22SgnEy12invw
j5sPDKjnLphaLdx6huvm1k5gS36glAIMuEYZzqiwTuQji13ms8QJz25Xr8XoPFbsIJnmbLLMfmt0
+Oi+uA4K+OJpnzFOlbarVOMOGEPcsLO3tBGL6GbhVxHjgu9V+QnY8KorHU0wwaAwClUC+LQMTnlY
Wf4sbftZwiRmoQ4tSmhY4pQOydjJhz9rclan56JbPMDYe7aGzfcnSIvv7T9Jxq/HQU9gCq7FFiQy
hso00KxUCTaQ+EwUiV2gbmrt1e/kC84GM3J8vFAi3dxYZjhK0FubF9i0R8pm4xX1TMTgyyBxE2TU
2aHAABo+cIk0JOMLqiXNxwBZdC0Ff8K7yJkSCPii+WG30ZMbL3PQYtwlv8SozfW3qrfkQRI+t8NS
/k8P7uM0v0lmRq0N6K8XeeC20l3Ail+aDx98a8pHgGOL7WNmolSHT8TfoqS5RTUdk5VeNyY8ML+U
8zUiXxIoynOYj0L7RVLuYYopPeUbc7j4/jXU8gSgxh9XOmimLPYSKphvkR2J30IIM4fhlsNJ+MZo
dcWNFWBWKF+XVUtxgpE9tqf4QHBE+kVHrCybCkep+6Zs8oW25xoRDTwFnwqb+GuvbHQdUOVmhA8n
GXhoWESch9feRoZ7HiHwdKQIMqXX8VuWgAhieMDsUYHYzlA2jecrrZcLunJ/4GBNrlaqVTLEaI+9
hTGLxDkzXImgtzf181Xhsjc9Rtpv/bvxqbxspCpdAaTn9id6kX0WAa10/jPku9y7lYITJwfg/5TO
kkhGk7LpoQ6kDkMEAflQzDHhqTa100SERVxfcX9DfdBzmYppTegryaiWBl1eXWNRsQ1NViVdYqtf
uSo41UjnmNNqs0HY5p0XhhmijAzRvzwV7ZxwfTOqeFDNMx+Rt/sx8ePGbvdhoEKSJuA/s/JFwXHy
rjYyRrg+ThzkonLuZTRCkQFsXv7AUQSk7VHVnzSRogllogRAi7NGz2HoOSyDj6iR20THMKprhf7S
2ucJqh5hOneJ7Uz/KE99MyJ+OwTkmuedSL2S+Vb5BE+pCMDBwubtJ54Wv8wWTIvr0SfrfwUnad9o
Le5gl8WZQUkHjn0n/5hMu294sYhEal73B+qcGQCIjyvkmypUWH2iA5c9fiBAIXeiAUiYhkIV+n1R
+7GZ5R5L/VkvLNYkNk+5B0G9xAArVMSi6GcxEX9RcbW43tHapmw05bBZ+iHbDeZM+Yj8RhJuY+FY
yJJtAz6ndHwoqhRHp6CYCQE9VaQkpF5x2mgi34psqzmyfL4MVthxJUU4wpEbaTik9Mc9DdTNC5e3
vkVtZXthYekwUhJ2IhZ+J3ZHkR1GB1qHpUHp5fU6udyEYet8UxsCbMuuUsX76+I+5H7WnnAWRZkT
oXWqBRZFGcKpS9Magh/iImQn+RtsNzj5lfewHpJkJbSrNOQ1VURHngBpn1hM9o0mI2WMT1KcIy+y
AV3Xelq2hfwMMWFrfgjjDRWtUwEod0PhLomVMICihicighY+YqKz/8ER8g6mqoYwzjaCOlep57z3
PnweeZTVliNBgzLjneCi+HEMYvAb5QeBtjRXSZYStf2fc/kqbEjT/2thVr3p7wxnDh8RmaFzF/CZ
s/yPbu6/XM9UUhD36WSE9z6//XaMXTDuWu9/TKxhxP+8kMVuYhAHCygXkdanUIwzcS/dnAsP8DlP
wrf8f83oI9CWG7lhtUKbAIanXDBSzCHMMFgsy5rqjhnLhvu2OjoJi1HQW/bI1CXmNsoZ3aOS82D8
K5hXLwqgpGXOnsl//5iOlBhHh3q58pqwfrTuyKkKVNTzsb/tw/20YmOFe01Zk0sOOG77Di53jaY7
BVJFl1sNOGc5UYRGRhuVJkh/bfH55GSYheEHyPHlxvg9BTby6W8qlOWDr0iadUvs106EQmb/Ij1t
30+3C97+paLxQnm3iQScQussOUBzUk1pyVqstjm/AfgcbEFuKH7cGo77nG3K9R94gN/UatfVUunX
5fuSAE6Fv9icnI9kJfKNUYTpy0tsaEiMu9pYrBRVzutQ0lhazIBZBrgVveNbl8rreLqe7ERbUmve
Y0CGYmNhxoKu2yHHaPWEOEqOvyQ/teQl4cAV8I1K5+IMBus7nu+gj+O5s5c79dkjQjKOolaTRRpO
gbmmKlVChIvQXEt4R310ENWDg032bomzm2NBfaqHkr0D3Kz7fGXegdrtnmFBi8/YtPwiP1Jg8WTR
JwETCLekfLSquOGK8RPloKHBwygqBQbVRjEs+VWCV6jIyIaAh4FBYfu9v24jRu+mGf2xxpCSo+xl
lnQBf7Rkdmq/wdKu4X5M0t0CtNosLcWeHrVOOSatB+nvqEHqobO+zEj0YvWB/CQJuVLPCUVQw/wN
Axa4orvAIgJ9L6k9z11DwfByWx2jmAsT/PBkjOjbgNT813ECXPDU1C7NCQEZWuqRk622FOePXlKW
gvJARURv6dKksQx3S/f8QjlOAdmrJ+6of1kcUmLtfea5SDdMbNXjBOVCH/yTzEDl1ftYt6BFMbvd
BALzvO/fWuxUPYVAwY40+5x73OxfX4ckpY+E8Y55yVhGUJUaO4mqek7dJjn30gY8vCfbuv85qmEQ
LoZuZRrOjg+KgPEA4M/TMiJADDVIsvHpXV6W1sSxr6mAFAR+cN8XTeYe9Ob0fH7SRZhCdNOR60wO
0nbwAK8t7GLBtI05NbagLWez4NyVtjewHJ4KIl8ov/gTnMlOKB+BI/AfLHfR8v1Q4fFheRRMQOw4
yNgfLkC9VbE5gR8mjoNLUXhtcDFAIaSnrOr0YCagUr06sLc8GndM99aM8z/p2Mk+FoRKRU5cQNlt
65unt8ITyMFJEeNlYKFhhmFqPj8mRi6zW6TCx5NG2h+Rvz1WFRLrGqYxCLmZzOiBWngq4PDlGJuz
KCmtNNQIoQp0pWAhDSwGdbxWjrMrnLWhrAfUYEY4D+kM3Y4sSY0Sr/DVGOTvVpwPDxPz1fQCyN9u
02wCv0G30Vf1ABiEk60n65EvLzcHiqyCMMtVxCkxsDDGhiwXFUm1J/SPhQ2vH3esRy/ffbtvErxc
FtFvgH0bd/xd16/IZpugh3G7ADsdwjNrIZU/CHhIR9WD4mPgcEf0s0naMSh0qAZMJZuOkCOtQjT7
f9vhgsy2RemVqsOdR/Z32asWAUM3YDZIdlXOKmLdcd7t47yRqiZb4PH3jfSY7oWyhP4UBWgJSCIg
4296ieshoNb1PfGbY2V8o4H3xUv7FXLaV/ZCR0BZqcVyasZ0D5Iaiq68T9xdTQwFtrjdUvmn3xej
eUX/OeVLDVw7PLEFan81GRI/XzCIjQ/p4e3Mzcmi+9KnySI2dklVIvzlfANIIKrq3Fg+EQAPq5Lv
uCTLeSvpJEam7/0S5b/kwzlOHmQbWesUsje6bG5sfo6BC8RgZUPlKfqL42vTXlkSo8NUAqMw7Esq
4rUFZwVdSsry4J3d/aAS/lb0FOs7u+lwD+qzWnSY81t5ZQrPHriXAZJr6AyxvhuYgkf4eQZ0rqRv
rBmSYGhhKX1QmqmhnGsCnF9NMjOYOqphJZQaDkXkmlM1SDEwOPAW59EVpFe0tPsGOeUQPq1NW7tf
YkGRJwcfvTJqYJIMcIVVZns8TBuAwxWJQ2nvLeSXrvvf4ps3nKEy9Li/g01IIcK2MP9DB5M8b3fL
GPRZ3YmtXet3AUGKG6Ypbu0pXDFnkDFXV9gWb4Um85/Ed3N/4b0qmGI5w2KjfaFza2wtsBlO/RPQ
QohAb+YV6abipTF6PnpdkEIUQS3I4xj/o34MFNkSLb4m1Datav5tfd5oUa5gT51Gm0ZUW/afumPF
p9NFB2BDbRmxMn4re7uLrTTVmV6r94ZHobJSoROVooG2SeWn83Xf/UhfecG5Ye+65OD7kok7kCxA
JnPq7BYjKwXijV4d9s8hJppVObUOWuQdJdsZZtLD6yjlhFzgkXWDWvkyFwA5Bp5LCr+cYwETlfmQ
s9rJmKBI+N6+MZjyg/T7c/yTFRPiAU6IrWe5k+6I+9qq4h2bwuYCWHfikBOacllnci31tIU7RJ4E
2sbMdJ5upoxjQl3QVvuE6FmETi+9eCSZr2GIMnXAatQ3N3XwgqYjj3yu88WzpXAFjin9HsPIlE67
I2qB6Omb6fhjOyQYlww3L6J+DGzJwNnAOj2LCfz1/S5OOQxulf2TGXyoN8v8FIvPzL6cXiYxwhg/
u12pY9/rhs3vQRQvS87s+ML1ZUB5UJG5Embz5rsv8Bl0taXQdlspVntihcCBAZj1XZsH5zaraQ1t
xmLTjOTp865+IYMwA5IKjFFE4I9bS4JDWrRpiR7NKi36URIb7Ro6Ghyxu/Tt0GY0aaONndj898Xz
lAN61toOTsH4l4C4yHSK1COJgPWb/LdtC4OX719SmqID7YylZYWG3kiz7kIknOfLjkHWDRNoeaNk
MIsmmWdfYI+z5S4vL18KZ1B/d2XXJ7YLLCqbLWlv1lq/lsEm79xyTj1uK9qBe73ql8nwhDZBcpv4
LthRH0mJSIaoOHPTNDxH8GzN+9nbNfx2iSn0Y8blP/yUKCgsYOR3rdG0YZ/wxY78uxjsqTGhFNTP
AYnFZlRR/grZglMcE3w54/64NdtOVuCz34UnVZzGyZLZnveau1eOMYdLUxBFfh1a+Bgnj0UuKHqX
4zRv799B6MeFgCZZ/2+GzzkpZ9Zx601OusMEOB6zzUMpZ++KU6qMK6ISyCs1H8maiKMK+HDgd3Pu
mUfWXd74bxANKrPIr+Y4U8qu5nwAF6GIbIKULDrvtNXmkwCR407OPHLbXL7ZJzDukGunlsDk4HGp
DlQisB1lhvT3aE1T9RJlcV5qSq8g3ZLr3pNFf/eq9sAGeAwaH/CEqWw/dsQwvfGZ5cuz6ojd8bA/
UviFCWBJk8y+d7z1EzZg/6vmbs11Ok601mvlAjcUtUxxCKtsB8ij29XMXJMNyTYgaFuiiB9uMaqt
zRklB6SwIvsbYjH7r6UcXFVATcNR6OK4/w2jLsHm6auxNrmPPe6iSz3BCbMI1XoTyigBBflw9nf5
Hn4BF4xnhhYDf2P34+8QT3SQVjw2Ft+66GgHgkrAJNDQ/b1utQD3XlhFGV6+yjA1HdaCw+30Quyi
VmYNqXcEfN4h4n5ntJJ85cb21i7OUanauUiYF20dHLLWS7YEDeGAMjoRNd5arZ2hR64Z2uk4HMXD
bCyhnaFf4hixxO2gCZ5pjaoEeYreEUNUg7FwitK0iVNXJr3sxKahrqgxifXBCuDQezKQJxsTlt77
0GVl55IajRHmlHWKDkuH6VrhwX/ntDQrFDpWWSKCKWAItBLtk33bowaQvRptmpwy4puGRC1Uzv/N
jd7YXBnhkMKXpKxNBr3NwM4BF6tZJCSg4ERjk2r6AsLjJ1iRLXoTROvPzIoa1c8bpv+aWggDjm10
QkL/DqSSxUHxL3xSQbCxR5qbRW8nR7M536ebhkEedlKoZkI9Gu3dNG3HiSbGaGgbL7/2W6xu9+/t
5ZqZsYNb/4kQowyC0cfHa7PW6RojM2iVOlLmBzLThcIQ851xnWKSrQwgndODYOZxNCo77mztFucY
+L1dlXPVy+HPBXmLPyvxj/kFyTien/8mH8wqls6UgorKE4te9gtU//OaA45lfW6tCvRnvdys5HK2
MUSum6/bGoCe497oGOya1fumQigqmyiXyEciCsb93NcZS5ZtrN9+4D/yEW2L0bpWI0myNAfKufmK
lF2quBTM6bBCLFWsqZSlkrXbiN5knL3pm6CtvxY3ZysOADlmmtaqMwzi7y4uHmTqWv7Y1aHx6tEN
T66p5JgArUjr47ktzNWYGZykb7vaw8D6WIxHOChPnjP+kz3xPsls51o4GEdLq/jSfa7yPKhkazRK
FVplkG2aRJn+gfj4u2WtjyJLEK5o4Jb5E807BIuWPZsCFos9ZCIG1Fvfemc681pTZRThdCT7kvPh
K7n+WHJ4kkRkLkVWLJXV5fi1u+cy6a7rfbpi8M5/P51j+gVX2cDYuRqEoFtEAfnZvW8RN/BU7PJO
+Eq6/heymG1r22lgdJjyiQ+ML9llsqwnPZONbRkTez82WeLHEHGVjRQiVFQZQkiAxnW9TvWfzckK
2nTYgIK08Pudec92X9pCyfH6xarNkgAgHKi4zk7ChmtQkkeHc8YuPGTkq0CwE1YlejjPZG2jji46
QuSOackwbcK3TDtXlutA56hgMR+KNFUuPglrlrfhXxOWGgl7Mv/niQhwrObNqHeytCinuCiC0n1Z
WmV6SP+5Dzdt5nq2kG+fAdv4FQYiHo0Zs81cbl0du36nJ/CpssWLHTivQmcKiTQyXPlsAygK+LQc
iZUFm9j7o+W1aiUeurXvKp8WrZpVa32V+uHbGCNo9fXX4rMmXjDoAwHzNixtncKjM0fXiNn5T2o1
MObogEFPYbBC/QYSdGAZset3areO/H3WCDDTFdkmr2NqYLYUCi2DdAhBFKJkdmgwFKEOCARC6dpo
8JyACq5NqcJJkgf+PaVceZZCEHohOi0izdu47PjBTgO0sK8MmvVgf4yYJ4cqBGNSz9qwzIVNxkQW
Xzt1MjSMAgP2VYKHgkXoEJSXTjzKrA9BcJ6JbmGpSuTXTKCiH405EoOoj+/4jLXgH9FmqO+Bb+/U
S4GZqIqqXTD7NZrvItYy25CdUn9PKedN+BVqSkPgLJFU7X8XCcnSS0VDtUyX6DzsAq+NAkJ6TXAS
Oy85yamU3JC4DDt+EhcgU0noR4P8AgO+Ee/dI2NsXCmosyxIla0gF9xEl4gwZR4BVd6EPeGQIgRU
6Iub+53KesKsm4g9I/v2OdXMXAQiFUkLZjjxCWu1GFgHcIdhDIJ35KguYiKOENXwcKNiiF0+950x
VfkmnRK2akbrP9A2HIQ4MHrtJYtpmxfGwdxIZNEozbhrl4R/9s64Bw+75lFZ6KuZcpnGgmZYMxKV
MoNWkmPnH5EykVSpzpMUoyFF6gpzXYzbXDHLxGRIYa/DUT4u8EJ3uDs8jWSTcnn+j8wD8fKCf+Jk
X0tDrt8L48hK7fF3PTZ52dt6+IG8FdSriymR6qFxuWNylaj7woy4HMQHrSwYeAhOq7ATmSyHA74L
oTORP9z76tPzd7LsSRokAUwqSPhQmyaGMJjuiWCYNO+GGLA1i1H6a7YC0hP3c8IZFSKmZUZXm0CL
Z0CFEuUd6lcU8hA90P7EaGW6QuDi9DrMyQN6KzB+HSTPKfhYyWrEe3VHHIHSM3FVI8o51r+99CdY
Hs59/QXpKxRZTkgaDxuFe+hnRW1Y9J1VxBM9cFDos/BWrT0sKyJri9Q3/MqvcRmwz1E95KgnZveI
TVcjwBUTv85G6TzueQDolEDHiSggTopKFVJvey6NixgjOwyqDnKnxePo3WTvww41R8pKGmrSttrQ
5iIztzk54kXrqW5NDTEA6hv5lGdkySW3qW6NkBE7ZNOxQboXOqSprioTQj0mRR5j4IlpEn7rDivu
EpjDYImdc6Zt11LLEskUachCIMCKTwQ1IzPCurpilm9+mPapg6OmkHmMB5YEB0CeHzzMwsnx0RoF
to+5Y/DCNBbj6aqaL2mEvaR2q6TliTFxp6dLFCda7/Vz0XDU2nN2iA25AEwD+NtTCGHUxuxGKacP
4tcCBErtD6KmSCvpqkGm9GBXSBMFnOjgAe1ZgIK6KzwWYNhu8XKyJI7SXngrmOkicKXcOIINGtgD
sVaPJn1GKvP4m2nkfmLYIFuKMX9a4EmBqm+E1U4s9lkFItFep/WLlhksu/rBXRUHWkkY2a1XzYk6
E3nrD1Xfi0Wnd/gzv1L1QsSa2g7nQmaetPL3ueWi7rzR6zQDd00NQTIPqvvytEQeI88SbdPskSOu
8eTsAWnVyreweebCvMlIlDDrFVpyHpfiGsD8CDwnVt9JovhMdi9T+2/9tG/Pc7/GzTy8HHc0lQad
f1KvT3UTI1IzRDU9xMuCOAzK/01PPtNPJyEGkLQkaocAHIY7zl9MX86kzsqUf5Z3chJGgXYtubyX
z5uoytYW04FqtENlXtKpPap8UxAHbZj5EQI6yDGRwSk+VkIoHcDtiD/Ch+6Yh7SKHr2sec83zbTS
G6i/SRiPulTfPZqrQmXHLfzf2qgv+nEh/7huc5dFdmMlvxhQ/hHROyMxV/3afCED6QnnNTWhKUGk
SpDTKNZjEaF0Qv7LxjHJu1xzO7di7Yq4hFxpbLOfOrVYvBpbEDuePBYqljiu0WhqAghbCLk4TVK+
ORMlehqRBARVnh6G2+MSGu7KUKk77nOubL+FaIVnJxzvKZNg4ax5wDeExOJgFiXrycxc48P92klt
hxaFCN1vOuD4v7TB3kq3VxU5d/rUj5WbbPrrDKeqHuTcSA0+qq4ZO8/47pDynSc9cYZ4iKN4WPAv
Yobs6OPdf1LVJiVTfTQidHzDYd13wVU5WNX1WIHCq//PCmFrFYgrbY+X4I6n5efU46iskfax3Bff
kMPIV9GcBmX1fruu7LCGnfChfEGH7Urse9AwUEvOSfMT+gm6tZP1F7pp1JlLfBVUsNZBUQMRTIds
UL4H8Ovmh63PYFyCaTUIaByjsRNfiYGy33DJztv6Ts2SJLsGRDfGCn0O8b0h5lP8LLDAy6Lj8jIb
37qSWpKf1d6OI1Ol75b/D0LTGeWZnzRiiTrHZf0nzCnrcpaft/+FVnOr0ci4BrX5Yx1SQq1w7wKk
G4Q2ifaUY/BtswfEay0hoJyu2zMD2HUwGrV8YRw/JLAJrUdNICcH1myy57jpTIOvKPDCRDodJW0F
DIVwn8WLmyjlWJMroVDoAO1NT3UEXVEeaQVQFQ4GvLpbruNEeidmEgol6hjEhi1quYIBNabjLpQ5
N8jsfFnatfaDeJ/5Ip46cUBwWruOnmkrGqvh3vO+debnUDu7f3qIcnF2IKcVGR3qANcZERCC//IH
Pm3xhoxuCbVaNy/Dgy/6EoWhF2DS171z8nIsMMVEUHNq98DDkiEoOtN9CKnp9vRY/eBjqV3FbqP5
xKhkIrmk82HcE6tPeMwvbgcIiwzhfg6zdASAtZVN6uX01pEqjMfZq45AGJ4A/RgEtFJ3kAsZR9KZ
qQCN/0k1Rt4mXd5UXi0xvpr3gAqyvCGm8/VRgX9GCod+PkEjbMQLL0796yqC1FPdmEe4zxlxdYO7
UgG/0ej6RU1x5MwtO763rnG1fDFA4A8qjZSMTlLaVa2SMwFFiqHWufJPPMa5LzBJCtPUKgILF19E
/Iaex0LZ4axpDj6bjBrpq/zXVFfPEtDVayjy2JmrZ4I9Xj8nVnNn9/wZ/ppdNZP2v/5HQAgBmbZV
9y/7CSfPyueYn3VdijoyAuhAdRw5HJkXh94i7TXu53UAeZcn9aeB2qMlBE3rXFgzrqoe+GmXglnM
6wDSe9AAk5KNyYlVLuFh0oSBKbK3rC0p2IM3sHGJG0sDnQ8Q2TXhGK9ZeqOeKVHQ9aqBB/N1kdD6
sQ6EZoq7tDHH735lPgjYJu0uvjM5FeMLqhafW2MBifR+ubF4ZyhL9LzcH3+Xm5uwJeMwZgb1/4Wr
NV+QCmHO32fUWb/nyNMJs1RdZF3k1zJGpfkblT1vmn+H6TPv/6nMpd+Sv6W2uJz6dXto2i/LpoPU
wTubrUTepWTW3jThlklagl42xMaRkki3knfUdyavcjlv3xBDBTUdf6Hr7t454BocEd1FplkPTTfg
j9SLu+IbwHEtRP531TOPu5gXqkRyawBISMowCFV4+lCBdNhUby1D7eKef5iRMI0h8w5eTbxX3GeK
N+3UA5H2bQK1L9NjkTem8fqPEq3BAspewUsmwmlj3hnt9Str7ONvOUmU39UbcsuleuIBNNQLIZ5P
GCNFCqEuCwC6QnZ/WqCgDaA3pY5NxZ6868O64dhmLKi1JnO35SG4lSL3qpwtgUkvtXbVAYPLzLSk
kjjHGvFDpO2ml2Xh1Vgl/OUjb2LU/CrDZJFssL0Ju6N7qRYhtvRRRrWpWRNLTgx+IWJUf+OehcXE
kVutKoxKLrJaWoz3dgS1jLOu42MpBtJhmv9qM04XZJMDqEbPqVO3YPxfjv/JeEdSh6OzM3sReiEV
eAo9eKJ2ay8Bfmjo+CfIY51DAvxju1QA30Xk2uY4AlXWpTSNk9U8BAMXFQmdGxiAo2lqZ3zoP+pw
Q29ihr2iXA32E2lUYiDfVr5PqLkSiDg8Kbe4kxx3x5s9+HP4Fcx6wKNUqOvbw5xZDp4NSjR8GEoz
BvsDVog2YEumiEfq9svoV1LZNxhMQ0fCKEpT+UuJVx9roXsAGDHFwYPBkJJrVWI0N4kfMqbj7k04
q5ZUqvLeOl6+65wwIkuqN61KBf969C/q+9I5TFtoCQks6k8KXNEU9yLPyh9QDbK9DSiV9Z3AaAHj
RbTLO6Jad/XEJZ4Ngj+AekHl9yiK7HkJzuGUFcyLf1TsmQP4VlsvGOfCSPJmqwirxIxTo0xr2TLV
reghU6KJ+A/3/lmUGU5nDU2N4N7eK9dz181SReoCNtX24O1cKp8RV1xviSxwj6ZaYPIWaTcj52mm
tdWSF2ij5UFyNRWx2QFEW0MhYaVAsot1px+lP2bytM8m3wTg1Y1ypLECN+ppDfJ0Ql+TlALk7/fR
AFM6GFo1V+UuK/LOPvT0pACHFLXIMCfU2KewZ0GpJsaQR5H+G2Z8qbr1InDI1Q0ZwsWHW3OFGzB4
8i9E1MyOC39ebnEr0x65p14MSwn933o+NokTiPT3XNdZ/AUszPmJgkf0wkBrBZf+vC062PiYCpAp
yfBCF1JXIcIzw2Emhbhcyfbu0ntDP7sLQ1dxIf7L9UDWboiUhFN2Mj96fLjgBy6CoT61M0Nz6P9y
RF/fTYiJFFeqReX3AIjoerrJZjVFHU9J6Azdb/dW+qimRN6I5g1LTzY9fr1A3IUJo67yhGZ2xYKb
BrCPnDrbNjyjvS00xr2QNQkWPLtYJfwVXkglcO3kGH5sJlc3SfZDLqoNXdXEMoj6LarRcyvkJJWa
pK8ceDNcWN6lUG0LDVJqpG3T+n4tjaBsH3XNoJQSmNtQocBwR/tYlT0bbe4kumcBuNOGOoFUsJWX
3DXTrJEuX39sIVJ/47+C5VJDae2j6rRFj8LD6smE4zyksTxccmJnA42mye6kMXgMr1wgIepW/b0l
F7qfH4kr5h0FHaC4oR7TJwARCdiP7uniWpSFYBn22Ox/77nR/AKAmgtgSSVh3pAu06SjjAciNimr
bSx15JelSfhN50lQR99cgGDUWg/+5HYTNlZtqrXN+vdRyGfTub0Irgtytg7RN9v8St9nMxkHwrR/
3ywxURFCUxeLKU9hlUVaDpUbfqJ+roY7KED90uJxn8UeOulpwbfcuRyGu2C4VB6xB7xgK04nyIe9
E9JUx++9qnFErtE8c3OZL6Do2tMi9WSx8PkTntTuHZN0sofePQnehQzyITBS4cpCSLfaAc4IcvJX
qOy3ozpvfNgsF1xlCA9WLLud7ZPwoyYQnB8TWOOSIBALg9J4ByPOi+EpoDBzoEoNCvbfDen6rhBJ
GKyIJcBDc0rOVLaLURWiURfxRcCBWzcoExQceggelQ5ByjvkxMW2e4VeSdHRUsCc75GwSZukP+XH
Z1fRarbimU4vcYlhbdcAHmiJk4yKTHs3pyXDsRmRQIpMv1MpNzLoPVoi29oSA33krN5SJO0gx6V1
g/Px1yR3cZH7ItLqHkugdVWsVg2gnyA7RgyIJ5fv6NCi9dRPVnyquChozTmZyvq1+JZj4NBtpoyd
0gFnwWS8VaTTDm32UatxYZzXwvxBH0IjWSbRS1bbpn8tUAHaq04Kf8Z21zInKZqKKoyqjhbuNIPY
i0oD/hc0APSnXVEHfX5/7w3ltdILzilFJY2Zg9Q+BO/nnpz8DHZygwUUy1+t1uGKz2vnmptq3UaG
3RjNofe4Q3L+hoeyG1rn3kpxZ7v+22W8/ZAg2zN1fVAHgAnHa5muoTvXVuZOSjWso0Vat6Ie9w/O
z59jc6FW/Bz1s8txRhoKmHbJoCw53Dj54bIswwusryNM8IGPmEnOCkX1aW9+vnaSqwMYTZ/juIZU
NHgEGFQEJssyG7RVkOWJapOIbTf0oqWUdbrQpuY6gYUEWHxprrsrWfPFvLbzIzIrYXqYqM4gAgv3
p4FMPeUg9yvLZJ1zfIU4HJTiw1EE664KicMfQmoxW9vFOOAKrWhK6tcIb+VofJ99KDRD9GKy+Ss3
bXR06nzxiVM2DIboTIOCQ0zELNgRJiEnoNwJMOH70bssNbw1XhWsXUlNwNbJJVcQquC9pUCwhX0q
fc8jmp24u4W/qSa9QTlYBioE+rFzCpngcC1MIji33xS6yNnQmNbSkANTn5jrwFztpstQlvCtiYl1
kMaEN5P/ceXXUNcmVpCA89g3nfwbgY1Gaajg+9KUNcx5nQaJGrieaq2ljXBkPOj4qjdydmMh1pIk
DZqcTJrGMJ6R0Kv1SdTPOn+jGjLfSX/li+MmGGX7irztguKhGOdGguw9bW8uUP/FKi9w0jZT1meQ
75vbrYlszZnAFXFax2Llvy9d+8mla76Icg1yUt9drD06I7aDfHGDxhluENmWQ0Bl+SPpJ5c5W3m/
DA3hCJepk7LuCiv869TiA/MKfINDXQYIyadFKNX9fICc2H/d0FY8BHgfhe1qq6cWdjX7SPgfks3g
t/4VYy8W/Q7YymonYYNMNNCuWnci9QCVmcrxXhXgY8u6MFhG1VkbjQ4BFx15Si9QMBZP2ZY+JtYY
zAWtrdRU8Y18PgRpQl0rK4THNeuPymXF+aVHa4rfTf5k1qCCvvEE45HuIe6gU9zUnm8v5aw3NVsu
h+HqlyBC2L5BiUAClXYDpkVWP8hh+YRC/RwUCPxJCDMoNU0z2ZjcPNyXotj12b59WOrwB1mOWq+n
nsKlmvqbQfq1z9ocqu5mZn2winrkTNLZ6Aqyls+ffna1nNofDTUrYfeuQ3/eUgT36sdiRfCkTO0J
G9JjNif97TQdnRtpFvPhAho5Jxgx5qAOAejGFETsb906LJlguaz12qEepvDTjvEvU3Rq01k172zT
kHrZhNUyis8bTCWj2hbcFLfdl7Qv6TUXRv65zyFs5hfTkuVyEnkvho5PeBOlthBABEZIVYQf3pAd
WpjgEpQrvbYzf8r1TilrLpUVT4JBjc51NWlmsMqFD0851E+T+iSI6aBLrjvIkSJ6TMNQoj+ux0+r
GSLA/MIATrCW0yNDNIKkH0GfUpcdUHMFgO6DKCCUFqM6ZB1+IWR8Tk+wYXi9rBlfhU+Rxv4KhysI
MWaefVGRoLjZ4FFTQeUiwqcpWJ/q39NABFXW5e+QdqkQ3mBAChkOA4nejTZzA9BBtplbWkBfGA+E
4QaP+ZTGlmhFVffjAMfElKrjcloM+fZGPTcJhEWu0gFkciM3x/QWj2ubkeBEQ7T5PBMkOMbhJTlz
guqVJdEY+zmQos6lJ2V3EJtLaIGztPFtl19unypsOtMDBT5Xthe5CKvcq8q4AYLNnsN8YEsaos99
YaDO1UTy1jCzzw6g3s7mphxQxCA43fr/cWNei8EgRqaEp+e63IW3qmy1QFQCE/Ir8J8I7LgualIB
PSPQgoTnS7JTQc182N/YYTTG09jCa7/B5GAyxHXLy0rnLg3HHgUGZhwgEG5wLrJJgf2nxFsukk+M
jQvaooesAODlNX4eEBZMz/RJiRD1WmZ78RSzMh0fmKkI0FIOMhrQp87HiMigmHcnjWuyerBICNi9
Un26D6DEy3vZnOTjrIshuosUgRu9AD4cnD8KOT0/+KH76yYCh663gKR9YmQnEu8sstbt/4mfaoIb
HLukZZlJIS1CDaMnYshZeLSjToNzzc0qOzlk18iiy8nteXAImfsgxe/SEZv+6+COxMhs4XoDe3nX
M/qmgORlUpQokDUVe+Jfq5eiQfUYcBgn+gz8z00FZjwBXhDUnPJYZgxcz8QpWLYMjKobJA7gX4VU
y9YE/bFSATdkbgdBl54XubQspsjZc8kXlqUurhLKYIWVzSZ2IAu08GvNYZ3EoeZDoPNhCMLVgFpj
hSzRz5De4qxl4uRkdEl2wcHVDg0hWllPKIG0O3oNWhw0RB73GWQGqUexqBgnWLWH2NjJm377H8A2
/Wwpcm0VJVCum8B8nxIxPMbFmXexQBj8ggUQm5+URc/Bo8K3t+HK4/Y7wixjm/pxG94tYsaqgmbe
KVNCLJ9f8K2CBJH9X0TRxgDBs8yYQEVf1QW+yjtCwTeDHmBTCjsUo+zyPEhXvKQUYb/133HPHGRv
U9U5ckvS3FMEOVxC39by5VXMISNZ4Pz69Aj7aVW+UISXLeo/jMj66Ls6iX1HjiF9T3eRa046sejh
4cYWgvG+22S77t4KV6TtbPjQMYnGhLdTfBJyWe/F9m9JHBfZzFolyHgi9+EXT5ctxugmVJAHCSXe
PZRsZ3ZImWOONKvpycSLRXo1vjjdMtVwSPoiwLVDxjtKm62BOupG7GN0KpgKxiean+hc7wO8j8co
6ui/AbPYupJ0RdrDAW77w0LkvFI7h0V171BAkK8u6FWJj5lOkQ4Pxlm+r+B1zwNH6iF3n+2vkkDf
UGrHVJFKzDTr10MWYKbAQJBTNWysjOJiQmkeFj60lv8mCGexSlGJTXYuuTaYm6VE+PI5cNjJqy49
3JqJ2dQhO0oYtMY1qXsMqYqHNeqlNN3WJirVu6lGdnpn5V2bv5jC3ncf818bLqSKz7oGZKwk8g5g
3ttsVq1LF48OgCAGyV7occf5TrdHCmaK3TNkl7StDOZ75TYqunCEvGMvjR/QxzSgLinCW7h2nYat
gyhxqp6j1qfVLCcby1yQmds8jjwcCJM5JyEiCwIMmkSNWTuyqd9S2oag/z65zfBUaqj6yQT9dYsX
aFloMdBq3Z1HcS5V3dojnVyQ+4thYlQG4JJWLk5gnWG8UGm6WVcNRkU27Gqyg/N1EnPGXixsLlC+
s/dEjh3ziI0vA8O2aw0KCwmR/qMhRF/um8S/XZiH9eYqjhd3PYS7rEQIgwtiKxcITOsG27IEKv5n
IDKKPoCC2ht+9qlTMIgs12P9at9CFXooP/vBAk73tUq95LVZ4IhTEsZmnyMTopJPuGUkemYDpRmX
2PkGBL6V8zJKWmGiNbwY7E9GiQUIezjvz/MkqIhSMyImhJ9+BFJwNE64clS+9bz6oYnWPZJV4ypX
AVAt5kkcvcSP0A+JpZsQt11sEGDNNifDq8Z3wi/oFjvcJnTEAdmnPESyS+Mj1xg/wCtwCEXtHZe7
8KWYNROtf4OYH6BfA83L+/MdUq1o+jQUrosrXPXBO4iOqnrjfLGuwE+e1yF2O+++mKEIVdbquc10
b14iqAMCWZOxyL8GLwCTkaUEa3QbzGkfOSpvRzPDOmD4ZVTm6sxivLbwOhTzV6mOVq/Gh8t41YE4
SH5pPlQfw3wl4xill3H4Sxk3Wpuv5kCc/ybWEZdGlzgVjJqtIwlOr05idrBnEp8x6EgARWauqT7V
iGCOVRUPwMkhWuRvO9sVecqM6lqov9+GJYMUYvXUHL31A7P1DsdCpTX4xNhd+7slUqZI+2yl0F+4
hsjo3lE7/41Tmpeanb1BkFYokaGbMwTrVF3E3yEZRPfYb2a0BIE/DgnDJzWuKpXRjH5BNOXcxZ/F
QUaO54lpe6+6rL131LUQqqf2KE60fvfgYYJIYKhXz8HX7iXGV/07aI+vMq579WJbeiclBrPgLIkg
KPnZh/ufbU7A12NBGUWzuLpcDLfFrDmX8cc7PlIHyIXWmEf2axApcXEop/LV0evgfCvB8auveeg1
IRdbWHNfPMaXSRqVBXxczZKTn8PKe3d7QWLGF4O0DdXOu5Xc+n7GzBmm61LqFHtsXV4+jAGTj7+T
dAathvGlhvUmtlN4MDVte3o8Ub2eC+9/dY7qnmECpVKBd3S1oqWb3BzpgTnU6siNuePmyxquS+AA
zkZKpRdXBCuDWFunbg9tr5t0BwgVPTXDCD/tNop/qdcNwYpO7pFyqw3UeRam4Wz7IMIPEC0KuX6F
Q8aS5gIiVXfW+7YnNZg2ffQeWbW9Zi7h4TsAxY5M5aLkaJOHQYD3KTvOoCcHpzbq9AADnR21FWjp
48BDlkumcZGWtxMHRKWxK/9omK88oW/aQSVaCx9ci1AqF8QBUh2Mrt/wXHtXouZjvZYH+N4zweJX
QXvmAu8Gi2yiBz4NRhBpJccrft5iNkCx1/OBk4m0TBqCFrQnNFe3bmwIq8+xU+3nQQ9OqZJHIJOx
wy4CrmX2B87hzUHcyE+U8iNXNZnRzyeYIoTnWO/+kyMVGGuoOGp/gZK5bx6cH3SQYyBN8c0bPrZN
3p1AYlQ5jJXFcmki7ClBINuN+rNavbcBP2s+M5+e63mWBUi3nZEen18Ysy53onIFvtE0ibXqBCNq
oBdCLzqaEHi7T2CE8RFAVvZN80D+71rAoWMBHjY/8TZjPExZ+25teYwjfjwb8g85o46tjIvTGdZQ
a4vhamZ0vHJVOz4VO5doFyNqQ0mN2TYZWJzGDfff89iwkdK1LRfBMsZ1vuePW+0Npl3XpULFUONf
Bu8sDCXdpsnHPapYqYsSQA9goWR1Dl0bLqcwJzQpV8EtyCrNFlTeBHkStKHAJlX8v1cWrorUHTKR
oVzoICYpNUDbT3BiY/sEZen96OzjtW2b/yjjMBi2T0zmkTxFkxekwVxxPSopeGF9+B0CHsgW1pKj
WguUa761tF1vPHhdtvtFug9Vse0q4xBj4zFHZbGz3YfyPVF6eXqk1jBII2xQ0M/dvYRuFGmc8FBA
0JtxhFs++R0tMdpmidTO9zv9qtQ5QdL0bhIzuYxJ4AGyoJIQOvTDt+esYx8COIZA2hSrmjcOFCR3
dqp6rrRRI9DpRQXdwMH1gDApGNygkqf8MRVN9taab1hnJvkxrCbUtV6WRiKN+qOwhdpbiVrVuEXb
bFTwsu69CM/qlwSNS0oTNVSzsKnutxHRyV3YraoC61YZB3MLhewfWVgfMId31pAXY45Zl2b5N0P2
4fmYGwfvU1Vf9Grtzz8PHa2YcL1sRJKaQLZJ1iPbK6QI83o5jGlWEIKxznYEdNHSVpcCLldeUcSJ
ceRuOywo6j3Pkt1zZZLvniXtbxZQWi++DlUzdQd/c9OoHJHr3fAg1FEepGwqt7UJ/gYnzrRdYKMs
o1FSAA3doRg0wtyKMVJyEsba684oWBlzXnXDjK+7aO8C/24dzpjCKzzSmKjJ+1srmyEwIHW9+aup
k499lEDdoGZkCgl+u0UOX1wbQM8mOCOaV24j1t/wf2C7lORxibVC4KGf1XZwBDZf9TBf0XST2M+F
5Pqc6h1DYzwcHtN16NNp602uIdzcl8dgAiBYl0W/cFwNAZeZssCNSgAiN8wt5CEz5rzgBmQBXAsY
j1GSdTbMLCzA7YSCb4CN+b3RJ7ildm7y5dTtpsOzesDP+eHrOsnyj470DpdVNoooMrIUpTR79rYT
czrQxkmM+Pu864liwEBlBfyv4n6qOyIFXDaYJJD1uA1UIj5xAYGhgHgY0Dl3glahsAZenPHgAcFw
8M3x4GzjQZCuHcZyqpjaW1ib8xUSPfcls8GP+TWZmdGWRj16dCAaAGaHwwBf3amevgZJxEouOszG
uUTOBpNRiRZxBeGdvbFD7mziz9Tif0RCS9sNzCe2PyCZd9ZYT1QeKU82Rle/Q5KXXxch8wwKrveo
JweOp/9PC2XkfZ/DKukW8D0z2KfWRRy/CmZGVX1idHEIPNaSI60E3UoAJEdB9zLrj3luRJT27zeH
0sN9AM9JScZhytjGPpMEr0tmYgB8/5J4SIUj0AayrM6mbxvhwYxUkI/vcAXdtE9wcwBvEwcZg/IG
h+DexiJvARODiBM1Y/0q+s74GPp/17V/zQY7UzXiHfKvhAbs+hlb9WnwjvNzSd2SX8CiCfyR6Jy5
h6To+8Q+kCUYsftxNRvJhxQOa5bOKLATmkxx7C/VpJJDoLvzYZlcDcBr5y22pY+hbEIEAsfFPgPq
cupw6TkM2yWhSYg66MlP4h/GyWA9cMrBO8dpoCd3pWs4yi3huQ1P+qNE193gsGD2/Mf6ZPj3HlS1
oSTJFSB3UVJyu+Yw6s0WDnG3Jr6pFsjY+QBt8WOHYGnCabh/8j8Pzfo1r/0zzov0b1RhTOQN4TnU
aTBMXgELQImJy8vfTBMlcDwzSMte6e18/VuAycOkR17VMQm5337qrytXXNmIXc36AnxEWISsYnne
0yfD3qZDTwOom91PayaJrhdypoD59qrYaBsEA8l6fImLbWLWCkyl5EbmFKN6rRuAmlr+5Yb8LnLI
kRg+kIm60TlIoKgRgEKB06Q1+w81DT0l2hn+W7XXvXiLzxOzXmpMhf6aYLG63T4l370fGdXhG+n7
/CGLkMoTmeGB5HKi0+ey2JaDncIw149o1koG0Ivd9P4s3vAMVwu0qil+M5QwnZnLCEBjVoHIG3T6
OVq1MevC+yjs4Jf2Kd6U22B1JlORvuJuaHiWmxvHhh8M0xJPn6ZKOtZlSHWXyAdQGCFz4n02nhwi
ZAOIlyoc7F1S1aGqjxuzu2O5UtLPwPPnu2Cf7S8+9LF+6cmrDq8+ibfuMXuxv6AjMGu7lV6Jnx4H
SsCJCacxZMcrTDk/DWDXwajyHNGe6DRVBui+mVQsYKLk2zGJTBX/L/OV5Kbk3bYp3BKCkNtTkZxU
r2BruYgxI3HXCmMyHTZz+spWf7Fva8UUFf76mShQhIUs83e5sgKW26n33HL/zVih+Crr0QURCKGC
ryZK9sHxD63fmRkuN/suywfzjMuV7xXb4iQZIgGeTkQtR9tLAG+IzRDoBEIjvOhblTya9BmIigua
Q+fRItk9jefoh6/nArjH3B6OMtgWxfhOObYA0swR1FyZFFCWETXnXo320rplWr04opENAavG5NtN
3lPmUCjFfObWrkrFK5izsD2wPrwSch4D+pO5GAB5k3bGQJGsRoEt4I1PZBr9zFF1tUdy5RPkHERE
OVgAnK8h3b+VwZsd5XLI5AcwYXrGc4t0KOKB2s5EYWQXvAh6yQ4qrHeN0Zx+G1FtISjasN9BHueJ
qG/6UmiA7QDTMCMpofB6F25w0DWY5XDhN6aBAHMP8slvif2sEV3NeX4YUzWsCRTpTv5qEWwy0yZW
sBkCfDtKOUi3GIwkCocWLRmXF9DPu13MugkEQvolMOn6cQgoVT61MbBbgL+MdJIKWtr9x3MEU53+
lcTBly16XAxaGsS21bXJzDZcM1jgCqR0cwhkKqF622CysZXjgls7OlicYL0INCqx/tluXZfNdzYY
iJ+1g+/kTeQfEDy9xroPJrZfkGhR4Kv9U/hxAIMLFKw/hm8HqY2GMTRN1WgzqDRNhp9e8PIB96sk
FE5K/tWPHczWJROwaHCXmQ2fejxILEvw75km3Hz2nJvB7+5ZOogagyoR7l51yVLO16m+6csCdork
5FxxaAeACqXEfrNsd8x6HrKmeOz0y9C/JWeqV9twAhS2lfLYDJoqraAXpyViYZPDFLcTQBxaWMzC
pFQgQNi09AaPiSlbRExVD26i8uN1Qs3KrDbsL6Kf7k1teOYePwKzmIeO7a9oQgtYLvGZa5qfhB6z
gQuH+/L/ocfUaVKCFaoQ8PkXU3LuCDy0Qp8Bo4qxVWk8HcqPqCuqLh1JyM3CCLBoUEVMM9y5mRjs
3PT4GiOhHw5wJWsexvd71AL3XBHe1KTGUG6xuoTBVVWIwQfaorB3/dgdIomteClO65EfaxWMp7TS
peVjxZ2llig2KWv+2+9c+Qcm/GlxkVfJFRxG9eMiD8PtRxpLjJPrgXptm8Si/r3GuIIIeYFn5BLB
Kh3V4QTMuM1kV/tWgwcWg7VOTm9XPuqmUaglzFlKfLwm4Fx3n4OiyLbZYO9l0fG3vwhQ1dICiVsy
ecyWfGAwkbU1unPkPVI5AW3JMjYfpVLdY11j
`pragma protect end_protected
