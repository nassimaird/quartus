`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nDJqMF1+ev13MCi4ZSCdtJE9Bu/S51tijI5JvDRM5Oy0UiehrcU3wyJNGp3uckeO
TPYhgHR1VXQhvEvqO7qmO8wuIOtrJ48oIbH/3RaGClBkRSN3qmefLjlTn9F/rWJk
ug6EYaZi/bEnFo86zZeIFZEj8dlYrSRluLV35dAfzU0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5968)
ekaIsZXiLcRc/dIWGhD6eSmdCpYwtk9BAr8644iTvnU4oN4XPqnfpf7mHYU0WgNW
Cl0rmx4QabWHEZs5Sh12i3aB9BYC7DcyhaGfhi8ZZLiQXDiYSUahu5XfXuDWgvtF
dMdR8YXCA0woTCqYh5sTZdkXSOiVTcaufsuQLYluJeh92OEQL10WLZxK3zaxtJSy
BxuIDTWkntixn6i/oCHr5hRm6iiZ57URgX53+C/8L5+n1DqdhukTbaBGTB5x3XZZ
QpaGGcyZJ8pOCilfMDqN92TdCGMH2d5ffxmfq+ESuzpymf0q6r5FIg/pWQS8JUCD
xHrd8kPeVVzwWqSYwmNPdPN9tvjMYSN7Wo0VhrMhhhFtmmgzVv/6Yui/0sWsj1pM
dMwYSt5BDQgcJ59Ge235kmFaGf+l5zheEtPzNhdBW1X22peQni8s6eFurLr5sRy0
hznfOj71y2iZf6GgVlRITEeaeOKN+ou3+gM2Vy3NT22Ri0/SirWD4Ci0A3wOXfnS
XmqoFnMNSwA3BEPLjEXKuicQbKbpvDgDAmkeFlfaiXkwubWfGuc+uwNjeQSL0AWd
Uhfz9E5K0i5nZSic/VS42RcJSKDYa59AVN6YYSORWyMlAvSRyCx6UzFqIYdM5cEa
AC7tQIyoqRe9xlC3DBREYrCvrMB6Sj/dM5B9IF/ZZKN+jAI/QmADNAg6Cos+spTF
we++lNyX7Gxs+kwedLysD1tqNiVGHGFHy00OgzxZ+W/Y7Q2zp1X5Dp3ADfeg64vR
LIQCuviyJ0n/4FL8myb1doootMr01E9ZeIk7OSmxY8HmwNRLFDjgget2lQEzf+Ck
LqVHwKbi7l9o0O7sgZWtXCqT9pupo+FMlKP/ZciIUnpwXYOfLa4izI8206R7Xs36
SfwAoluLqy2ieevKnTcMO/9RS+fwCOjgDZfl2B2Xx2Dj72K5RT3Ds/3wUt5Sk7/H
haW1BW6ETRHBWgMNl+XEWOhURRE25bZAluKdIQytDIIelpzAdAm2+aBXMUJ7iW8h
MlQV1/mZH2PyjOKga6sLkQgTZZyZlrFljaSicpEOZ3WYh4xOuUbGFvpaFoDrSqTD
n2C5WbTiGeq7hGIHIHM24M9aP/vo37xW6IlakeSGx9D/tFFcX78uKTzKChf7i51S
WkiisGbCfG5uVTyKnHtTgf3GZpoTVTofhnBPh5SXvfRDgs55I/gQe7dCGtTNFgTs
OiXqSaQCVVFMBRkbOVgVGQE3ir2ArW6RjpnZdIQkH4dzUbfm5OuTyjVH/SK8mijA
gmE79c+pqCNJzVmv3W5qElM2fsjUiQoJ1IOierToAYIc7TgvCnUZW02gr2BX3O0b
m34PTiVZfdfvMWr2+CWU0Wchn+DR8O+gvVTGsSn+Xr4nvAzJ782FxSrAHcdQzM65
83sftf4le3oiJ+RAX0N3f7iJJ62gK4QUjRcLRQ101MtGhDQ6N+QDIVxWYySXy9gy
sCpOFWgKpf5V85MDanYXy4Q/Roe/pQlykw3mJo2fGw/hVAQi3LGNnq7S9gFMN2rQ
y1k9aHJldvUud5r8ouM7jCHfQHEAc5lIj4mdyMQECr8SiUoIo/mHauMkfDC9NKno
iOFhCxg0F5dUzQcdolHaymaC8PfGfZfJ4UXmxCOb2lTvytESm6d4TiXoHtybCUez
Mtr0CMOp0a6eE4nKdMql0QNcPOifZpKahAnDaVc9oJKrmhsenGWwY8rai7azCk/g
/6O2LGERr1rhs3JdKTUqgRgl1yMp1E4K3nTxWAUORYLpAiMgUsBe9l+0Lhb05jrS
To+X2hhCG+yWc/0DguVNRiiH5kP8l3jjYdnyEpuROl/EJ8FCYkEnyiLl2kJ4CTGt
VsLND8FGYz9/EHPyIHpI71W7IMGbdIOCP3KOI+PKzTZS2e2zXbuESEou6PLp2ETM
7n8DwQAX19rTBlXwTgIgIJl3vNhxiip6ySJVWVsBnQ7waw/d6sO3C7EAuhOVosyN
4K/UBLTHHc4PMW+jAN23Ty7PBdCL32iu8PAwpTVDE8S4CEX7/vFK91Rc0LtwbjEf
xQXm3MYmTEfXpY3bfvjHoDJ4QQlCGqMGdpdYFDW6B4Q4XwZfxDkuPiOBYGaPGMFJ
UFDDKfH43AnEuiUTFtwqFaCe8Vpz0YuDY6nnVXusiOVOHZ3QrL4Ihr+fIJXFVPhC
EaYccPq8Tl9cjLTST6+lNVE443DGVrEgA9AH3eIeJN4FYIET8FaPcEAlCCzEvhDP
lSMqNClgcWL1fp8VMSlIq9GrhmdAoYzWWBxx5nZDcvLFRcKFgAphoJykwQCdrx9S
vUIhEXrgyJlgAg/264BHckxfdPafIFETaJl6DYClwC7W0h69/uKkTgtuzXQbmAby
FrYxdyWKQPudXoeO7au02xQtUyBEaZLT/MIxNnK/kd+4QVTgMyR7Or9H4J+MTwi4
MfFVKnPNp3LfFluTEkhETDIBz7bE4FUX/GqbwVde7FQ9AkS3+0iEx3868j0PXFfl
Pm06qsZBSvRfrmXvi1H8RiwRLKN7jXEXb/52PAfvtG/2/558iVwSJEnJa3JxIP3B
/c8O1NjXOHQPJwLjghOqIiUyRvg/q/bnB72dIAUBYRf/wefQ/dYvl6mWlhurRu6e
pvIjg1IfGmkUGn99fthnkK0Lhg6Nj+japqqtuFgvxkWooNrnzM4t13JaUu7nbi0Q
5E1wvHwkgNo72y9gIOsAhoiY3eNriMecsrNRFo+sLEBAJvjcAod2h5H/U2BKRJmh
MuVBxHdOlDaG03nv7gQTNd1FZkhmXIWCP+eN0e9FXTMJk+uZ+HSosMwVE3S0hHoK
XPdVxO3/Fvb+s2UAMsEO2M7WBGDXPLLTZokF1m+PNHaK1aUAenctW02sf7jKjw4n
wvUNz+5RFMCwU9xRQeaeZrFRsABUcnVrQC8hjfnnGL9nknNdqy4hyFF3LwBCHMdF
juopTvzMSYJ83/q9B7xtFPp3D8HP9hvYLl0ygcA1vkMjR4n8YMs4gJaWnHaMW8O8
xplIzXkmBhmXxpgKP7yuQL2btpDA9QxlzXMe+FwiI5dpg1XFe8OSMQcx3ZIAEpxo
T6qnE/PQGM8mIRk8HU1Q8Hk710py9fis6zXIDa/rr2geoINU9PreL/h/yDH7aRux
VwVxsuw+xm1bAuFLlOj/90RgeEWUeDlCZ6WHdOxmXXopE6wtOCF29lbqUXSSvFnR
izxeg/nyX/fKVbk7peZaWGUT9km4iXDW6vvaQMO1Ww5LeY+XoRxECtaWt4paSY6b
X8gqoDNEpLXhvGNB812BuwcA0ToSENpecz9Ra0lGj9zhlWHNvAgWjVwN2GreSoPN
/Vqd5jtR912GB9duSzQBhd9kwIYvdUlB5DmUm3j1eU31WfQxU+HaYz680ZlQJ+Pa
jAaBU/56iE6N35mscUii9m9LV8iBQeZZjVxzxu/nre7Rqjmc5LtL83bmdj9yli8d
3IpkWbgJRJk6/9B3tum82oF04b57ObF5XfB5t1oLBP9Y1sKvb3bd7a+AcfvmKLln
y8XKfWQIWnKEQmjhPPEjwckbD8OVTGHwT7h+4FsGdHeubf255LDV9zQ/3OdZOho3
ALhfwMkbijL9xw4TpRh1ug1iaHPiO3Hri+0CaBmNgSxNV8YaYwW0Lwm2pcdaWWGD
mUfRx8t4280rExkAssbnMA3Z36Nb87WlnWtXBd5z9k8Q5+zFmOp5WoaOS01uLk10
ZsBxdDxhyGx94ABkWwcp7gUXQ95Nzjgv5Uuu3umzRYxzIcDmlmISInpulhwfkA0M
UBrP/SN/e8NnRNQmijW7d4eDJuiJgk1qajGQdkieDAdAZKLTwzdxGOciDDGOJUQ7
CQdLN6Z/e2cwivgbdFW0nF5pOKElumZIhWImiXFVp8x2gTTJ9ucO+SeEmkZmLSSf
h1kP4WQBgYeip0/hlOVAIKPHDcxPD9spDF98AToAEYI+Ytxjrz333osoP1iv78An
j99kF8ogtsMzLacmd24aXLjHwXK1PmKeuvv44Po00VN2v+Yihuhos7fBz7Vqa1ai
g/2OrDIvq3iQoT5Qo7bnk0PGnkRBwMh0bdqkaUQX2UcxxHvUN8/yUsFvysFK6Yuj
KAr05TAvU7rEme0r5f/x/p8Gn4g/1i3a6uBz5yXhIp0ta20LwWT8uDuyjS9iq+nk
MpKbrqOfu6UJbPFlpzNtnx80x8cI3mKbrEzlS3KDaPf+/aaCW14wjkJingsDm7bt
GeJjuPoQrqvMyM+ZM5ApEMF07JOXk6ajuAnKt0eYvJ9YvOd4OM0QqAZOiO92Mfnd
iLWVInFO9TInktLyuhq16UsWG8wDD7M4xNBPBMTNFb3fzHQptKHceYgowQbW8XwU
atsNk5UEBhOV6UWAPQzyT+icXNeNHl8Fa5lGs/1Tnbl5mhv8q9Covjl+Lyot0bZp
/HtgcZVnofxjCWOa//TvAw7uYlcdlW6puc0GJhlrxx1/vmz0cAPVXo/0sUCbuwP+
2VrPG16t/p/1ir5l3NitJTLLF/Av6QEpPw+l4xvvPuixcRWzxyPYoYtgOlScdLUY
IMB0BkABk9aANEF0erb6JiafIfVCjEInnTNlh0Le4QiW22SouHzINnT9Eqf9fbTX
CS3Z4YpvVRQ94s7JXj9WMmuT5rAxmt2quqQFGDWlC+D2h6EOPHeTt+wLZKfzUTKJ
92VE3LVSiSqAUL+aVUcJjXu47o/jea2hrHDOw0UDbxDpjToobBEkGW2ksxpbXCa7
+gs9nYyIVPL9s5ov+cLMm7l0sTpCvVjt/oGymjai/JgWGz8vWcEsuv87FO95Ozsp
Hc/vWnJAjyu4alRdBUsUHsauKOm7r+h07XAKYAr9qpxZtQd3jFQDRN9ZMWDKUA+a
h7T1Q6V34R5cgj4zb45cfkrbldOxNw4sznEQP9iqYRF9UbtEnsXCHLWj3YP2vxdZ
SXQbc0mo0MLKBWZ71ZhkCbI6ZN2ezWZRCN0+PhariqnjMW201Rv0CMnGTW/x2qSC
j7BrSNJXwQm+wm29dzEqI9Kh+3Rqu0HYpUjWXC/GY2dggGZv/2mRAsRVEmGo/mdi
1YN43cugK+cdNJqrx+jhu9haVfSMafaI6pGjiljn+4df1BJIWniw6tH1n1NFZlFT
uLcU1DNaQi0WTOKC7IsSajp5LXXmi4fhX2N/qCtSg8D6usWyLhgawnS6uvuF7hmz
DApQ6qoqsi5JQS3OGgCXIfkDats07VmBJ2UUmpz1TFOpjGBbcaT/mQCRUo/2PirI
mb3Zb9UIPUElwqOWxocDcmGT+EIia4oN6sVrhY4srNhPLOnDu6/Sj0XvSb3yjXiw
M0AWBDjaSzieJLTE4ZkEp3Y6StDlPlpggxl6SOMGXbBHpIaA3W3yHixBoSS+Qo9q
yPU2gy/SM4AHU1vwJlLt+anlIQYdBKd1/9XcRQwaEp4+XcHLcWcusO3RXGrZCrZj
6kGafsnTShJBpM4Jq9YGY6TrpQ/cJPx96dgw1emU4DD3sAkfqyiDkNv5oVu+f2P0
XZNNw17W3fx4MxrCQY1yngHfGm6lG6o6fwGFgEXSnfF3/P2kk3ecglXTBp2v5Q8G
B9Lt8W75GDnNvDigeEg1/Ue8mU05TZCF/GoGdSbMW+IGnhsqgBcVpPhOIcGIKnnH
FA1aORW2N+68/1qNpnPxZ6g4eg/f/+6cA7iYuhZzZplRO4z+GRMmmlZ92FQEbuOM
q1txOxm/zsonvSw9851H4uu6pfkMDAKlZc+6P7ndt1CB0TRH53dGfiFHwXEBFRND
ZgqVGDZODPz3Q3JTRyTUptKeCa2hf+++A6rwM6+Vs7PCdELYz4c51n+Iqm5oruLs
ajvjFd+INJVi7EahP5PAKTKfCvQ9CYAULR9DsXYgtbljcLuE4dng/QL50yi08GNZ
GqUykVk90ScMKpTJ3WLrDre/w1i+aXCbxP9bmUHGJFPRzCRO5UaDxE9D54gzT2M3
LLo8URI+EXRtA+A1qxKLG1JS2Eiigy08rda7qEQGssQpSwo4FBBFQyLeR5Qdwwxc
kgYkAtTIq25QG1rRjxUiVuGeFe20LayERwlLpelnc8hK33DFqPj+OKSRrM2RupOS
e/DipP+R3G/4LgxKk+yq1BS1O3o8EyRYGCXr+DNFTYnD/XDK8dL5YszNy8Nn1pMT
qli2Hb7KmJzXpYc387DaDezDoSCAHAj8d034PjFt5ri17Akyjx2bP/IPEMSKN2ex
9dvHreTM41sugrDlaE67dlXqqNcl18lnF/q/+GfJ9TumGiT14G7k59TYy5zxefiw
k2cqN+8hKGxs7sCRMLY02hOqf2AF/R1AcRHhVdakxbivpqmPB9sU5AGk9dsj21Xc
dXBjwFEHDFT3RVlZuxpOnzSu4MkCKqhjUD90Nvp/F/IoGLtoMhfcXQaJCm24Eg0v
s9TlnnOQTkpa6l124kQdTz9+Pbxpknt5z7OGfmwkA177r3tcpa+KXfbXlJ1s9xlD
HLO3sFVrrs4bkZqRDVPSSNHuVMdYchbgtUlGvbVTHFJHF7eoXH9QvyiM8XuOlm7U
LkZAwko4Tl3oFLJomXQ0zjU0WzoWAyABbfkr/socrZpgr3qk8GYY0pfnwm/ghryF
jTGZn+mRq3SN/lZZyoWWuA36x86nSzwPXOOucT0FM4ycZ9tS3DA0ViYPB13wqS1d
CO5ZUtQ9fV/TyqI27E8v1RFt3q13pqX0N3njMYSwAA92yXAsY4J16uDgPEEyfqVa
DBVzW1r9saPA5cfMJCqGC+E3ayepNbzNHOUomhLJ96i1JYicldyoSjW9N5z9QgA+
qCCHBfrAsQXX21eMI9dd3ekZ3wRsGsoU79wEPPXKaBhCLKkBZo0c2+jqwxGg06D/
GH8A7ELfE8MzTPTPKuI4xJA463Bkhn8ruBVO8sjkmrpVki8a/Nkw2nJ5g2eU4usl
qlEaFAeUQwszGzsiwPWMHSom2iPyUgeJgNdKHST6d1TF0CR6x7RuPbcg9owA+XBh
KnfEI1YPHwEmIHoolScDe6KOVmVwgybH+BiQXIS/GOVqDwrzEJc3xsMFI8S1otvr
4SdGpiLc9xRbEEHnDe+2xmfohkve+N0v5/XYYuHchPLzFgzjb8yjR7PLKg6XEY5C
Xhla/17lppeIeYauMjJciJch47eFOMpK7wmytaQBoLdZG73zGAPKETZvEP/xgOa0
7w/wRVYRjgSFr1SwpcRNNQV71IcWieqo7unxNjj/FKIAMoJ9cznulnpdRf/99ibJ
mjbIhysdFHl6a4BixMs7y16h4P8iXWM6RtJL2gn7UgCRFfBwWGTDCZs3xzhRZtOP
TwnwcYLNgu/QNhTOqqLKOYjCRDQey5Mp2mIBWF87L/d7zagWLKOb8VWAwbpLY3oU
dcri7eO+ooUHdRtY2gf09YOqMVsKGeUqioZ+XPPEtNqOR6G2x+czeISpvaKWG81z
fnqfNi+gcjA0xXZYY2EYNfP6YNbSx/Oz7jOD7B7RxKPho+TLS93lS2iU+j3Z2WOO
tSXmg9lhNeYciynbGoFNUQJRwqS+nSUNxcj5kKjT882zwnhXrwRSNSrPwt2v2Ygr
wB3TdS53ZKpyM6+qqS6a0YOXvj5bX/++ZX7wu9f8i64azAS2/dywmZoaJ+nZnixf
gBdKTdr/aYuaIyDk5oUwfXQHSdonVRjigi5dXloamNhowwP/ciXA0CPygnc1J+7m
jDQGKeGYN1oF1k6cqzz/NlWVbs8zsBhUX75ge7xJ7TIarQCdIVx+tUGR4n4hTYKg
C2AsSYmSvXWTRTuLMV9J4qCL12UHbdoRJzcQaLbiAG2HAwk+nYuskXnKywDxCRRg
XrBEx5UkG1Huo93uekf9FLibdICqJcWxpDc+M9h1ovRcxEqGminp9czPXbLLlKIi
49sG2NzDQATsSNXMpUEIGX37OtGXuohRiUqp2kRUC+IOOvl65Z41c09dqa5JddKh
UtVrh6Jua2NvVaWnM58aVg==
`pragma protect end_protected
