// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
blyjUmPVrliY4unGHnpxTXX2w6DIDXgO7j/v0VWIiIOY6sTqS5EvdvN4bH32+C+DPD+duDFzrW6E
pO9j8wRcCtvshjiZ72fI7ZqOhnu65q5/iTlWV/bqew5SB76J2+/VB4xZxIbEJZ1R6Oo2s8/cAUbe
GNFbDQoFwE+ZeRBTYjoQC7QMYmFHBJ94oGjMdANh9S5MFrHevid4LB3zrUHqw6dqTJHUZRL13NH1
nw6tXMTxN9PgDfMshkVC9cm8+x/sbvv1luaOUteJjiG81T0pVm6MBG001TBSo0A7pJBZ+JF7iHHf
eBgcrtc7d40SmOp3QbBBKaJ5caiRntKFnzBnew==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21056)
okw0py37IzReG8STnLwHy+BytRSnlobUyyn6Im4k2WWeDahxJQJ5yEroAcDthTqrFO2xlMhE+hXa
XviSSYekrvy0afmKaqe6b5mgmrPcxeCB4kRg1XyB7a5k//R9zj+cfThkWUXAVAxTDyH2bIkrgz+m
w/kA+UZn3rY2QnvK/HH5tm+LhV5wJEDkH2UspsTy6yY5DCA57jyq9/zgYkgYLvT7LJGRK+QWk2uz
OU4Q+c09M39DuxKvGoeqawFzF30ucpWy53/SopPxVvCuTDuHpM+deG71a6Mi0WpuFUF+HDwcWlwv
r43eeYozSXzRJR75JuixtigwhtPUqbuQXM+dbmfQzxe31Oyf7SKrTcKXUMormoYhlAXC0FSbEahO
mpl1Ekdb77hSC2M+wB0m1X3Jc0175w9CHWWNlfrX+6xGGnaxav+GS9C5uLYZMsYdL2la5wA0c0zl
UMAIaqEwBz+xb96IIx2J9+ccTXWIiW7pxhbI6x+3cInJm8azlkY+gX4+3xE7qlmOdQq0WIYr0oH4
aQZlrYpEY99skQ8uKbDpdtLbUcyVZVncfN/RmAqEf4wWvuycG+xRBpkcVE4PlJRYfFkrUygP8gpm
bm+iXv1IYaG2pM7QlYEX1Vh4NeugxncuvrPI0OsjAAhin7ru38VSHjZXu4aoXb28DBy2/Qcm4U7o
NSYR1LkW2VuBKIJDxjOoaMKxhXKQrbqSsccLiS+nBo8/VSv3/SK93i8kQZwSKwJhZ0tI2CeATALy
9eBPJQsRp3SuYgnzhaCm+/N3YGGuTAyjPfNjIijd4XiJPZ7ABVUlYYwJ2BHAlVhLyYfHAD/BOH+f
vDaV0QdqyNKvL7D/dVziB0xcy6hcKKnDTN15uFtH37SA6sr4okRzIohZ4zkvlOhXUCZsJFj5s2QO
0Sb+M2Ox7n74JX/5eNiYUZuAKtFlMyw7bSEJZKZr3L8R0HVbWZbs5qg4P0R+2OOyInL5+NTS0OXG
kR6+gTSmnDCKnRkFbdIWK7kTkyfuXGOwp7Hm1KYp+dcYG2jvFL3orQN1FfZPxERn3yvNlZbq1EBQ
dT0jk27VWEZl2FRahIka802pHR3qEBntcHoFOFMdNm63lHKXtc4BgzeQvr9MxG7UH5NPvphVWtU/
rnZi4H8L/uMxJ2w/lbiRMfUOkanAcKUAihsnA2ibKXVJUCRgJjyUTMxTDwXi5WiFo/i6FCDuhvAM
IgnyayFAwaotC0mW23yjHb52AcJi0hIfEL5jWBIzGrNOjKqMARrZ6ZSe0aGqvbBn2ZcWqxTgbRM2
gj33JHievyau0BqQR1jBhf9CzsCfajjM+G6A5AicnXt6lmywy9QSaEP9BE8oCdiV0oKoyhf2IkV2
ltdeBvdKkWw1aphlSM4LaLtVwDCeR69LD3W09faXe24+PUx5l9N2uKG4zkoYiEPjnxdZvzkH1615
IVeOCDgOE3qLXQDnJ5ovVC0cINTxQsoksuWIHmAQxaE68lbA6+igoYoXeuEvUnPIXg4hptwq40+Y
m//0hohbhZc+yvpnvv9pNk/IiLTH0sn9pyvmBu/aPMXUp2VckXnBM0uDZH3SdrOn0bnuTbpCfHaG
T0L4uX9Wj2peFAnXfX9bHwrZVOqrb3QXlrltbe9+k691BtdQEK6PNqcGcjDmkv1lnl96icFClE3G
xsT378a7aw6q56XFiPtTVNN+OijNhNwna59TK5P4vYe0mA6KqN/82gx2V/4uS2Sjkp3zUNiY/qiU
z97ACw8Ud1jlFQaCF/cdzd13UDR1M072TXEubSGoPPknq5xB9BGaDdin24p2CFo7bIG89ms/2ddw
3lwcNrbUyqyyN3ql3pVAyls0TT13sz2ut4nyYGNcMM1nxVoOsBg0TllLihLmTslUAYvmZ1S3Hmwo
izYwMOPj46HpdMHtzgmCiCxzkFkDve2r13Q0VQOKoEpNiDammrvRjnMBzba/MlQPmXOU0GdV9Dz4
QuX/HO6LGnz6+ycg8BV8plECH11V1wpGNZORmU/i+XnMQdWYhZ/KtntW7lsIjXgIFaNOkLZLHuA3
9fVfRclGApY8e+3Xu+1sUc8CUFwxRu6Web2lr25uBhvQk/R1otNXGBVeKHk9KFol/Y3LAkcJQ2kN
Nv7FjqqTL69T+N69frtv/UpsyAoUbJGE/CI7QK6OoqkmxRXeIlONUSaPgSnhECTCdqm08saPJhH3
JTN7MYlnavZ6MgYfoGcLmTpPhrjN5CCK2evwKWdukB65VvZYhIgKs8g0BWk8+NTr3uBYvOppAezL
GLqz2l3FD6goiU27yRgibxhRlM26st0BihX8EzYQshrLSEPOJZOFxQA0jiO9u68+/BcmTH0f1UXf
SwCZphTYvBemvrlPiCw3jYyFT73USExk5lR2h38EHgOKAmG+Z14Z1U/4WJ8Pgm1+4wgH2nRjH5Ea
1km0V8TFnni0BoMY/AgEtYrBsIUrAf+cIXoCh9F/tqAn4zHAcWN5XLB2nAYXyHRM/qDZxwEXdK9/
4f8gTFh/ZBwAl2+RTsSDHFUrQcxYqnEWq01OJcc6yJdVCR+dVtvBHWrTr/V1yhNIJm8Q1bUMvCEn
fU2L5KqP+E7lcw+ltCRd69rryB8ytTn7kIbsHou6nkEibai6DDCtEelUQdLSVtfHAWsxOsWv9vu9
c0uN8ontXFX9w2n8teq1hJs+eVdVTD16BPAIlPf38l5zP72pk2kR7rcmhmakrWyYHHQWOG3YY1/x
g8RWckB9xO9iM2WdpOAzFlpKvdIqGb+8k3RQQsQVtYB7kKnhKt7LY/nzrXl8HDzJiyZTocTlkhLi
ZdwlmRW8d2Xyq6bdx70WKaBIZ2Mq2pxpUM03O8qsMK79/APQYDhcm1LGn84CIrxd1KxRH3T4L9Id
9MslLX7RL4JjonBDI8ilAhvayI/rPJcotbYIoGPsHlReMbxLQTyF7DgRWZMBn47JpN+eqrw9RYDc
/t2ttN1+LtHy6SpkFtzQeKjTlaX3CTCCSo7/E1/I2lKbxo+A37AiJ/4Ts2cSk5Lpa7ThqOZzhyhv
PyEnl+Tvr9Y+oYLLx3myaA3r2ZpkliCuS450gnaDNahtf1cCuZbhsL6FwI6FhTzMlgnZYfuNMwyp
CJ3WYCFgFsCC867vg1go+JxXkDybOVKzDIv/ySsqrDZdIZevtXJ0Q7wNG8esN9pp/9a87qF4bPtt
rQVJNqT1JURBcMQFBsXWf4IMQmmkuE2eO74jFwfuUlIyj9Iq51TtRSfGsBJrPp506Eq4KBXiOBO6
R9xQxeeQRVLU3Ma6Rok+PrIrB6JyMfCciGLIGKC9Yn7pEHOCmHXeSZKVhVq68jk3lfHqghVw/t8O
mxzO5FGDIxKhb8cw6MX89vLissYV248xAn7/kAuOO+bnDWHbljpHLvbmtc7ZBnu9YN6mlPbqeUii
zb5uolm4pSf7gTbz1X//ZJtAvHU/Px6/chHBXNUGx4zjENd2SN8aOYvpDVDAe3LIWdTDATQdMTK4
Ps3/ugNU1PnnDMI1t7ACwpnR73ABN4MWg9hGSN/RLe3KcMnQhBXWsNCqz6KFv9I/MiDl56hD/hnX
7JkVHzsh55g2fcgNat5eXPizSP2TVGZf8kW+0FfRC83PjBiygBN5ZMioGx4asyGT/FnYD1cgmmAr
5kHZZU3E1z0iFSkMOOwu7kTFEH8lc1riyrvl0b8ObS08RvhzwdDPb9vVQrDFfaImf42jP6oCQcaT
bsRxFIT9VqXg0T1StE3nsXvotuJwj51dvxCKM3psjekPKCRQ+jTRlCvTBTWP6cF0S+E54etVefpS
2iF4bEJC9FW6SCbwapRCD0GZlaFBLt8fF8j/TBsfsFt7iasbLTOArjaNpXmhAfB+2/reWA20JyWp
TJNrKajC8X4iERWqfzhCmCezIvu53ZwPETnrxXTw9PBGUPbFk45/7i88HWsgEyDfAOhgpnelIH+w
KgOKZ1uUS/7dbCl9X2suTUITEXoVbOGjsaXXfcXxbYsST02YLJtaYAX+ljCEUlZfm+eB0XGgj8Iu
TJRI5PzBBeNDB7wvidmo98yf4pps0mq3WWSrBsCSDVNQuimwPx2ZbkeqzN/U8YelEfJ4kJGljil/
w2B7euwU1KDnxEIYj7B5HcVtMv0/BupI3+qc1kYouw5ua81M8tqDyHkFv1W1i20nyOPqFHoPjxcn
bbl0qOrL14c40XqcWTsCgFiCXJVog8AamN7cWieAXadEwPL/56U7vVxJegUwWvo6COMNJ5kqiuov
9NJi/wFFqk5zXXJKWmDXiu4PTpjbbluO5dLWmYD0Rrv59Ct0kbZWw7E8nr+QcHp2Q97/Mg43ly9e
BBz2ulhRURBOoMIbWuXvq01ob75cPBUxjBpQ8emOxL9iYeVbMhJxSkrtngA9Tc4JhM/WbjAZ87hS
xxjgqwozS+HAkfJYMan05o0i7FsQ5C6E7SW607c55yQvOw5dR7FRmiVgxb0fX1tdS/v0EJ2rk4C7
28ZjpjY2UlDM5v5W/4q51rxrRuirmcs9SySjdk6bNzUibQerzpJpKXdqzprhG7kVlukr0vP94N5j
ibI5KqI9fLTeqRvpMAoWrXX1kR0rcxZLsrIo5Vl2X59wPqNy9VIqFeq/ZgdBC8SXRc+5jesPG4eu
sqJH1KxpI1U8CeTeCp29cSs4sfsA5fcqgMBXBo7a7MHPZZvWtv3obiLrxOJzPFVNCs3FGlKPlGeM
oN1rrO23FkY32APh4NCr8YpGkggJkEniwrPpagLom5gIVnI++DSmO/iCbLZEAvl211AVZGa4hiiN
FCRsYFO56+O41MLG2bAZvuvZ+wCwJIFIjIwGoz+YGRpmxNDNf6Mu1p2j6otrkIuVXjXFHQDevF77
yaPTCq5rQONNnHgXIrvMGVy52lnla6DK0lWT5oujnyCyzWZytg537CBOS2THzzuze1+UwZvwtpHG
yevmUBTTTAAxGiRsFb/+pV3NAcSKC+zN5+RBaQvwmg44SC3rggL/Y/yoNANKhGWovNNJ0z4onrc9
owZe0Z+M1W/feY12Kzj5xao78/LV8nxOJybwEzeok5lB0Top9g0u9/Zz/9ym8eo3dZ+/Pfo74kOz
n2dHBz0kxl+ZgfVVF1+Qa5geqBYuGd2iHQlxbbmXHn5bjjrufUdzAb5mMgAzvVAESTP6GeDECn5+
Ti7EFRAGosspCzSdyeXjd3W7AUH0gjzYwsqeYiwoFR6D/dehA0wBsKAFqJC7/jpKdV+zzJ5j/2TQ
mKJoqFdNgA0lEtfo1y3T7405D5s1PG9nKUXlbOSRhqXU/LHwZHk9CtFwHgDoR34rW5xAe79Bikj3
ssQCg5lStQrWafAcFdvFZLtJe61ZJUXy+OQc4bWaVl4t+E+xlkbtrfSdOLz/utByy9Le9AK+3VZg
CQw6I9kp+bTNhbMeh5iUpBmYBCBWl0awR9+SjrogwCrBI932YIMPnG/oKROcEBwFnmgm29D5xBeM
DT0ArAUk5MZizMWvXj9B6vK9CgVmoCfVE0SpEFCM4LurQ802SHPnSLuE6jnX1Je7IBI7FaEpbcl/
R/9yHFnwaiO21qgszYXe9mwWED8SPDg/JmBupcZtjIwsFG1tNLGHeQLJcwRGe3IeIEJeTv9c2mqG
LPLOoLB90EjDvDpesKzd4IiiN51EGh6tyjyczNV+SAAmRQYPr3VvB5YHldeguey3TwPxyFfNYaZT
N50l4T6i463eQPtVcJkKWj3eaKI0VdLlY986Tcjc1t7EZ7gV0rbF0wGT8bgllpyGuBtvF0LmoP3k
u9QjLOhz/AA/wVisxtKCbTz7rm/Zx9RsOvc/0t6xE0JSVkvvIVx2xx+2THjhjPf1gIhDlt558pGn
J0ai5eLNJkOLNZHc7aCaib3r3BV82nMMljuf8ShrY5aKsTk3hxoz0NfB2dppGDuRNz0zlw3zizTS
ii5ZL4TTLDsDkWU02Dp70u/CE+IGEpEbVmxmqBvH1X7++GOQ7yErbVU0sWJMhwzXPR4vnS0k187q
1tS1nJGReJh/SWKQ5zFUjOe5QXsz4PPNUECIqHYF+0a1jpPc7815vT0F24N6Fu5eC2NfXuUD+EsK
SKVox+cG1/oM+T191e9MA/IPq4W5I1tlxdVvwJKnTRmZO52NIDW+dvHKnhmhHLR/Oc8AgoEGcBeV
qanf+mBvirqro9U3LFBDV+F6EknNQVKhOVQK8KKjMvr4+GIMKGLjeQwhJL39z9boaVOCZ5kPyb12
C9YbnZMMY4fo6ZF32CmNFkF9GHWwlrOr/Yihu9ANqEsL8dFgCSg3h8j45EhxyOOIpOYGp43Z999Q
Cl4K0mbn4VsTPaQELffVmMQvf4acaU32YmWwLbbrk2P5yXOjnrh+QWR4YKUCi9Q7P3B0Y8KCn+05
2Nas071H71blaNyHLVzLPX+SKPYSvzoPtsYDbCBXnE59Pdo7WoWtV1AjqFmIava/FmHtrxxoUELe
9YvQEy3Vnpv4bLnlNZyqiOqbQXoKg7e803di3BxPabClMWbWNdxJNR++nnnbvY34325JHM0/HByG
qXyjKW3CZC+UpfnX97HLdpXDB5R6CtOjPcL5as6A+k17P4ZWGS9iinjhzkx5pcpY3jEVc4NM9OlV
qHCaAj33Ta+GmCyhwHFkpQSGSUX00DCl3rf7PhQNSHgH4/O82Ov2TNGXPF3KGbXK30mLJYVjC6I6
bIUBRJmz2WJggsBsX2bGLvHEhYQ6+VZQE/e9rXIcFu30s4oWcq3NcxeCFCNfUxuaXYi6UsY7cbIG
HS07DTVENVKF86KWwJvcNV92ydp7/O2GIil5otIVlCB3qhbvtmgVc2/I6oMki/cFsVL6L3+op+a5
iwh96F6I+BvokXX3G+/yj60pbDnpZpa5e08EHxMTAxyxCfPIVyPZs90+O99Qr4UgDxpow2Fn1wxP
lReo2+xUhPoM5wb0vn/uWHXEHAKUpzjKvWXwLCped3EYqAma0yan/24C777E0wUr/4V2leDs3T9d
C0Z/0j6/0AkjFMoEmObBW1Keo0jmmMSTxD+ynRr7iIfBl5GYwn3QJ7i0GaC1hM2heVcc0nzbZ+BR
VaPpGxKDZ7RvvIFDg7GrPpDCaDI5ACpkQqddZTT+HRDMfnwb0dk6oIK6P8g0cWLTDoZ50pjkBS1m
fSuW2zgVeBI+KCrliuMzz4ackt4s+C5lxjDp8kXAHQxG290TLTc19wQlXXP7dJ3qNs8wdQBtTuWL
a1SIVjBloMYayAuBvMhkN4twdaCKLDIA2TpI/mRjDAvQSefSEyealyz2f/cz5nTAuetL74+lu4Gn
oMrFIK3RQoG/YhAJBa9MoDLgK7zgER8cHJfs0QAalOpu1BCVlRwaPuNP6O+7QKeJ1jzSVX4jL+Oh
84QRvk3X+O7zORyOMJOFqG9lpguRAQ785Fu8y2JYmMZfXtphYhPuwn+yq1HIo5SX3SvTNr7yifSz
0J5G2A/2bRn9WQFzDwiDXAe2GcH927W8VlzpyODJC9y3mnFXF/cy7Hv/PWCTBaLwUoMXXi7tIohT
0vJ0tPJbh7gQ+eYVPqdDXyz5X59atvgBaxld1y7xAjDcNVWFT9Uav2FDzxOIoL2OpIXV/mKYvH+g
HLxfO0BGH5HuE+smmIZrHfZUsJT7bbC+XrgeB5ARE3Zol+rH/zi0P0/2bm171hZVEesx6J1tRm46
7U3U/NwulmvG+PVVH73e4RaF+P7vAWqecm2JVFE6PElk3bXZAwAxjy3flwuyEBiYtlwZa7sRh9oH
jp33uRCVO94wr+vrjmQgZm5zaH/Kj/F/sg4gX/BMJ8uIwki/k4wsE9iYmSdtANNmN8XISIk4GAs2
j6IZFSQWjcTeT4VF+f4nBmlDGsUtL5097cHBLSr0kGindmauziumM/WWKRpYv2ZOC4P2xO7KSr7o
ThE4am7kN6MdkcMW0bu+2CHZ8TcsGFAPxv/rw0rMWn4dc5UQqVbU/QM1VkGedOsBX33/Dbx4mz0Q
vSN1A02WQYhGYP8tvmzUR89aOchzfeHCCy+MeMGQF0HqDYQdpNVSCE/GMY5mYTcggeKxaD2Tpf0Q
6gHgRCI1GN9oVON75H/HJ69mB4mpp4lbaDiAD8QFm87Zz3UppPH7BsX5c8pG/LqK1DQc2kTax3A9
cNqEcN3ZJGdMusypinBIUe1/j6SPDjvObScwi2ISQcWOIjR0IQeYazxcXit8dwyVmONZB2ZFeYUX
cRTAAokQD3Ml7KixomqoVlQ9OUiXVJJ7O5t8X2zn+TDs//lH2V7Ing645CSw+Wv6Hgxll/sj+y6S
AxhsXJ9p8KlCrWzACgIa/77LdU1PoEN4M3ToW5v37HOtaNLgOzMs6SlyJk8xs2TPSxqROt+sIw8T
oeAI2K2f58yOskM0NxZnO6C8m0drA3P+DyE+BmnS6YjhVtoSRhJZ/Bvx1UN5PTEUg8vblzS4vRnr
pNTzj3QpZ/N6v0oWng8CXmFeTw3Q7WupUtZAaJNfJJ9yNdqFASEYi5LGfINXxMB2UeFoDeQuWsSh
IkRyl6EsVMfARwj8ZDt1znjexcZYWTK0NhECDx5nerBY+5tXggWSKGujIKPr/yd6FyMmKYA72poE
WCzFv6JO17am51nMa45SuZsF55T77pZojY32Xlo02kRRLd4oWUBWc34nUKdWuq2w81XSSM/hiU7x
lziMHUN6DkmwJ2e+1nj5pR4vls3i0/Th5TumX/Ih+w3NYITqnyGAizBPh5U8r5aKzfsnHuXhjvIt
US/6HthAVdKPYfblJ8FJUOLVL62dTkK6vKVzi6FMVGUVJL36PDwPBtcbU7MVYay561RMBZkg0+ts
mmS9pq7Goxm3LFo0Flaylvl7YtyDta6/O45pZ8P8tVGMqJ+Yq7EK/F1B2SLHhZuj+r5h4GgZmAyG
6ScV788VDfxvmia5t6DotADRbkNeI+osNcWX6DX66zaunj3KdwB+rx+xras/62/6pwKCnsRl+YzZ
b7ww1am33IMGqoWttMzHjVu4qcNYy0tyeSO1RktQtD9ieZG8YX0OOS/W8OLJJGpJXH3fKetWS2EQ
PSBlaIo1PrA30L673dff4rzCBsTUK8vf5DiJsZ8/rhN+a2oChWU7YwJiqqdgJrph0R9ErJZAdwoH
ifZuXcT2XyjJ4OpSg+XIY5+gUM6FpWyP0jZPSOkHN7O+P3w62QynvG+4yDc35pUIY7dNRLjRq4dU
hAFn7Oym9o9RggSngyzLHCJXncjfXv/TMFuFAr6VN2QrWPzJ8P8ldgX/mp5oum4G6Bg/nLT5oeJk
VVSWcCAwcy07007E9NUGNN1KZxOcLLIsS059ncT+pRfs26t16Hu0Erb0E5H6UYPcgadl+FKNS2np
9P36IGEqhfY0HXfNbkT61jJR0LTU5Z2tKtdgPV4bG5UsZIpLl79BSfNtwT2YQrZnbL5EJWrZqfuL
LTWflVCuKUHe89QAgwGxnOJEs/yT9amVK3Qpv3JhtT1gsO07EYq/E80T09t8WYJLsK5MX+SKTkt2
eNwhede9jRGyEnC8+xQGbYKVkGvVtDzUjNUr9Shu0GViFhA1WWb1lBHcaGbTibin+6gEc+M14e4j
XXHYy3U2lP0X3Z/eD61S4HOogJsNqj1pjKaVWCw5iDxoXcfOa0VK2wWfcg9da9mtmmlqEGsrhEZc
UswP1TO44oTJ3iwZos5+A03QRfKEKIX+s08rCSV7/Mtd28tfo/riuNHRb0/8iWcS4amV2KQ/G3GL
B3YJZ9OxzIRNCY9DAXu0y0Gk6eVmwAUBGxW/qFon4NdPeBTzsbBj33Wey5gh/HAqHs8akT3gBcsO
JBNpad4w+6jmVKbbqRsgkktpw9YYsx0SqYExLYGaMRTSQcWTpn12hVFUvwKpacAmoLqoW7tvhfRm
LWm6CZLpxqyKdVwI+6vivB7UDSt9WP3zVk9Rpsn6o7UhxhQCQGt8pJPMHH9x71anq+kHXOLf2slN
nkVF2fHs1Q4AFujotUJGv20xH/5TnlmlOqPfZ1NzcY4Xao4KI2NCiFnUzXatOO/suI8nb7O7uHNK
eSDH/SFGKWoYVGsqsfy/Inl5BOy5/6dlAVc4f/1q2AoQyVcIZUZCeuVA/OPJkRwefHX70zv5Kcpx
7Ug6g456KWrrJGagGq3KZCKJq88kGHeoZ5jtUSxEvZw290w8sJ6tlkq36rN3U+wqcrKCLaFKPBJA
uptZX2svv+3j7Pc/0le52USQPcJGDlSjrkGS5nCCFV7wxAT1XuYttWVyqZeqhVPoVTVrx29Wt1Ts
WFvP2CxmY86ggiXgrrKh0hrhooUAVjDbZl7dvgfcvsOxSVAZBVOrDA/dQf1KMMtHBjuQw4eslZV9
Rn+WyM9NzQ0DrYTMQZ1oTWQ+WawBGRpi2Lw/nwbFQJWcsOg9WTJf8NttrahtZlJW2aAubseQLfIB
9iSLMzENvI65fibM/6xqjQkBkq9q6iEtz2DJq/cEf7c/8xtRp72hgLVWR8dYqb/f1TQWaSFKpAZE
uzUVqNItN4uTgJYS2BBsXrhFlFwQDdsChjtJTxZ7Xlbd6fZUlyxoWxSkbcrkS3Twnnk0tvoTNaLX
hahpAjMu797wdnkwiMYtOXSS3/hx49nhS1HgKj5t2hgAs4OrQtQahi7Z7FcXJdSwLRWh3go7yJFY
SbLHvNMmxob5jftoxvmNGbqKGaquEdMdHP+hwbT/Txpt5tDHlqCHuTfQXe/Gd9EJWvmzna0eryJv
DEvwaRrtEf1n2TK1G5yX+CtsLHGi796nE5LFNxwAAlTfI5KUGd4CIwK12JMJ/Hnmzo9uCLO4E2vX
gtume7YGEpsSEoSl4ztmExTfPy7VFFzkmQAw0BjBi8ak+X+TT2P7ULzCBClA+O2vZ6JohO3d3BEs
7AFbzJK7EK/tedYOFKm9uxjfpW969zNmvrFSzih/nwIzadywyAv+MMe5Ij9wqccB0iAvyyCPymdX
MYkgPeYhBUvkWpc4u4Y0NmKWXV8sraUHn+5AOPmS9cz0jqf91ZVThJY6bopQTqErxQQT6pmj1Oj3
V7gOI8bnE9DqrFRcQZSH4KIU4pwWN5e0edwyTpWMO4SGTH7BjimGDuybrSnXkzuPmH4WwSMj56rc
3S3HnB4zVnQUIuYF6C0/rtTZ1khumJ0EqtsPH+3rG3OlmDCs17Mgt/BJvFlPaxzEePzXH2FwCSwR
cW+FD0JJkts9ROBBYV4XQXNjVygexWHnd0H5rzxlM4vercahhTox8YPXiC8MAt9dFImKoxY6GvdK
Dv3q8nuUPMkpIc8a8zg44icSjPTXcKcwFNDjMkIbP3NizTvHYt5CIqU7RAEuNNQUunvNEwNJyQ3q
qjyWCn0EkP+ujKbEDmXUVJt5Z9ak3SAhuoCOHbq+nOKPSQEKAvmuC3EWKqxDMZfrOpFzw/vODG6O
Q4NqRGH/k7wNzVuLmOG8sIYsFgyLiM2UubpplvAttn3FqhxTSyR3ma9/NWpWrQkq0iYEfC7PvgrE
w5WFMk3p/zflagy6lVIhrSJ0ruH7yXYtH38Q9DzeCP9UUWQsZqx8GBF23dfTbthLBxchv2BtwJRz
+CbTXhuzRs5sBKlZVAIsDPE64gFVPfoxU1qbf8NRJIju8I5/AFqpz9ci32tsqBXMpfamY+MWMPZA
FKX3R3HR/GUBv/7SPFmn19CH6IiA7aid5HmZNsmxwt2YBPGutMvpKiM+HCR7XMeq3tCMyeTIbOvO
I423QRjzQVC5O5GdiwrMNdMa5HmTJgbdOIbDNE6FHxE3pzS7NNN9BTfhWHCRdy+XP+B5teD+jaIa
165/eRatNS5zUlT6ROqFVB3ZD9aqOWRHNC9bmwP7GYAcuqWybBQ18qbpe4igw8Xle3GQJXgZHmXJ
9VpAomQ7WjWUcoYZTxtsSP0C77+aJO/NxBgE2Y2ertOwp/aOXws67bDk4H66jhUDio2TGKK5CPlj
/Zk5mGs8aAfeey4rt963kS20fXy2W95KUhpjZ2J0+7pU+G5q+AwunUcVqrXd44bKHioeUOkXwZZ3
TLoVlu3zeUlOPnS9zMsL/9JXzGh7blaw2/n8WY29keWbgnQ+hhGtJqw/8HRs+Gyp6pGzHt/yPLWn
i9B6nNnHRKtxqWLNe3l3sS2lWtUFYkfs+icNANLWPLvX4QRwY8NQCQy64lbbLzwQYKz1eo4Afz6H
8E40Kw6da/g8apwkRng1LZwdGr75xLiWeCerYmckDtMpOm9TzwXqqJsZjDWLMOMxNe6jYNjUb3vy
wCL/fRZNp7CIl0cq7zd512V3Yx0E2gO0ZFICORbWqO1ao6+P9OqVAKKQRQ/V5ozCwh+q9V/3S4oe
pGxUlO8IwLBHEnRFYXwiiqlxaLET+m9KcO602Ji7I6kH99MW7A7GRGh0qP7nDT6xL9lnsCuvmlcm
f+5ip+qzVnuYSAzeIuctEqGZqi9ynP04r7PskK/t5BeDrWgqm8IaSibTotpi7vXOo7PrPPzSgRTc
xecV9NFvA38gBdByspMsXNQokW1viOtmQ9Ljc0D4lMo5umgdMz3TDdyf9AnE9tjPrcKHWmSRgHvF
JUbfXgSt7VmtfsgIZC/MW1NU2E2/FLwabV2uI2n282IzJunv3+klnCc+pQD0RKt20ynCSbpceVOz
0ZylvDFGzl/kM2/65VwH0sZlRg/hH7CycOB9CTb9KWMNatV2TcikskcXxcUQ+46/hPiyuIL4XzzM
E30kQ3JHTUawlws4pP2KitoiYO1y0m9uwZFQbHtSOVuFFWuTXlJZVnkk8c2BjsuoazZzstsu37YD
lWEQx+Eaz4dKWl3IIKYIw2UKLYPd6Gi7qX7umwl/gnv2LOo/7I0nlNnY9yXOwWQTZGmFRxGQM7AH
5rgrFOIQOyYvqnQ8o1JZdM6wi7BP1L2tEoM9NAHlTvP+qdRWpPBoDNoP8l4DpSAQL9VFfSAB8BpP
RK0goMZBs4eT6MSNE0vS1e5eLrvhKiSTStqgSHGkRe2rV13lSYlQ7flnZnenJFwjlgGiqw/TAcpp
SVTRJ4dVVQPNXztR+vx9iLOfmq6jlQp4GOsi6X6+iosti/pOPeFrgnw+kZPoMhqOpzlqolz3fgqz
Iy6rZ6ueNkVMPFsk7ChwcKwseoLR2bx5tNxc8bDOGSTE+zXZL7mswiOGXM7eCFrSLhuMTYA9Q/Gl
ozfkxiuYKwweiO5ke/T+S9h9FQPZa28tSu59/8fynGOz1cqxNiitaKrm9Qp1gVxBAG3OZE0j7APH
U6vQdHjbUUA1DFLdpDPycc2wWPJJpefj/fbej9e//Qxb7ZqQAZuih5v6eJIqfdvyjckMzU0nUNo7
M040qHd5eNJ/2PtDxwoQvvCsJ2bxH+M9fBT9RooltE6rBploYuzPuBQ39Q77b4S97PsJrNlUg6Sd
8ZVjCZS2NDP8Ku5+fzpF25In3dTeRL26P2P+MhKZ01XAlJwbZyRM5GfEBmLu4zp0Df3QMcBHzxlL
iqGJcdSjFJ3PPg1gqcd5XnxUQMbSyB9nkGoT8oIyOTIQW+fGvFxcK1lR8iA+CDI8nZmsO4z1roBw
MmyPipuMK2YUQYbuzA4I1eXN5GTfTM5D9nc9+tBMy0plvlWCstpSP5rhIJhnceY9HsjDAf7Jq+hZ
OtnXjel92/oDwU/gnJVNqIrfBoWUBmhQpu8TRtllwu+WaRFp/Atxj2LmPjIN9whvpXRfwpaYqQh6
wFztCKF7ZnOX3pBESkbO2CRCYpoRWN3+YfuY23RdT/yQBsIAzcPNZXrhoiZuyvCKd37c5c5eu5+i
09UoBVzcAiCQdOj4+9W2RADR3s+bPGKPH2Pj41iYTtay6LK46rF4cf7/wx6B6yTfLhVGP7Xs4Qdh
K/qT7BQjZxX1mJBQwAYa1atc7FPs4JufH6ABnSrNfGN7p5bk1Hi6oPVOUbSLnQ6SciUJsvoe1Oz+
jr3C1TONIwtgx6wdavIHlC2iMqtIBcsp38PKSaCd6Yy6ywMAei4fPcCYLJXsAd1FFcBYB41bs7mA
yMAaXCXPNdFshzHg0Vfw7ZZUGtId+vKiyihQMNaNu9N8P2RHNG3PDNaiFTW1U4gL2+ycVfaInKH7
FTSLZYioct63CWsacutgBJnf/zUOgVxjyVX7UmxflbtkXPfigu/fi8hGGRhNfr3tKVWsyQAawUvN
MQ6TenH0QzY9aGPVYzhA0xaAqIYritNjV0t/dqJg5PyTYssASwvzejC1nIVo/NlQeHqqCbfYiyie
qfdeKlhRm2Rql7/vAaoSgtRqEVz7TZjt9PYgVp+8CvFonoWKcBYA0DBHcDHog5tQSLMgKQd9JbGf
3+TFgYzSZ7srjEV0tmgsDJVIn53wQjU7GXCBo+vbhg+wyKqV1IG+Qy0qV7hTNNPLNIXfo78mcL0F
fuAMhPIzv5a6iBbX8WTu9j5/ClIdZmcbNi7Tr3YyixXRVlbadlkHj+5pKNUBw0wehK5co5QpJ7qa
8ZF1AU7ZdUWSqqTJJ6YBhumJYIGOI3+QgplPav8wpWsu6RqKExpWdz4xcLysey8/jpXa0rRyE91b
8A3tnaJ++MQVD0gky49XBZXhH0nJPFzdSiG/Uo83RRVg6t72YSyvPqJ3SQwfAwPofgLgKf08cSBI
lD72ORb+VyihlkMgh8rF+gmjAhu+UPU02bLaYr1sDBNKM6LCFmHMP0BI3GtIJZOSNoiVKcir1bYa
Q9qDAnf4izApIg5ZNjNHy8HdWpC8LE6qAI0n1ZW7Lm/TjYUCEJs+3LUHJDamrwEzX6BULtD1RNG9
bELxXvLteEMO1tGP9Yz1062wsZSrRxnJ7EVx1DwJPgAOqxWfk7ALgSoTTrknJi6/0gYYqSgRhrO1
9J3gxmCofNsRP+wQTRjfKjIVe8a40teJAltoXDAV75VuvN2JOonlc0vlFEQuIbofr29U7YqVvB36
gMn5qlRXqszvGTWLK7R4L/lxJHyZ/AqLJg0wfYFTqEAX0iJlBrCJAURSGgMDau+/vk9CStIMJuDS
EBD/nV7D4x2amd4zuX5S03fAmUrLHK5WM4mAnN708RQQRhNRoKgDvOdtKib/imxz6spKc+BuluLl
TXiQIX5SsXU28wkY+dJf3RvwoMdBUnxaIJ2OitGmeJBc8Vyb7B+uUBPS/UfuE4A1G3CsV/w2LHCy
oXVU7WSMpVZVSYaCuQ9Pe5+YsmbXIm5mkA6rqIN6hAoCXa0NaA0opC4xLBtPZ34f1EQv5EqCqmMX
aYxdb7Tz9A24PSP+JwyyrQn06p12O5Zo5JBJBBSQ7R5vbjar3Gb2TjU4bWCTvkZhI8f/RGDDDpGr
l47UHF0gPbqwrivq96Q+0LU7RMCMoUWB6BOp58VjxA3N76fXzec98zvKRbvEdzBIkd2QIw1uM3lI
tnp10mwWNdKF0wBsKIo9RYhsgVG8ZjbYJ+IBrWdvgfHMqnPu+aY7TsDJWJW6f0NQ+LW76ViqC69B
MzgSsJ0doYwuRV2Lbl5qp1Ww5Y60x5CJdLGapzrHhrunOaTNblA4JagCxlQvnT04yTZS2f2RyeS/
iBnZCHOjOj9sSNMqutIz93Rpbz/a80FDkNE5nPQuIfPFDl/ppChdGF6eogWTg+OzLwSZBvNkIIri
MOD4h6QqmN/itbVqYcxqW6XAnAFiAnkzZIge4G3yIDj9WsYR4eoSqV4WXve4FhiA7Avg3ep0iAKU
C1ycckQG2m5VIaBbbrPRzIPKUUGnEwNpQVMhUrLNjIZrPkKRfkooJLJEvKA4axQ2iCfKrL4NRYEE
Nrpy3FnY4Yf5TbRCAXhGCDF802AlqLN41M+udwdWVW6oTotPMK/v3mjk+J34RYbLIexJkvGgwplQ
bGsGtutg9Xe9rgVjzF4ZtQAeblEtGcgW2Tl2RmxItpmOzWgRn2jyUC4+evZQqXa0OVmQxW3lI/rG
srCY8GThqU8ZSsc9BKhMEO4vZGwC7xD2P/yg9BrM1IbzGrw+FxSSWSAsTrqzkDsJOtDobZDU3HgZ
YbqiOGU7quulfHbPHSqjGgOhDbbpKUw88Y0m92OcnI+/U+Y+BMNAzzs8KalATNXgEDL9jRcnYUaL
F+We41X8hoo90l7F7yicYzE04XsPUXASF2HGkQxTpAUMXckgZlCfvUzvmSfbghfoJHbszzYXWi7X
CNHq2xNylck65K0NSK31thbiooanA2A6IMPF9ipMSBp4EQMw6QCOBER2FUBW/63bggiNdpUGqvGQ
1ZkYiAzEsxfCe1Gu4lddmnTd1b/ZXWWa8oYf/pim0/zlqhTZk9g0hffP3yramQr3PpcUPW4L/Yp4
Dpoac7fi3oH4WDd7KtDpSbV8WpUrdiSzOSfAlL8AjmhSSPYCaH+Ac2rlnugxzgl7M5304e6ZGRJG
Ebc/q2ODFXJC88FaDB6S6qZVKL1Z4mxGqbUHeEH9S3mVllH8c41zSf8pVB11cUcRVLYf3zCoJ8YV
yt8cN+2dlhwg4BgEdmxFANSAIDHTlyn2Ni6gn6PlHV1u81pIejLcNdVxIZCPWwuVs48NzwOQ5xDB
M257eS8LUAf9dB50E+BQKA7wKV771x1gRncZspXaaTw6oCAs63xhNtrnpjGJEZ0pEWrYvJ1hzkNc
N2WkQP5wId7mThN7oYncULYZJVlmH6MlXMxFsRA+NBAStHBjOXo64IBFmNj+N5wMZYCraZRVcYQl
MIZ6I2Bgs3H1Ha/4PQkNY/RCRZIGxaMGlNoCs20e9S1FnsCCgYE7RIxkehVdGrpRlUu7jySdQOxK
/Bt3aNzPEltenrdZjN3kQy9l7KYLBooeL8bT7SjYSdUrmyCQ/oaP627OtIhfe0TYt4Ohl2k2nlvl
0qjY8gzcHPs+vrDBngb9to4UTNRbPgUDe0u9xVrjqjkUXzuwdw7KFkJCcXupB8uw6AGti89rya8A
ZlRJW0iB5ariywfo9vpA8wRdfcTBSydS8O596hMl2raavV4zKX8i6DuwflEo+xeNGl0Vq7xs8rt9
zqHJpG8vwRO68R/BV3BQ9uaht86gWZzYGdvK76SzGrUwMKvSnDeSYf1PGHOHVcRNznINGG83pseo
/hbfhtOX2VEkVMlrHLrR5gCp7cTpV+HqcEoKe8YNOBhpwv9YjDUNogp5Cbbsd5WyvrASgP2zNFvx
BBkUy+Oug473TC5QWZvcUeiGsYilAFGFPVUjp8Pf6vne7losmYx/LvUhVXvRmBS7GyzrBjupC536
29XyniUQhOI4Kg3ixNgHrlGnFfMGeeYP8mhwf5f8LatX6KskX0kJ0u+5qXx+8fnwAkfdLeAaWvto
wSVjjnA4XrIBwBExo9zt9ShZ3oJyhoQA0lu1TUNTCGsEbmbid26x81dMegQNS9ys2o6GHAu9YWw2
vxqit7E1R4+lqDnBshtEBjaG90zuznQ9r6zs0oG+w6mAU3P9az/sKAFaY3NT9OQAFdXDKPcgFz7p
SJzbuSpk2jLuyf3BsdlHBAc3xgITtE0poY5ULudkspSrYnfGIFfnW2emqiV01QU4roedwfB1AfRb
NKwGcKcuMfxSgstC4dMR+SiN3qzgI2Rcn7vwCja3/cyuzAqFtccnHGJCpbZpWwU60E0r7sKq4aT/
FRxpzXhUs/pB+muMcAumLSmovXedPcAc0SEJp+mqF/wDhiHlumzmvgLkT1jOuNn8JqOyLM/t9ock
Sz7j3EXJ50tsmN/NxF/eUX+27ihEHgq572oJxelE+RtoX14zsVlrHTm5tzZmWNyB7wJdv8Z3dTgp
3QhOnc6+V82pFALsDaPmehzQGrvZFvsb/VchDBLLqC1HNkVNLg7DVMzOSuBycU/MQLhv9PzHwU4l
pI2VgGnOPCfjPrWTuaAAVh/nyQZMmj0Imq+l7JsPfw+UcFfYVGUpYXgvOT3QtsEHawllSqB/+T+q
vtlXfdhgLlT5DBsv0f2drL7HcufeNUXn5M3XyUSUA3TdBKa935CFtBu2adkEnP8YIJYIiKc2LmwQ
TLHts8HHXVsNX1MCmc4pArbam0MN/UrDwTvb36LdsPcSqtAMwAWSHyHSM46j9NbdRumv1fIFfyR5
E7u12v4OXCk8P2/+DLLtnIfiZCbdno1k/DswXeLs3oqxDgQU/1qsrsj8yX5j3cmRhfFiBAOZ4b2X
RtpzxzurjWhmSiKI6hwwVOh7/kauQg2TfSLYCxg1QrTIf1tAVW1B3dSs0aix+QpA7NdyowI4jNTT
UMWUSbCKub5k7qK8UVD8kTB49tFY8iSWGqZyPDmekM1Bm7XSiarhcNq+Ii2f8U89CjGWfSEUk5Fc
7MkTvamBb/YebCnZSXn9R26Lq2GWBTSzdUSXC9Ry+P11GYPqP2op+BPP8ax6hzJz1hmo8RTFoUlP
PNtUGjirhTqvrFMZ2L4WW0u+SmrQoJpt2l9KXQQP30VWev5rF6w7FyIaMFW5tpyJZlUQze7tC9EM
UNibGzlv5lSt5m6vvXe9OPs+7wSpFgGCKRO2qV4OM+vMC7hMS6tAuWgvFFBQRLKWm8n/eOYe6Q8H
Ma16xGqZCNPTreJFVziWrqr4b/2VskCBPdJQWn5jJokSJpX6BxNO7WHtP02P4MWenVKfjUJghcAe
M/oUZw651kHkVGvOdwWDVODbw+rok5snyIv1G9UKZ7Rqt0akT7q6h+TEUTIZDeb/DgxjkQi2lhU2
jVvE9+xk1KsElv5YMbeiUKJlAwLYrbvcw1g/rPLGLSr2XIlM/Ty7YbbfXgGm0HUDtD2JJ1a3SbS5
GjklGBRsh+RrektX9Tvx5s/72cjJiqitn9GcDCjIR7SUzXW+SgzubAgpEGxH2XTAXv3IDhGjAr4/
qlxi/vwO/2ydgWTkde46HUQHJY2rzQ8dy090ll6blWfAGbdiMmi4NrzIew8Hzwyq+zRYCQRHRbrV
9WJqBi8KdIgcifdoxlgpMiFCfqHED1cK9BA4Y2oCmpd8RJlgsSYcWhicamKex8K/GCPW+tVqzxy8
u3yzd8i4i79OSHoFb2fvAcw6RLDCjhqb14f7SZ4LDDVCoe8yWpgVR4VrDtpR9t/B05FIGd2HfAHh
u/6hTF7qj0iQfkjdx4vo4DTkrcPegHar/DmUvkmE/JpjGpUgmkg0yWc+L0s3IidpQaYhqodS27+X
PP5stCzGEVU5wNE66mB3MOMQOG0tneGWgWEBfBFTrCCHjiqZUttaUjYK9yHEj2i7A3pmW8IteFxU
jjG5l0qwCNB9UQxj9BM81f7wk1RWCl2lAaaLHKpQw7g8weN3pb024IdEhYwL6R50copRv8STv85p
PE2KHMZBoHqwJczfp098VMZrkWnXYzJfQVGXwefGk/UyMuccfdY/OYt5YGuu04ohc6h15t5/aqsN
pNlGllHSrL1JMQEoCrSuvapRyrkq5tlNSlm3zL/dVkXGEDGcXHy3rI8yURyYf87VfJ1LgfKi9iJw
gAbEh6CcaDwS9u+RYhp1ECps9ky08hNgv0v7qhRzzttg1khi+zM+k1bm2OvKjOqFLlLZaHB831Z0
YLFZM6+5/KQoQkU5pXqnzrAWwnEQwhFuf0aBESpMCK1+Vu7d3FK+MGuHOr1d7TB5Yqr2uF2K/Tes
tGPyMA+c5qWpXXQVGAhVgv+7OQkjnXotxpzAnI1SP2x1TdF3taTbCuD6qNOv5ZqNMe/gRdFXCkN/
RMCtclDPFYpM3DQlzWB25tgZjZJzmMT+QzyL7egt2g/d4YwFj/7BX+xaNdvn1hG2aFfJSQt5cPVJ
/FLmNeq9Z6m5mqroJDtxX/JFUKWppdRPr+v6MnlAJ0Yx+ya6UPSsK7b1vDGE41h1dCoaJGCHqFg0
o8KIH5gyrlAVrd5gK0Bnyik69XqKtRR0Y/snBog9blMnip9AUr0Opab7HDQ8qlDXobjCSp8Z4LU5
Q3CmepYyX7n2LjL3c6GBNYFSIb4brgp8wCR121TjUo8IgVRN5DyxVfvpV6QEoLb+Y88PMruxvCbR
2Wr5e15vOJ9OJwJIvZMtD0kcUNCl4XwqcZZdWNOwmm9pLBHYRvjFG/2jCUrkCRSSEJ3SW2ljTxpu
5Fac+jPmqfRbUHCGuHmW9s5sQiwD3rVrlCZqvz+5naXwepQnrymdIsAqG+lbeA7iWi99gZDf1idI
WzOnULQe7992OqEBtHzWd4e/yyV53Dc0MbZNouMqk3FdksIXEfZT51paE81MGyNgSw00p4j1p8qU
U9qir8CNILzkO9KNQyz7nQGgaBAYWx+zuYHJqhrUdIMYkZrerDLQMMHZwWY9bXXCsgGke5SSMUwQ
QIHfiMeNk2TRgccYBuvT9zVcQshz55hXMhrXnRNRM7Q3LuuakZwjR49MkSIS9rdfrWN6om7qvTot
G4I5uAebmBBTsQTuYYtFwduCZNhmxQ1py9P8jMTYdk1q7kMSlXBdauExmKkhofB1HfZpZ2vlIWzU
3vm0orxDMxK2L6kks1Z9qr05q3bPmBBfVZ06df3Qy8V1YVM1IpHfn7ZpicZukaq1pFZ7tpVjTq7t
j7E5cXmF9poNz4arp2gK+b2DQCAIZSuwylHAgJhMQCTtXHXRyCSjbcsJXYwzYtoUpMBIq8rxIqMI
QDWdPnB+ofmLJGduuQ5GOznL+0+Qpz9f7EPiLrsIDat5Sr1ozH8gFsHhv0XtDXOi/sJHkoP1Ul2J
4dmsUSlg+LPB4RLNx2eZvbgsfyrvQblPIhg/I55Nm8oNliQU/Sm2P4Nw9sXLiB1yswE8zaIFO+wI
qWc4Oy3Kt0Znd2bLLiWgHbCQwk369jRf4mbnyHRQRRBfWTDBd0rFV0rl/pzbOCXme3QfUXI8wM2B
Xz6GigGoIShifQmhqjhl1KtBy1EQ7leFH0/8vNWnciRilrvz+OXuz83Qo2Rshv+qE+1z98nXAm8c
LaR/Udx+lI+UhlRCf3znj4hmVhGvtxWSdH1R2Aiu6fUMyyFA7RQ/O5tT0Qn87rWcTYJW/4lDzYQi
15xp/mtRHAweMVfeBRp9NajWINgkIcNPsJmMP3+suZpHEvCdM3OJ3gp290OKxRUW8qa0Bk00ZtEQ
yIJHS+cz40MkIsM0EH24p7wAANm30RMq59Hrfo4BotxMkx6t0RrTtkPvpW9EyvphQggCeYDReK+X
BF55PrJZjHW+kC2OrQ5enecqjblYoEAR4xunLoHF0hgE1Tr+huY1FQ/Wobxax/zAlr/d5oycZ1sT
F0cSmhkYiRFcNcgD9XdOT747/LM5LjxklJA1ELOBcQiiPpUasFV9H6fMUMzh3eTcnUzfE4ds/9kY
DhUtwuzXxF9wssy/LqworHPtjdCGvxjuMN1gncHs2yN26ECYBDOyUij18EZun0vNMTKlmqqs4NmO
7wcahuO0DG9eJgmet+tM/rfBJ8f7Ya/t8b7gdQzzx4/BGQcvzsDkehwje32jpFWuSbhUCL32nmvq
z9zIeYYziarf9xeQcrpFbmJkjEYSNN/vsritYqvjsteQd+ihv7uJdNCuYVIAc7AqraJ1C0gk26kv
yQFGoWY1dr2qqcQZiU8hm6kVV6lrZJk9rgNQYNiakSBlpbUVcTYUpCC0VVDYZyZlzSFbgl8PgvkN
G2DUPs52YymyO+YOWufHaq5951FxmA/bVYJZqgkdvN8at9TLAJ7JMTbzPwcXV/I0n0uAv414UsQP
Wg4EGp4CN5e0V9xFydCAnUUMsExzprFiKRQu3v46We8LCDz5YfpppyNXJNfrijzeoQTtq1tS0VgO
wnfQ4TsUOtAnlt5I3Rj44FS5AHmHGMeuO+er3jmek6cqk0FJwKmXJp8HIJOaxhAngDUjDZuegnSP
GvuyXF0nqJ/6gEvrBqnXzxW7/kW/UPr/YEj8s6EjOvG7ZVFgD382jqn0bsUBgotPdS/0hEwVMFwb
FQ9YRyAbJ3bC5KOAWq+eWB9269fg5r+nXxAgT3Gyqwqk6yp9v5sOrdKf3dQMW5j01sUCxO1xvHwc
FBkhEjKcep+aPEzKPcCTgnI1k8vYIu0mXtPAjjaP9UyYEW+GlszqEpoLJ78mzwtBLpEKRp/Xwv7C
D9KKNw2FLQDN0yoY2k8uHe+mKP3bTD/hKt9Y0uBQGiT9160RF11PRkeF4dEKSvXicdZ7aNUd2MdV
39OQU7XjXDIa0A+2/VzhazBqNJSjuHd3EZztvl+gjDgZOkPQP2MslEl/XuToQaMZfdBvBG7dZc2B
dAEpT+gal2Ws8dJ/50565H9LjKOdnSGwfqQIUhzvnRfmw4jy9iTiQYA343e2AgKaEEinCduqj+Dv
vlTEgMOXS1+b6cx8m9u+uObU+b1U11udsXM6YXOYDZ6onIShK0GA+cQjLNebu5mcfqHM0SDI23BG
D+VaNiENVAisNcCA2+7ALVABVGT0c24OVNn2CUPswK/C5qAWm1mbzuRjJUZs+vKWcS97fuELmtKv
ICYTcqy1oXixyrUcUnPnB8yTv3Kx4DsDZH4OA7v9nSeJi/o/Fw1S3b26ugmLxI395TAhoMpDjWqk
R2/cuKx2C4piSFhyTrKx7HmyJqcH62e8brI5KL66Cj/tEj6tqnuzpW5k6tSjp4aDABDsbnzJcW7s
AD5KBDzKpxNIIbYp0vWT5WicEJk3gYYWLJ619qaPV7ZfPdQJ4WIr8F4RB+GZs8lxgN0txp+RMPr8
erG6SKnTJxcWc2t17IaL/1sCaVqRGG1qE9xitbX8zav1B/uLI5eIQSpLuKogFEl9lRgijeANmlE4
Vq6fan1ej4/TJmNAC7FLwoE9DyEpATfjHFdN2JZplWuIrxMuSaitOTK946Vr9hLQ4Vm2xPcDy/Aj
PD6rL9oihKqD0q2E3zd1BquIT+4uSnxffv+d6/179gfFoBDZ/5TMXsCdVwXsRfH9T3ZW6JSgazp+
kUqCIdzKNL1/N5Z9/vO+r0CBKNRtF21AtW8SNlIEnJETmJVDQfNEWsHK6vh3htHtdG+bGW8NE780
oJdyFu8esLbKVT7OfrQWUwdRhilirwc9a9OtXpE1Cls05bJIylhb9vPO46a5iM2u1sZsgTopsALy
i913kkEQnWoDRMCPBeYglxGA/+BTEXD5L7xxT7K7vSG4cwfipViFtZqSN91eQIimzWcKjdHnwFbF
Xr+YHCwMSlxW/oVr5YuwmX4kUputl5+jxitX17cXYRl/A22O/RfdzOBIro/22XrHTbkbsN8MHwHk
7uUYOWzWYw2LxKoPOtq8bEVgDjRuXlVs/BCOjb8tqKuKeFRckKwm1rLUSrOlmAS6i05hj/0k8C9h
Je8d+xRt9M8fdr0ng4bpYEMsbMfN2Ko2e9gaYLjbcHrkRTau/5gxk3twiP/5Bz36PseT5/FVeMpQ
qiF3P5AnSyMJO+u0f/CmcBCfZXlPIyP/AWC4RLr9tcAW5ohItPyBLwsAEis59/6iOBjsTMUsQCEh
CSmlWbOqHXmEbk7kXfrJk9yIq0WCsfE3U7TreM5JnYFJxxiu4K1+K6EZB4vvXerKx30WAgxgeMga
YKEStUR7W1e+f0cwtCqtUvRu7bpZOmK8SY4cn2oB/4uUcOj3zzbez3/Q5YUT8UHTdU50HDfGEeUn
qDZQczqkxvVsR7fxYX2iWqYFf4FA4lYi9nBuV5txpJaOdR0EJBfONR//is6l7xGOnfT8nK5OkUw2
V5UppX9pIOLkldyBkOFCw2KXHvldLFTHCoH43IF0DfSlge1xTkGeM52ENjn6DJuZpNX5mqJjIhXs
CZppLCMb4nzup6Lq36VviGcf6i5w4mHgo/K9LMzrxTi4N2GDiQezzgpSd9FkVXFpXlNSEnfxEA3a
Nx5Ex/cjpp6wn59jS2UAZh/H2IkWB/H8oC7u2mEfSa/g1PQoZ7daBtKIqjdvaU5Td44nH18XhVGW
/qVPUkY2CiTY+JP3ym7xpzbBeU4pA3TfO5zZ3IoMOzEp1MAHpk79ME2shgIHKrh83oGZH90jZQbO
G6juh1CknYwvM4jWxx1OKI3c7XMDlsw8FBx/TCmbNCzRBqjhqe9gIWgu/eRMxx0DX9rzHIoAYpCS
j6cokmV6FCe1+28wLJFeH93uPI/ZQjOm6mOSpMs2EXoGiV8XhM5iPuj1pbfeRvfeZ/H/lMvw+q81
aQD1/bzQrj1myiewEVvr202YV/aLAMhtO6ZRvWV/35tAKFyXT6XMeB/z1r7At0kG3MJ9AbmeL+ju
cQp3cbBdBGN686XLUzS3As4Y2icw0Br5/J0j+DWe5SQlTIUeusBPLOffPdPItxdFcAAhpjBOnZCU
mrldAiK7VveY4p2APlJ4H7sd8zkYlOv/ikkFhSuGvBgRj3gnzAquhOmwZ4Kxj8LjyS+I79B1flMS
6ZmOuM2W9tkvBgdBIRlwqXzRBAP3kxiKxt5BR25K+IlyBXngdDI4aUWSYxfVOaPgxsua6aLZjvb5
+jzAUQmt1drewfgxb883ceavcUbHMLgwLWcoXRlMaR8yE+K5tU9B+rxZ5C0WpqmEANSWqC5IRTAf
HrOXQAkAnmdsXSTx/pIfk+p0ALD9HahjOvqQy8ctQNAhW+lAyGnTqVqo5YXXSoLQqgXFqocOhVE5
hFtFdxxxR+KxWQVarCtlgNlIZttxF8zEbL0ijygdOi8odSl9eqKdwfC89xKmaPAICYYhCnc5ktqh
3wIp8RyzNa9PJlqAFUgTOo1dqKd2mQVhs3/lhtv4TXCIa17+N2mLIa6HIHirKoIHTIV1YjbyJRzc
SKdP8FeqlrBSY/2gJHHYXOMwS55XRuRzGxhe18UgX1S13xAssLXnOx+2xa2eJphT5njOacHulriD
bO157Nm754uXjpmeCRPZwDXKCpV+biEGMgSYPrj8ooDbeRAKGbqATdWfI5p6qlz3Tj5nYCGdsxPe
PpogsnPXeA13kId/KVdJWB/sQ6jHE6LLM3usgIOzMsbmFOAuH7Z5gNcGa1WWZ02liGWbQgFduFLS
SA6CskP6BccYRKDpr6u5RjHE2OVRO8QXfw4O20nENogigLJo+SjWzipIKP49ZuckIznXWlAnMUrL
EU6C0zWyW/bUKnoqdKyC7zeqdLsSyzuqThTOMbnkeSCvJ8YyP26OfMsVx5l0Z67q+w2KQE2zwzVU
RofA6nWlb6gt6kT4ARu9M9PrIoYKVWbT4Ygo+VUYcH46YXLtgRDmq30C0TOeEz8B3piFUKV/qaOS
Y12q+tK3PdTa4f9PIK8RtjywDXZKnT9SJnZNMEdQfVZjohSxPD+I57tBY4iX3jUcIxB7qiwiJXdB
YqP+GBkIme0WUQPXmVI02d5jRFTuv+JxA3Lpp57lbKan7NTa3vzbJKQBFFAehtZQiKmHVJjwCSxr
vm9HMIc0tmwn+LEnSKvYuJyIoLLpZoA9Caq2oTdZYhOlrsHdalkyqFNxB/IwmbufqLVxNprZjE1l
MCHlNgYbqyejw8Gtcw1sG7UDy4JtmetpIRf+IgxEwZ4/sYTuQNtRY4EJlAC8OXc3646P0xGG2mam
eyNy+YV9Vu3OTN+VqFEimEXQZiJohgtvUbgikX8gdtIiY4DFsTN50oSs21kw4W+LxEeK8lx6jdiv
16OLc4BzeDqsycQfaZtlSzZ3MG8b8AJGm/KKeVSfQ0V/a0h1JwxrjolBcH1n+aUgy8XoAg57DrH1
sgzLyvVJ2ZdfvNqFvV6UtRU9wEsL61s/GMM45GV14/3188vbjxxEwV4JsSES0ccXfPrRmBahAVQq
mRAsrjfTptLYm+jB+/PESOEYghrnScZJrna/iMU4Irog5VpcQ3JCIq18qP099m+vh+5186CFNk6p
HTnN19svE+RnGSX7ZBtbfWLUVOBPK5+d5sxn8g7BJ2bigHFOnamHTEiLGAe0VsZRmILfFn1pq9Gl
ZR/nU1VBw3bJ4MyAYQgdQwuxONI18UOTGSsLHL1bpPxYPT3s0feUAU1KEOu3oSMVirJkI9zIsK3d
2BA+3EBTy2bi6z8xkJnjrpBrA/6ErMJjk2dQeRNrNV+xvVMxaPJsXFE4zBFEHNoFC442bnAJI+Do
PoM1SwyvY1MVDg58IChTdSkt9uFRaW0QWJNisQzI5ATwnieQs3rT5vPDkkC5vSpHZxBnotog4Opb
O2WRWxjbcpZpqzmryWZcuhhTYLgrUf8rhgNdaQMLrtB3l6rN+XCBX/ncBhBMaVwJ4+1Fqp64EniP
+a9oh/GZxBwadm2e7jN9oVbXl80zNoePv6V4fDaWnU1fowX6cYvxAisGtBgYi9a2wwTuX45xhxan
vDwsdjCsoF4o6aM6dIQa0c5S8S4Bi/fiO80K3sbwSjnGqULHFSVCUEokzMNfNPBqx2UFgs2b/Gxx
xOL750VHh7yLnAYnziMgtmADax3QRAcARFe6BLCJSYZzorxgMUS6t0ZTCyOR5PBiXQZtDXMOxKrJ
uEHRU5+G+sv9cH1/v7Tax15lFSJ/odz6ixwoyHWsDYhIEeeR6XlA4RFg3eDPQOe5zF5ofL+j14hU
XKaZ431XVsom0ycGQ5uHEmteEpjOpBT9bj0FCVxfXo09lTYnMwByTW5yg2dhm5qcdBrAQIAywtDk
2Cow0KVxrCNeQITpNDdNyaDbLRSonhZQ9Bu6VwZb6GBoiYlRNzTZZOhvBRpHmg9kWT+I0JEecOQ4
LxMNLAhrtLD6JBUeYLwaAWbKF0Ck33k+jO+KGODFu2KXwVetYCqCLY9TOQYn75gO1S0/5T7cOTZj
jCugMBeyzcVFoihg4h+4Tj5QiXMjqAMFbDxbrZLCdVAyxDIaiX5gWhxT69m7agZEXHMne8HFYOHo
isS6TvYdSDayAEccJJi7UISmomRVLsQcuD8PTMuxuvbIvvPsscYeqfaOlzNsVz5HraSh2pvajoJc
aEWj/pQE+G0RXTKXVEyCy4KmyG7l6BjAVLOHScr771SDMXDx/BZKJi+WlBiVwmnk2PVnz+bn+/vX
bj5dh+jfP5QDOH9/F9qlbte1f27NbCxLmc+Kr/iyDRld0jgEMNN6FufwU/kIR9B1ZdbBNYHEz5mi
C7CF1IJN5FB4xujF2bT/fWd0wCFusSW3Zi1mDbOnowRgv8Yg6H8qSF2PE3x1WeM6BqQwAoyFNr+x
jSNscrbmdR2yt7NEhDec+eBPiY5tDJiJt8iiZE5pNh1ONJdiwT9xwg4o8fRkg++ZLjmbh9mH32ZE
/cVNTJNefjHOlT29Mo7MaN+GsrXZjFatyfPtjXX/atxsbsKAF2Xsu9GrWCFDfbh4CImRAdx2rRPw
N0OwoYHQiz3EdtBt6fX/USPxzR3+kh1Wn4ztXcbQlE1qhL4+OZdoEb/GLmYRKEP2qkQ7FslDo+Ru
y5bswI4e7M9s8VbCL5aO4kKrBO8JHaBoAdM22t+ksc1klP6P4Z5l3YtreV6OVWD0Rgtp3opYdIMN
WfCiEAVycA6tLWTVsZwVhRxtACkPO0rvjdOM3217xn5QnxUHews8T3uPyWcnDoIC/7OUWneT6kbL
e8o7JUxkRhkTmxCQ9ECIDFR1YNKy7LBPnwQ5mi0m5xgGYXY6u7OR9e2a4tinpIA+lwIwkd1JdY5Q
9tVN5Ab4juEluKB9g9JV9wvcCg9BtwEF4s1FBN6Nl9FsXrn/zUbK7xwWE9TEW1uAuPHrN+7tJlPd
nVKRl1e+tFF8Wpx0/S+riC3bvAY8r0ZP+1IyANlsP0PPLZMjmP2CIJVnDD1kHj2O6OfOAvvewDhZ
HjBPibOQfZ/9o3fIHiIlcqjKjDqcb2Gd61F9+yP9FIKATj+19xCvzHWKJEL9QePeZePKnf8FD26P
H8ZWGc4a53hVlzctSyljXDHiHH/rP0JfpfLnG+RHfAj07YrGJyx67hvBTwCeK5i6IA1U6cAvQYol
WH5qr5alutXMXlAvNlbh0MWnvYdr1pXFlLuoKl/xw3rhj4jHXCl6zxYGYd2Zvhty+t7YyE3/JnT8
s9rOG0H1Pg0kQshSA+Noc7WiPDSuGehJa09nySw859hCk3fla0Tl83UDJitvFKsXKiZKvFhi2G64
1HrRrxfu/9GFWf3mtNlxck20QsMYWTrH/JX48ejWTMN+c4Z3WDsoI5YiHyXoHVh64/5ERrOongn0
bGtqpzesvH9tfc4DvfuCiATxXhAh0XSIPw9SN3bnYhgGxOUi+dEJC3S+syeVPfoCVlG7rqNxKdJp
7ofZ1yC4E9nhrBivFmT1v+LLxhbm9Jc=
`pragma protect end_protected
