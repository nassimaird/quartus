��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�˅������d�xp� �5��B�{�	e��Hk�Z�徒��{��\�83,�p�)V2V"'������'v�{��A��L�J��ʖsk�eRGAO<M��a.p�b��@�@a�;Dep�r�p	1��"32G º��*ڦ���ƫ�r`�c�}_1������	H?���}� ol4,n����������\p�kх���F�y��f�T%���^5�����8
�2j��pVq��zK۴N��@� 0 �	��ev����m���z_ws�=����#͑��]�Ţ���FC$����
�4o��3[�Y3�v��� r�'��̷�l���S���W�v����E���1��_���Ѵ~���;�ﺴ(ܢ]9�\h-m蹞����3���Q�ó�?�A����Ƶ�̟(|����g��~�Q��6�tg��}Q>�CW��k�9����ΨˡI6I���OS5No��k*�D��p�(ޚ8�5���6����I�0�~����ǏFA�2�;ҩ7^&�'UNg7���ZE(�����
J�E��B�:w���'���W���;/�R��y�p����r��Q���Ĺ�х��9�v|e��E��(h�,k�NNk��xL9ӌe�9:-cJ� ,��[��.����r�A����eA�v�)����8j1�A�ƨg���o��������Ƨ[cP��^��r�Qfm&�ؿ����I@��3Ml����Ɗd/��gčZM��H|,*-�r|��bo{��@C��P�eV�c����C�u�μ0�3�,������N�X�WBC-���2St6�8� �7Uƃ��rX�p����4�P��V 涱�P�n��)\��*՚�S
��V����RO�����d�׾�����P�䈾��*�A� 3�b�S�|�>|0�X���w�g�g=/�CmL�~q��4|S"�p�Ń�%Dd��E���5��@}�n4��`���/�z4�5@���Y��R���ѕS<.���Ö���D6y��X�����K��;Y�aH�V�ik��p0�P��˚(B��Ȫ�����q�����d�\�С��J�MцQF�3�G��jUQ�Y��TU ���Gh���5?e�0� NV��2�;I��6�i7�e���Dsc��ӻA�S��'�SqY��EX��J�X�2v��vB@�El,ZT����յ��l�d�"m��󀡼�M,��~F����������Y1
�Tr0�90�����[�6�5��nI+��q�Ē��ֱ_��(v�	Ea���2�-�(<❬������7͸i��'�����T���A��В����ݺ�fQt�E)jd��L�'��'\��CG��@��s9��2/�T7J�4���1���sYb.��Q]���њ�bd�����d�~贖� %����2�l漯��~KX���l�Y�Z���J��h�P`s�lS��,k�GƐ�x������|�E����}�x�ސzZ��|%�S�
Pdr�|`�e�0 8MI����L{����Z���>����� ���e�x�ؒQ3_��?���������,|�q���ɩeXNFUo�}��r�dp�M�̒�m��.FHH$x�8}�ByO#����A�?`���h�-�C'o�e	��/v�y!xQ�������n�������E�n�c���gM�`�y��g�P�D6d�"��ԅ��6����īM�x5� �W����	��L��X��᠝ ��y�pV�q�^uo7�u���k8��߾�4K��Z�����pٮ�}��4^���/��(;��v�_��{���ލNe�S��r���˕X݊��1)G����H� ��\�/�Eܩ��h��A�����+͸���|5��!������W�	���� I�Og �"�鹪�
8"z��9�2�R��塓J�i��.��b�A)_ؿ�L��uW�g2#ރM2�͑ک��w}�E�� �@+}�_f�|YZ����5���a1O�@����u���W���P�q�	��m�!�n�ix �T�Y��N�/�a3��@(�Z�!���DKM�a:<g�Ȩ�e0H�H�t� !vX�w�͍��4����ұ��thn�^�q��#W������ǝP�L7	t�"�B����ɜ�����RT!O8s�[�MN��}iI�yHQ����!wveggt���l��C�������ޓ;�����ZR�_�\Q��tk��>#B�V�x�Sc�N�e6��)�.�X7 v���F! C5���Vo�g�����J����,�]�8s@�l�9J(�,X����d�^��v�/�E���F��h� %��3�w/1RK�0�)��ŉ����k�� ۰/�ưl��=�7X6
�έ72��A%���I��^�K�b+4�^IOcE�_q]5HP@Y2����Cwt=��5��!o�%(�������˚��\�"4�wÂ�MI�K>崲���{�U�9�8�+�#9�ۻ�e���=��Ht�;RJ�ɪ]�_�bp���*�!	�8�����f�찄 �Uխ��ɱ��`�@���ԓ����],��W��H�r��	j���yꤴ>�k�����/���]�5Z<�n���@�_E��%9�yd �M�4dQ�O  OZ����οgO9%�U\t��A�|�r��Q��vX��h��O.N�|��L�r�S[���\��?�+/�������"�x n#�v��+vҿk{q���^��BߺJ���(�r6��ߊpօ�Keγ���c���
�1E���!9��4���%��D�Q������+3S	޳ ����LKX��Œ�<� c�u�`����������Ä0x�[���t�L�y2��6�D�M���������-�o�T*7�Czˉ�Y���R���J�T��^��{_M��D�,�$U�.�vxҏᰯ6�+���4�a9M|���U�JaQ��3��I���|]�:�!��9V�jLP�e�����8a]Eqq� k��Sȿ_���d����"�^�=B��z��N]�/�b`s�>'�tT=���׻��i`v�y�V�,�Y�֏`�J���Ex��]��f1iFn����@�ݥS5�{�ѳ��ӹ�Y?r�5@:+�K� 8�՚Ҷ�K
����H�3/����\����ut0�ܯ,���F�0�	�#5ZHT�&����5�pV�;Av\K�I�`��J��š4��o�f������à��5��A��$��75LF����清@��9:^c>LK��9�����Dk���_�	���r1���Am��7��6�k~]�����&W�_$o:�Fl�F��`��SGw���;Y/�4FP�V)4��7�E�!�ۮ�~�L��h��W�����
�:���z쨵��'\X �Ne��r��\�����x���!NX��H�h�b�I��0�[��`J\,l^70�J��1�	��?�L�vI�&���`\a�Ӫ3�BI��X/��)5L7GZ'}X�qI����h�^|�3?-�G���`���'����s`��h��B%i����l�����[�v��X`���:��IS�ٮ��c����� �]����e)�a����f�b�tkc+׎����#�KڐA���*��H�X�(z�=���K�v���A)D�j�+���x�CXI*��	�马���e�*�A5'GcЧ|�A�'�( Yƅk�@�0��J�J�'l�R��7��aj�O���4�`�I0CǏ榾����n-@d��T��5{X�4�p�*9�숣L�m���Z��L� ��G�ص-��y�-GB���<�����pUe�̙������R����J�y�W�����4uCu½�X��EF����w)*;֧�k>� %Bw�K@P}�~�@5��Ȗ�S�Rr����/�4��	�:��ޯ'�[D%��쇊� ������^��� P i����X�l}s�,ΗD�����-VBȩD��>�9�n��H���y�j�*����U�����)��s�;�TFTU��`�y��Rhc�b�_�+I�r��b��*��1����j:O�'/���'O���l��^P���w���:��,�Mܺ*	m�p&,��S0��s*�C/�	�l~�p�(�g����~cm��/4�G����ϥ)��EC.�>�� w���v�λu{�������J͚����n��cr��K��!s!��{�2s~{�]�3o�Qj�U��)|�m~8W��X����\
*�|�� �>Y��[08xu��5rN�L��ł~��,�dBy�da�do�>ݢʂ���NT�a�R�3���O�ǈ}�(�k��
��"���Ħ �g��v"�*zcF��mɕ���,�o2"��WևV� �ar{�n���:��;��*v�&Y	&�w�����mwe%oo_����ʵz�iY��3�7SY5��B�D�J��W{�k\���LØ�r�[��ל�r �l�(�Vxr&�a�Wm����&�;zhJ�)̉gl���v�]G�\˂N��bt�rh~e[��p��g/�\�gpi����@�k�̂��V�����l��h�*�QmH�"&�Xρ�����y+7�I�uu�LE�a�]m���6L�D�Q=��s��0�)��$$r�(�j�#E�o�ϑ�$���Y|��f������;ĹQq��r*�Zg1�yUM�\��@]l��9kv��ܚ+Y�d���U�ꤍ����E6,n�]�-d�3�A~Õ�d0v���x�n䳋�y����.:G��g�4�aƌ���1QqiJ��'�ƴ(��j\�"����jgX��C�|��Ȁ�4�
�������.��Hf�Q�����j 	{���6y���d��ٓh�1�>�[t-���T�X�.�����`iJ�AG|E��M�SꌕE���'�(�Qi����&���oM�X2��LP�F����@ݳ�7�mQ1Jˑ3�,}�Ԇ���ɠ���Lȸf�s��cڞ14�ꗇ-���G����!*IԘ� :yx���JW9�Ԋ�HP�uD�	Λ9))o�~�����d�M>��l����Oj	��ޝ���g�u��Q��Ct���a{���(�9i]ĚWK�.��t[����x��H�z�ܹ��T>TXł�_l�>�.�j�6`��{g���t�j�-���!�s2��ncc��A��5z����,�Q���MKK�z����9p�8 �I���D�s��^��C#�T�({8���@[~������[�}���cy�Ұ�B���B����P��>ϥ�Z�W���V�Ew$�\��>y�]7���ڧ})̏H:�ޗ��#�4��P�I)m�$�V����_>�Pxtk��j�&����e=Д�']x;7�����ߠm��G�F �P�=Dϵ4�;5��`��fo۲؂(�P,OZ��s3[+����������菱D�5xUN�j�@B�J�L5ܬ�B�6�t�#|�Y��87��n�zV%�T%'�g챱,x&3^0���]̽�_<އ�'D���BA�G�?.�)��*p&:q}7@S�zyL��dM�_���(t��ri3�|�8�(1��H�֧��\�1�$:������]�"��� �׎	����[N7_�#aT��p�2�o�mO��tbH Mr�p}d��c��bFЕ�C�;���w7;�oe��9�Rv���}��M[�Pj�J����.�YN�Nςy��W���}�񇠔{���Y��c;ދ�~�MZ�}eu�5)�$3�k��򵪃��J��:��9�D��v�ɖ�R�Ɛ���v����o������ۖ�g[y������Q��j��e:���f�` ס��eOlӧ4��E��C9���GM������1���-��,W���l(�O��К!2��W�ߥk�s�	_�qJ�<����#W 5�c�|g��v�B��Õ���C��Y���ܖ\к��(!��E�I�dl����x`C��6̩��M1z�D�pw��&�4��	��x@�9�0M-�M��D�L˖o4kU�|�̜�g �Jb��f�<*6�yc
�>�Q��0Q'8>B����н�i�o��	��{�4LM<��݉�^�m�.o�-��uS��0#l�L��g�#�PB:�l�klU����?l�٥t%�v����xTN�b�~t:׀cB��C��8��Y5 P���]T�4�">"�t�Z(D�dvJޝf��=�{��J2a0�Y>�,�m��U����R�S�\6�sW���f�_�YX�7Y���(w
�^p�@r�������`���ȓb	��"�𻲯� �z%�v��]�2L0���N����Z3c��ߴ�;��B�\o�	���""�(����	{C�T���/WL�*��mG���%4 ��+����
D��{�n���돲��"7�aF��/�Ia�5ޱ8E�g܉^M�:�{�7bnT�(F/͹��ӝ�<����`c��>ZmXq�%rM Xm�L2Z	64���RK���a0,�\�vR��؛�%l��ӞG�B=IkI�,��_ï��&��Ȳ�s�c�Ǹ��(U�:��;�{�{G��J�DW��_�"L�2�D�Y�n����H2ߕݑ-�&Q�F_�r�3��{=m� �8;U�h> 7��ʛТaF��'�~�v�OHk�w��,��c���wB"G��zD�w����z"A����H/?}L��ٴ=���*��NQ��I&�+�o=_w�����L�D�$����@?!"��Hȼk#�jBNό���?`���n>��YvAF��|Nj�-$�D��a\y���T[����x]d>^��$�W��mw1A�B�`����CP+����TZ��	=s�}3���*:66/�e 	Ѐ��|,͏�u�����;H[���,�?����V�Ş�1�˃mw#�M�/�
���>�J��=PX6����ЩQ��Z�z[�F��A����#0�wL� ŶRuc.��X m&�R�1�	��l�|��^���t�V-��B�V��O��Ύxԯ����9� OƦ,���;���IŅi%��fRH'0�P��~�K <�+�c �l���� �O�_��W*�r���y��['�9�\`���1��Q%���3���d�p'*<M��V�/^�=���k,����օ�Lf����������ɱsM�4���U��e:��/oa�M��s50�V��RT��ˊ-�4}���&�rͺ%;�����~�VR#	K>��2XG�N���@����]����#��J�h�
�T\��S<� �m��D������C䜖��-:��݁>
M���0�4�vݫ�MD�b9��t��ѹ:F(���&f#j�v��4<u��{k�bL�������G�z+�V_���j<��v�H6�JP~�z�9WG7�2xim�U+Rp1x؎±���X�/�a��6:��pa��0e�[vk�T��Y��'����I?w��=�q�k7w�LxCV�6&��J�b�k��S+�iĈy4�n7��\lM�Ҿ%��0���S�ڿd�1�!��yAȹK���>�,�zҷ���)ng�����t� �G'ϧ
GX�:�򐰿1����z[,��ʴ�n���oL/|�FÕ�Zm$�U=l�+2�w�j/�UP_�%3�g��q�G�~�ھ�N.�=����r���	s����t�yvb	�6󂽿0*k�PK�T�i��%-��B��{��P�#�x����ȷ�sr��� �"Y�{h�b%�B�c.�L�v�gwmrGzTN�����?sF�����σ4^�j��2�+������!��qY�4]�*�����Pp6�[aஉ:CW��!����kp Q��=���
M�b9���3��/~���L����Ԝ�*)���o�j3�zA�-�W�/b}d��ៅ��X$x	�H���,���Ĳ{	��s���*����eTଠ�5(�'��z�þV�_��ۀ!���8�����rK���c���!�%hk�6x�H�ٹ��앩`���l�E����������#�OY����I�2�)>:��\]���X�p0��O���E��I�D�q��^ˁ@g�Z�)��*�{������`�s ��`~���y�^J.Px��]y�w��L��w����K�����UØ�3���;Z��E綔� ��%���u��{����4_�c�(�`F��U:�X��Z4	S�ȏE`���c�$�i�����c��n:>`�*���8{�V2Q5��	a�&�6���0���[��qqV�uW���_�O�D��L�4M��h;�)l\�o@���jx�A$��YV=�k�{�W���U&�� ��@�6��iд4#����\�l�"6���T:`���ĺ=��,*�b�59� OW�CIF�*�����.#wޠ+�Ӷ1+e�
\�1��q=`�<�]^O��o��}菴��E�Ĭ���f����P�c+3Wlq�{�z,l��4'��b�q�j�p���|BO_�[��k&mf@
3�^�*x�����a�1�&|������qR���KpzW���pf��|�i�A�Q��L<���5�˫d���-6��-m�����V��ihMBD�[�y���g1�T|�@��+l�jU��;�ٿ�.R����y�h'��FM	E��%h�6���F@3�UP]/Z���e�Dm���5�E&A��9��{��w�!jbv/`���ξ^��5��*�l�������
Y�"�������oz;"4�Xo�{�}�E�(�'����{�w��b)l�~~IK�	Hu:wڤ���d�jj�|�/'��n��|�W�����q����	�������!���BT}k0�eI��z)��} v��Nip^��V��;�A���Ў�2�,��9��V��)�3�n$w��H���BP����L|B��kB�fn��ͫ�C�	�r����K[vpgՇM�k�yg�J�A1V�<�Jʩ}���$f��B-��eΧ~
�H���i52w�5�|������_��o:Z���4'���WR�`�oX�<������w� t3���hXU��3O]N��!Q�Z������U��L�(rsk2��V3k�:�?2�W��	 MQ�ϛo0U%� Y�iAp[%}�]z;Y��|W6?�R�	��ɇw ��w֋s�Ŏ�r�Ͱ����!"�Zkbn?�B�x����b9�E=��)5$��"�x�;���y������p�x��|��3�c�|n*��ӒhB����Qc(�'�S��qL�E��砶�>�g��] XݠUi���	�pg�l��਎���w�*�v�����-C�\�ǪQ���5��v�Z��9xb*��4�DŅp�+7�РK���g����n�Ň��qW,A�,WB�3��8�U/��$U�;1M�.Z���_�7/��Z��Hx8O�9%��.ڿ�s��$�Eߑ����w/�M�6R��]�n��T�zL����>)vM5�
 �;@�w��%>�9��6��f����뾠�=PN۲ՁnL����(�:."���f�s���Ӻ_A�m���?��Bj:/RuoKm������Lw��/S-��i ���zS�~\d�B�~�9K����^��w�`�5�����
�z�L��Kv}$��}�eU������[�I�Q3
�'�Bcv���=��!�}��â��vYNg�JrN�yw�0��H�%6����H<���Pc��!jd*��f������|�}L~v��i�Fߜ���4-�/$(�\#C� 0��]�[�3���3�щO&�&�y�K���f�D�IG2��F�'ϣ�^O��1U��G/%�{|O��,�xA`�	N��l(��c�<8(7�f
��i�VY�=��w�Qf�*�:^�N�	U���74��u�:�{/���RYa5��e6gf_s��9���ae��K%@�S�%u���f���y[l��+����J�0r�5�+|��X
���>�����X�bFY$�)\|$"�ޟ�P&~6��\'F���'���}e-��h��ˣ!W>�`�3���e1�%F���oV�=�RF�y��v��r�o	Z�^O�S�q�x}�x��M�=�̊���Int��IFi>�.qB@�j�1��!��B���e7�=�ꖮ�T���y�\�;��#�Y��K"��P�3n� ÓbO���r�F;�����vT-��a"�E��)�%H?�2�������t
L&,װm�za�s=![ǹI�=��]���c?p!����]q�Ќ횏=����[8�AH|�,�U1��oj�����-b�$��m�ۘI�@���V�����%/�%��=9F�o��wٱ��ŷ�J�Yq4�@ e���ʀ$��1M�J�����ڌ�k�S��e��3p!�6�~A�`y�;>�����y�L�C��B)^O��Ⱦ%K�b~�\��U�Gu�N�O5�n���_mL���%�3p8�U�3#BՏ�%��$�Ƅ\��d�W�7pW������'���t.2�yQ�}Xz�&H�`wQA�H�?�\��P %	�)�7\bA��V��M0	n�Z'^o.e��ѩ/��PoW�+^�e�_z�>Tx� �U��ȺI�V���	;��qB� �RϠ{�mv�l��2KJ�|c�1V�{� 	�����4�ʶ\� �DGƮ��;j��ud����f�I̘ٌG
`/�v:P�d �Z�� ,y�s,�
���tm)�K>�����^LtsEE��|�[���	c@.!�֯�ڕ��-�?��H���=�Q+wf�@je�l�j-��vʆ��]��un���s�3sp0���Af��k�;�jYZ��fL�c/�⥁��~� %W<�bn�S�n|/++���_nj��S���NKʦ���GA�o�;Tf	b�vh��He/�Y�����4��B��~�e=9�ґ�YSc(�J�10�%UnSAy��Iʞ:����-���l�9ˢ�I�5H�����[��Tu���6���([�U)���`���J�������|\e��W�\�J���\����H�;{3����H��	ݎH�@����j:��*��ʌ�&�����8��O�"�����#���&{�����&��?�lO�A�:��w��Q<�̿"��*�ݠf�Z�9s��Y,��J�1�z�+#"��jdB�����FP��M/=?�)Y^��"��?��$"P���55���z��~d�8�3��SY�R��z<�.n����q?Btew|���L�x�ns&��
J�^e���h�/?G.��Ǝk��k�j���Ini����υn��F���j0�&I��w��rn�-��v{��v'��xs�cxz���>3V�X�l򄞡�L���\� ٧w1W(d���vG�&�3��5Cy��c�XSJ�/�w�xgM�=��,��6�H���O���Z$ˊ�w��ga����w�����X�DX�&��RXu��ɻ��̑neY�M6���A/�i���+�ت1�[']q�;S< �%M�:W�s�*��CF���$v-�("=X�[�2�x1�����:��B�`\h����j{?���[A�TG0��W�����Un�xB�5z�S"���%��fR�n,��&����hO����C(�%/wi�����o�-�Ģdၷ��S8z��H���ʔbY;:x��nG��`��'�b�ڜTۡ��7V����"�,��ku�e�z��Uac�+	,e�@�]�K4˾�/�#�$XS���e�-���0�����A+�pi�I˜F�&~`O2�$x���_� �$}�?/��qF��q�㙗D�3�J݉ǧy�r��{���Ns�-WS��G��Ѱ����\�MO��ë�Je����S�����+M=#�vr���w�GK���vjL�l[;O}>	�͸	��Q�ĳ8�δ��	�ʛ$h���h}�3|�n�3ƍ�w[�z�Gz�D�jv�9���dH��֩"&��r�W����^̤�AZ��*VwJ ���Uo'��X�� ���M���	^��W9����[<Z��X�q��H��c|�zP ^H��-�-c����J�d����$��5� �h�7��V&M&+�_��i�.о�iWe��=!�D�`�7�PI�^�i���:�O����6~Zc.�`��c���V�#��@�j�w
��،�K���t��0Q�m�cF�d�<cJ`���ڧ9ɜcf�������*q6&d+|vz�*j�L��Az�<q� ��.�T�Kx�7V��������]�1$ѵWǲ��q຀�����8Y�gi�EgC��yA-��.N���#%'���#��M�U��4�����i�W�b�^Hv�It[���h�#���'�~v�����é+��C��z2A�� �����J��A��?�s�^�p���!uNRF�����FP� |��̣���t����ƨ���h���`�<��E���_�4�e�ҕ���M&E&ȠRe�|?������9���j��
�Of;����&�7�G�cVs-(�֓�w;��ƍr$�҉Y
u70�c}����N��DH5�9<,	9���Կ7�v��8�*����SA�Ĉ��tϖ�g�j
��(HC܇*>D~q	��Ǹy��K��I�㯆�SP`�������dZ!�]�5�y"�|�,����ʢ��o�]��OJ�6�6��N��qO��d�h6�g�%e��g�n:�z�^�X��)=dk����}��^����}��f��,�7,$Ǘr��շ+7L��7�y���&����"���G�=$�p�-�%i�owL��쓚�{|+�o���
b���y7�Y3�+ZA�'�b����9mx&��8��^�5��IF�Bw�)��cE��e��0+���ALMj�[w�9-Er�=�/�,d$9��ƹR?@�)�nu�.��'w�1��A2ܔh4���:���Ē�M�,������X�/s�+�������)��OI��ì�1:j��E�;��{��)��˜*;����+֝Ȓ��~; GF��Q�i���5���K�A^��ϗO�ǦA�[Sd|�?ߥ��UN�a���oo�}{٥����G�g�������F��/D�#τ]����/"���e��7~T��̈́΢'�k�	F0�#���q�6����C��Rњ���� �8�$�X�>������p��aP�D�
�����F�)��E��n	�Ճ�n��a��6VҤ�"��/���ؿp����15C��'��n��aP_FE'LL���0���8�lbht��Ⅹ�%i��m,X�Y/��|�e�t_�>�mlP���e�
Q3eڻ��%�񣜛a2X��t�@	͎+���o�~��Cκ���Z6�����s�:>R;��;a�
�F������x ��L_q�Ї���{�쯂6���K�[�}h���3��ar�J��tArX��W����7-�r�a`��q��}�b"�R(����~]{�?��P�ZS��x��b1p��p��,���:��(�ψ���1r�,��y
CQ
��\_o�8@{��G̗��!,�7m�?A!��z3�:�7������罢jR8B@d×��Tݕ���j���5�<:�G�ʶ}�j�뭫܁;�S'�'�$�0���O�ݕ�Z:�G����k[� bL"r��.��\�2�N58�h����&����uw�e߂��6�/���g�!�"�x�ʹ\���`p����*����ƭ�J�A��x��߅,�u�K/
e�YՓ��ɏ|����s��e_Ix�[$T���
{(�Ut�2>��R����S+�,Ts��?�]�hқ��3�����M�n�͐RK]���3N>����z�vy!��'�/�͇4�%Ï�S'! �J�F/{liDbI�iq��o������{}�(��Y��o���n�_T���<��z���% ���q8�5W�l�O+gd^��X��NC�7$4o�x���.&�m�4G��<J?�-�x2R8o��%�=߼���`r/���Oi�>P�6����<��b������Ԟ�?�q{�O�;�O80�\S���#��u4z�v�Z��	�+ՊC��W�;�[�`6��+̝���Wِ�k��1�ë�u���G�����w��2n#����m	w ��j���MNs�yk(�q[^u���ހYC�uF�^�d��E��]�k	TK��-�I�C�4��J���y�$#T�x����.H��P{L>��y�Wy�������Զ�34Z�/Ȭ�v@뱶�`��)��!���҆�f(@�eP�%���onY���h��"�?����Y��VWQ�Z �Y7݅�2����g 	ca�;3ch=x��'>D������c,3��c�o��n2#�	ڢ���S.��WU�%�(�� �~3�8���+�Z��,�-I�{5�$��sE��b	,eĂ�b�a�y���.e����['�>a��Ub8t�q^���|�A��h'�; 1=�Q����V���de��qGz��0��$��h*�Ѫ�w�J
�i�>d$%�T�B>�ж(�{��i��ȇ*nޔx��ʲZ�g��~}5oT*�?�tɾ\,�ᗐ���͜�{J @K���mݽ؝���!��X�w�7�����W	��$M@�Tә��~F�����$��=Pl��	�1����'�&��0/N%&����VG�F���v=�����?��;񔛨�kQQ�p�0C��N�Ħo�8�;[�G!�I���!r�ص]+^c��AC�y��*��`����qVO 	�T��8M1�A�蟲|F���otڬR���i��4��Ӂ�-k?���SsoX�5n�3��e�~K�x��7
t�n��=�ceD��(�-�)����EAI�os�'r��7��Y%�2c�N2�	C�ћ�Ӆ���\��tyԲT��e'�f��t*��B�l�J`������On9�㹼�3��(���rd�	�>��#�-��hk9{��&{K4*��{���a�tS#����c���?�,�I=_�������u���p�ŭ�m�;�%6˃��]�yOƹ%�<�8M'$���9�8��c�;�SC�@�+T��j�m_n eNe	�oɇO��HV��Q��㨢n�P��+�y�Ъ�ګ�ff��*]�A�gꝺ19H��T�$R�;O2Lo��
��
�*XkF�!��o��"�>���D�U�O���C�-V�Չ��L���K��B�{;@l�wٯ!"g:�[���j,)�d{L���؁C+tG�pz��+�8m�*�>�@�@�4���/�IPE7�K߾��T�F��B<�]g#Tə*�?D �/�wIa��|���ˡ)`�	5�1�أ�'�s�V��@�ھ>��H�����G�8Z��'�ږ��F���ZW�5X�1Fm+V���Jy8RT�D���T��ӏ�P���\��o�(�A������YS����ˀ�5�u�R�Vp��~�	�ߜ:��~?�N5�ǀ-3�Lhbb`���`NI�|˖��a����N����T�}�ϳ R;^������i�����,�Ed�(��'�K�S�.é�/s����MN��	P�(T�@kS�=u�U�/d��ۘ�ِ�N�3b�80�6��:��/26;��=���b�]�y�i��t�㦲m!�0�ȯ<�i��e���&��Γ���U��+lW��8k�m�`�ŵ�;\����A��7o������2\�	�� �4F]š�\�A���ŝQw}|o��ױ&����<��3��7�w;�+�&����XW&*RC@lW"lz�_�e��2do��՗����B����-'Q'�<)�7E�#"jU�!�&��K�;�{�3���j� S��hݻ�a@��j5�n��tq��.�VM(8t�L�%�͡(|Gi� \�zQF|�YyH8��Z�:��O�Q:�.�u�MZ�&�=�A�j�8��E=�O8Qk�bL��*�\lDpV�C{�{Vb#ߖ� PӍ|l�=4�Q�����e�M��I�(�W����<(�2D�3ԑ��W�v
 S��zr�Z}�u��:���Cd����+Sُvt�:� �uY��>`Fe�p����,��9���3���ZA�J�I���_e��"�"QrZ�W�0����S���u��n�B	A ,������idv��w����
.9D��Q�-e��=�G����
e��Y~�?���_|�Lh��P��|����D��~6�6����"������1Y1N�WK��X�_����/�v�W���Nr����EǼ��d���$������@��[U���A<�9�W�4@��`N�?�	'����e�G��b(�Xb��!An37�A�U]��N�!�:[jY3$���xc��/�a�
Wf D�7��gٗ��YXM�����O  L���G�Y$��5����M�8G�	2���/�����7Z +* �܎.+y�OOQ�&�r�{��V�7	�U���:��ѷvIg�j����E]�����m��^cMg.�g��QgF<����C�!��	�K�̸\���箓�f�>9Ǫ������w6{��9�i� U	��P�PO*?�����lAq�U9��HB�Y�[�fS�Ps7�"�����rļw.��&�=����үP�o�S�u�e�E���!�<E�AY��M��f��g��f��!�����,?F:N��� ������i~H�ӎ�$�:ɌN�TP��^<0p��=~������D۝C��*_^�$� j\󑒬p"E�ѳ��):��آ���!%*���<` ��!0�ga��`�	���+���:�w۪���?�����IqS���3R����>��}_ {���)���7Ti3�tÉ��G%�;o۞!yw���0��<�Q�����2�ŧ����Y�����ɐ������Ҋ���EK�d��#"��rK�.��yy�h&b��Ípѝl����Z��(��bԵ�z�ܸ�Q��V���be�G�Y�R!p���{��؎��n�V����
2K�V��^R�+v4˜#�Ϛt%�o��n55hu
Ig���Ό�E6AP�)`�F�ߝY�iON��a�8��3��fS]�Ş�� E��>�m����߸�m�1��@~�z�\���A���Q��E���G���ǣeت\T�8�8��}���8�g�-�n��/��Fp
��N���?�p~��^�Q�
�R]����(��ط��-V̻k�w��N߉��ٕOǞ8�D �8��c�R�M(���Ȭޅ�-g�o"2�mF�Zx!���Y�b��6A�S��Y�ym�,J�YR��y܃��]C1Y�)������ݢ�FQi5}U#�d���p���Ο�,���Dȼ��h仼�4N=�чO�@�k-`�)O)P�Z)��ql;/ޯ�w{i�X��">�r1��7#�8��h;�|N�^�3�@�?�q��c�A����J���+1 	��� d��X 	;�o��h��=����jL2��ݻ�Qvi{	j[6	���ǐR��/���{�p7���8ܴ���dM.Tev�/QKM�2������y�h�~�p��}�L�quz�S7�trݵ�Zka� �>6� ��ZkLhW��%�_{��7V�X�ݎo	 !�y�neds ����E�G�Q� ��ʝ�,<�'����A쇶�'�;���+]�����������2v��M��ƗI0=r>����ś2�!`~�V^:���\d�U���y�蜨��~���J=�*aпd�*��y>�f2H3�W#̧��-�6�Fbj*�{���j�Î?r�4=�xY=�q��jӀ�e2�B�IfD�u�-1�L�0ǚ����������� cv/��2Ϸ��H^�=��d�����!nz�j�����jY�袶��8�t�ի�����]�S&�Rk_N�&[�������E���p��V /�{z��p�眥f��t�tz�NT������8=|m�t5#�ӏ�v8[]?��� �c)�$����"���)3ߗ{%�"U���
�0�H`����h��e%��ʂ�/(=}���"�i	y�Z�w��@��)u��x!��/�V�(��ؗ�4��m�Y������e?ø�3��ea�W��Ki�eJ\XE���B(9��Ȼ�Q���E��e��.,�蘨[H����&�L�L^����|Mp�zl"WӜE�p���U.G��X��֗��3�Բ��ph ̿�D��-���4�c`n'd�	���Ǩ�Rt��A|S�*�|A��.B
hNUyY�e��:*P�P�3㤑��i8m�I5j�ϣ2��7﫪�kutԡ9~�[�?�ۆ�³Z�$�ݎ��>w݊D|Dț�ڍr�3z�_��ln�v��5e�.w���vn@�횒����A��6��ġ����>�W@{���^p QV�׸}W'�U�g���[�����Qw�U�>-�!ט(�ߓ��V����Vm����9�������� �8Q��y�����'1�f(Γa��9�w�{�m���}�@l��>���ud�tE��{���I7")W%'	Jwȣڀ"�lG-�t�|���QK�~M�A�0ȕ �R��I��GCb
~�6���*=�E)�̙���:�WF�0A���#�:[��U���nu�R"-����d�+���%��	�Ւ�7�yAphG�W>R�y�p���I�W��φS�!U��_I�|-!7��S��dB8Ⱥ���;¹�u�F��u�Ѕ�sH6����N���^@d� <I@�'�h|$Dn�����-�ǣ�$;42�v���#h���7�S�W��5�N������X��#�����&���}�֋�+�Wx��K]����
J�B�Wi9��7WzV3�qZƚ�Q�G��s�[�3%�φ%1�7��/�imy�Ўc�<�p0F��_&���G���� �+�)$g)O9I5C7�<��,T:89���+�}0�s	�m?�O�?i4�U��	�S���K�e���t9вS ��Ro�c�I-�_��=>����x!)�Ja_��q61xR��Ë�Tu-�q�ԝ�Ef�?6��J�X�����(�Z����k6];Y�2��e�b]�˿�]��+�V�:=���qI���E��xW�dÿ��7�ٱ��|�*�ѧ�
���}����x���Q�mVy_6��r���KB�N���Z'�A�v�x�,�KAH��;y�����������w��Y��Ydg��|��5�4�V�����&}��g>���h���5[��jwS�l�6)$�K숒8D�����;׵�����-���=K}�����'̤+f���65�Z�3��L9��,5��H�v)%y)5(��^+v�pNE���<mQ]^0��8���7}���$�
�K���6�R�0̤�謳�L/(פm�P|Y�^��0����o��i@�v�Z��vt���1������=(nTD��V��l��tخkI����U޻���-]~�n��aE@�h��n-�dy ��B$�g��m)S�=3�~9�T�	����H��;e�u[��7����`rKt�����k^�B�W���l�Đ$foW
N/�11CF��Ѷ�PZ�{�r^Y�p8����&c�|VUxE�����u�eXH=(b$�1\�j����Wl�
��P'�-4ﳒvﳣ_�y�l)Fe��/ KXB�G� �ɳQ���`��xPyhj��o��R0����~tM�?�8�j�y�Ɇd��"�?�L�_2�eq���@��X��!x�9i�n�����0q�uU2�w���:�~ �cgZ($7��xۀ�P�O8H�j���d��r/GK����������^���&�`�����.ԣ���@Z��V�̜�����(�D���ҮHO
��/TD�.u��CcC��zΜ��K���[vUGO��a��.$��0K{��q����0'���GؗX��Q׾���;��k�n�*�g��\�b��+��be�̤�o���,r���?g�����@�Ǟ)���\�b�tR�_$c�)�_�0����X����0~�
4�'U*7V���bJt�M3�b��WT5��u�ý;)��~��{�v�[�.%T�b�Dx��%B�X�^D0l�e�ɂL���W��OE��4���g(o2�+a&����֝f��3�Ҋ��!��O��y<=���y!,�8�8(�	�ӯ��MQ�v�)��w������&���yP�D�oQ<3�؝�V-���%�d��lS�a6�5+\���C�=SWdi�n+�n{����SF{�MW5����tb_��:Z"svf!mp��,�w� ��_ɠ����3 ,g�_Kq�]����\�"g9lo��n�`�:��_�s`��!^�P�p2���O�,�W�N���%j�������v�&�"���Yʥx6�Q,i$�fCW\m7/=E ����<g�n����e�FChq�}��|�d�~ � y'jd�w ׍�Bk��Y���v�{c��&�4�BC(�8���	�Rv����P��|O7�7��bו���+S (��C緧�N"�r��x�0�M���'73I/7���&�����dkaU�3�;��*�~�X"�$g|�5Azە���=��ȃ�Ay%S0Έt}��T�C�����p(����j$kFd���D�ݛ� s7��"
X�okӤ��%,DN��.3����Ǥ	�T-/Jz�b�ȼ��x�zI	��+�=Bx�T_���蓈�i�C���j���̢����)2Xɼ�ϗ��ڥqG�h��if!��x|&U�鋣��IQ�\ ����q!��LJ�?Ë`��5p�u,⓬����� �К�.f��C�&����N��Nucӎ�K-�}�����lp�YNkF\�[��Ö����Y��U2۔��8 bwR5��q?�ר��!�u_1.tcm�m��7��_�&�W�ui�p|��5;~�����������*���C���(t6F�ٶ�xnr"|[<�+�xx���~�ϵ�)��PB�X�f�s�]ɨR��� ߶Pi�߲� �	��L�e=Вy�����j$�D��C46zbƩ6�E�}	!a�zc6�&�t]��K��Q80r�؜�2?�w!퐍Q��Dk|C�w������B��^�H�w}*+u�g&{J���y�][Dц����T�-����p��j]Z��O�, �ej^���a�4s������XW� ��`rۦso����ϕ��ǹ=�07���VfnH�;R�Pˋ����K�b��_��;� N�!�|�L��4������0�w�|�-$2�����"U�C5|��6/p!z:�s�j�H�$Z��kaQ�^1VP�1��Ё'�}���߈���X��y�Ǫ�2p�q�#��rU#����Fi������td�[�s�uS;�@�`h�S��҅�=���g9f���8��Xr���ʜJ�X!2l�!u���t�G�q,��	��o`b����	_%܈�!��� ߊ��_�\��|d�|���"�2OI-�j���/�V�j��8n��T�C��L�ԌFhLp,~��0��Cߥ�k�[L�ok����w*��K!�5{M�o~w<c
�%%��6����U*��a	w닅��K���߾^���AhMD7����A�I_�
j�Ǉ�i�Y��P(n*���ga����洚d�z8�M�/S�R@W��vF8�[`{8>��:���T)�I���[G�0{�����`
u�k!Z�p���&���$���P�%r� ����A�L��.:w<�=8Q+Ś#v`'mV���5�uǅ�A­V �tJ��?]]�<�D�K�s��	ڽ柃u�0ޯ�:/s�L$�H�.��ik���ݕ%z8Џث���*!�Ŧ��YQ��yn��� <�C��݀TiN�h6��5a-� ~��Zw*�^���X��U��x�hi��q�:���1�e߸J�{3���� ֢p�o���U#^Z�d[�)&��n~���x�J��>���
Q�:�(b.��N���6���}�����p��t5F^s�olr��ba����Mc�]DD�R�(��%M
��Eށ�X���9è�s�������΀� a�úR?\������+��k�	�Sy�� ��OHaLAL�~�L���0�ÛY��� �6M�&G˵nӻXѺ�g�D�%��]�(4!��l?ia	��P���~~���n_ƶ��	�
3�f�1���=�z�ߦˆX�0g!·��k�S��]Ӗr�P��E}����P�F�E`���	�r�bs>�%����q��	3}^�$�*������^)e���KƜ\q��*�1/膫��*w��<�Y�S�6����9�f���]dzY���]���擈Fkcl�̥s����� [ k�r�N��D�]A1��,��h�F�]��Z/�YwY}��r_�1o�>�b�)8Q��f��./�������̛� �M����s�R�-�X1�*��=����2��y��>4��7��_s��S������-D:��n�ץ�s���$��=o��)2��x��F_�+�c�L.��I$i_�5�;Q̎��0 �� ��/��d|{�sס,&��(ͷ������7/Y��F#s��Կ.{7�1[n�ʚ�j3OG�Ԉ�z�"�����[Ɵ$���|��4���rR^�_HjԍKü�:���ؒ
F�5W���2�+��٣vd����N���:aoqWY�}���$L�	t�#���ħ��0�Bjy��5S�L[�cʼ��˟B������Z�Z:ay@�x-E��>8�Q]���4��`��f@l��6K����VǶ�E\���̰�Bd|d�(�0 ~1�U�i@`{�������XN�����:�E9ft����SY�³v��!��|�,x\������tRUEiU���F��"���m���]jM[}�ҭ�_õ-�`st��Z���)��zn�z�0�b��ړp���I�7�R0��k�G�����,LM�Wx��u�SCd*&�<���]�۝`K���a�5����v=S���i0w�Y>D(U��54��H�^�e�@�f�;���d3�߼��h��eB��[���$i��R�%��!`���h	iB��[�P�4��e푰fsy����h�c~8����M�5�(�����Ѭ숻��D�Z�ۨ�!�λ7�}��t����8iH碥ZOł61���G��iG��1dB����qD��d�eż�_��ă��~t�G���A��/�q�$�����'���8|>疋�� �Z��A
��O�>o��#�:�Kenf�@�^@kGS����ܒ̃x��4����:���|�J�X�qKPI4ě"�W���AQ�m	�䆬�+��/_��@����_��F(_ń�y©��� {�"ە���>:��u�g7B���\MTl�S�}?�������_F��E��@��Y����ϭ�yb'��W"�	�o��u{M]��~�E?Y�X��A�n)�k��\nN��K�/=0W������	s}���l!]+1F�&!�R����n����y��7k�� ]��n�a#�=�����/ 3�6y'�}����.���W
*I�vk�̎2+�n�`n7O-7a-���Ѧ��������qu!��Y��A	p��2�t�F�Δ��G�@��,��ĩ@!�آ�O���?�� �����5�?�+4��@V"�jd#�D=��⾮��-�!��dgڀ��s_̴�}�ѿ�ۦl�,#4l��RL� da��
�e$�I���e9_yb�˩ۀ��%���H�1^W��~D,�qw�9ͤ�s�һ>u����YKIg"�ߟ ֢��C���ߡ$����:Z۳���oN��kTo`'�O6T������B�+O��u���
���{:ϫ��o?е��'��=��&w�]�<p�����V���x}g�Y����s_��Z��;�`�+gJP��ju�|�3'H��ߝp��x��H�ۍC�6�y�omc�]K4��mY�eXqF�E����X3���U�h�z�}ω�!�� R����Qc�Mo	�P|��?�(��Àڰ��'�ߝ#P�]�R���*\�V��d�\:n\�T���0�z#˨GntZm�:dU���\���������i�I\R��u�g`6s?�c��G
��nu��S�SW�?/�ζ��-+8�ɐ�A�U�+����|>C��ˊ�JK��� EP9i�ܺ��&�tD B�2�ɫ�@����X�4�lf�%������6�/D�@&�/�������._��T�.g �T��+�ʃ�x�:��~��L��Ec[o�>����{���a
�����]��N���jb�񄜨dJ/�)���b�^u�6��и#���15&^V��MGH!��V���=�<���d'���vV;Y�����՞�/ۖ�&��g��񘳟JP ^}o�Eʎ�%X�e�����/���E;��� *��h�*lE/�>�D�^�i�;Ak��Ϩ���c��=񖤢��s�Z�O�Cj��h$j�w:^�A=��]�ST�+ʎ~ ��A�G�x��Mj��C��̾g��̹�7��zL(��-�\�W!����KA��^	�������-���)�3,����|_+a��H�~Y���2*nń�
��M�'�݃��4:`�ROr3������&����P(�
r��d9g�'�l��{Q�S2n���R�t���2S��I�d![��Yj�w�_MV���*~W�����YyS��y�k�p>+�ܶM-"�;bع�$��p�98!��}~+��t�7Z�w�ٳ.X�x��g��F�Z:'�Nqt]���Z`v̻�4|�d��r���2n�)ڥlk@|DG�MV�L�5���~+W_u&,8��c������-ӷ�h@�/x$b����.��>9�� H�I���?c����7k	k�"UOE�<���x���jr|z;~c�O��oiul�7:��x�/�7���`QGH��ހr�d^�m�,�T�JJj��Jһ��7�,m���WJ�]�Km5l�^���7�9��&�n�ЌzK ���������~��j�(�_�)�|<^U��� f�\���
�
·�g���2�w"뫟�m��ͭ'/+V����;mф������(�,~�Xm�9�	�~ۋ��]��/9I���0(y�[���}�����y��sݭ2JTO�i�OL��"�w��*�����e�m����l�V2���F�RmN�/-�`�u4���4��5�r�؀�D�8�8G����踏O��Y�v���a�S�g�[]i ��J8փ�������OD��\��W���V�(˱b���J�����# �c�yGu}wD�Qߠ�R�OB�/��_C��d�h+|��΀Ɠ:.!�}Q�ٺ�9���
�pa�Z��?�nU��w?�i���NU��)|�D�_�i������ӨB_w����=p��J�\�kx�T�PFs[*��1��ZX�,_��[K����	�q�m�<���\�AF%���$Ƽ�rv-Ы��ⅷ��q�d�6R�a�6���4hց��OCMEL6�iB�'�ɨ'�_���o$l��y�(]��-7(!�E���4{��k�M#!�i��Xf���*?�ޝyt�Uҭ��}#�#�M��% �C}�J0�H�G��I3�V�ĸ����3����I=�:$�	�b�0�F��3�����o*R��A���#�?A�5Cc���p�򛑙�h�LD�j�2jn��?@��/��Y�)
s�E+ӍD��q���݁�ze��-Xgt�q�����U|�B
�Zvu`:W�� 4�x,b��+��uF��e3�1KF�i�E��T��=Z5��ږ=�l��')g�;{��t.�V"$�:!�p��0(X�����%�Q��J&�K5��[?й/L��Pg�u�7AC/ؓ��D�Jm�7z�[��ʥ�F�����7F&�A�9��K�K�7�n��ۋ�}s��n��,��`�l�@WY�AJ���F0C��,$M�U�ﴕ���D.*���-@#�ȋ?z3Z���Ea՚v<$���J�/��]���hX�ل��;Yzwb��slA�g,-��aq"��u����%B��Y9��z�(��m��ؘ�v�\�7 �Iֹ�����@̼����CV��u�I���HőFTZ���b���l7u��Qڇ�W lԤ��[H�K��wmV���$\�XBi�v4�6~��}yJ�� K"���2=b!z���;+��������&�q��1;++3��+-Z���2�u��Q8��,��?�ۧ7���N��+%�P���2����R�q*-	S�G(f@�m����Co3m��0��J=z�1}���0��/���MRv]q�^��Af{��-H׿A�Py8��b.� �+�-S������yj�$	��^���b��e��10��(Y%�mnفZ�Id���}��Bo��ǵ�3ChB��rr~��<9��7�9��a�`�1�vΆnjV\��D!�5�a����B�� ����IE��0��DZ5��0�#G.�0+�����L�����%�z���<�=r���Z�V)��PL�qXkڻ3�/S�r�@�v��yN@c˷(��e�	'�Ji
ڨ-*f��4�m]MM7�����6<
Ph�O�����G��c�B;���7�(�ឍ�=�7)�7�yBޯ6ۮ'�Vu`�"u:"E0#��v�ƉǢ��Y+)�̥�v���RU�/�R���b	��B8���S�ؠ�d}``R5frL���1`��{.���WO8�LL/.ٝͯc����$��)A@�rd�"� ���?|~��6�A���# �%�)���Y����D{:�E�ۜ��;���n;Wm;��T�O�5s�<�\Lf��WJ�H���d��{@%T��u���l����.��:�a��^�bQpA����T�WH�P"5z{�I����`���� NT�z�>pCu��E7�v�|�\���ֲ��>9��δ��[x��
���Ku�-6@X�~k@����W����#3��tEC�d��_NfN2D�D}�(r_�����[� �<���o��a��t���PhM�b��2�ԏ�������*�����Κ�#�[k�+Ny�֖�_�K���|�C}~�a�V�m�xhk�g���!m¡��M�*H����wȦM�Z����j��5B�hD�uR��]w�f}��s�9��t���m�G��Ǫ�4fA���Ʊ�K�X2�y��
�F�ٟ��&~���Y?My�,25X�)�UJYW�4�r�3�l	^��r��]����t%��,s�s�;�4���D��$�{�x0�rg�>��I��5Hql��0֛Ɂ�(��+�,3,�����S�>Hบ�a���uC���=ߏ^�_t\�P�5���R����i 7�d����k@����F�ғT���o�\C�?��ᙗ��1�]ɡؒ�N��uoE:��ʷOU_8`��o�B{/a%��ˢ���hj�i�Go�<h���&�T���v-kn��g�r�&�@%�?�ev
��ǧ�嚈��E$X��yK�e\���a�{º5�m>eLKq��k�SZ��|�Ԛ�����b���ˇ��Eٟ��pT��m�NO��|�EoX'P�?#�W�z�?t|�8ie��HU_��˼����n��#��
4yG�L��n����O��E,h�*,�5m��El�K�~m��Ve2�W��E[߈��lk{�:���j�5������||\a:+�@���y.w�-�Ձ�_���d{�`�\�I �*�4�13�N_O�%�X�H��� ��e��K��)���q�H��'��>A�A]b���[�w��R6p8X�A)��s���[h$��y���R���k�Ǭ@�Ct�76�0��(�c=vZ��i��MA�(�	`���\ 6uH�P�Z�
I�i%��q��7+r�=t�P�ƐԠPc�Wˀx�!Ǉ���m��i�d��������ʅ�Ӝ>��%����ۜ�[bt�G*8���=K������oR={g9�%$������`#J���x���ƿ���Hm�_\�h����0�I�޷�����y˷M���PP뷺0,��sR�	Z�K�P��Da�K���Ȯ�A���]� �O�\���^!	8wg��1Q+�kh�0�pE��Q�E��O�f����Ұ0�K�d����9(�=��A8���䩢�LH/˛��y�Xh��QM7m�h
�����9���'�E��I/f "��Y�{�t�=NM����n�	 �������+��U��HD�m|��U�_ �8PM�	�*���ZQ�� .O�Ff��4����K�T-��MN��+�pw������V]�Ư���a�q$��:?�b�Dԅ�Sŧ����������	-`s̢=n��Եu�*��EM� �M�U�pE!�Lvh�a��"̗:վ\r9�q	N�L?SȖ.����xiPN��g �;:l�l{�L��-2Ȣ��a�a��ʐ��d�0��N�^]&�^�S��`��4V孺�j���Äo��7��h82,���d��0�G>$V)�����*�M	�y^��}Gz�m3q��6�O�.Ī@���`d��4���m�r�ݭ�z�~�7	�p�E��;jZ����s�������S_J���V��
���)L0>�]Z���r�:nI��u�=Y�%�I˙f��{�&o��X bs��������n	�)�Lɦ�/��T����$/����?BF�����1m�flT��ܘ!ͣ=�/D�M�X��\e>m�5'��u`���R��<V,Xκ�y�����6���Yԇl�׷F�bb�/*�т)�%����Ws�fmҏ�88?���w�v)�����-�{��m�b,����P��/s�R~�Þt�Y�#��U��Uf���b=�R1?�4�k��p�A�d�"x�5Sd��J�����PwӢ������/Ƨ�c���R[od��r|���E����^hrK�,հ�qӐ�	V�ҐOU�jl���Y
�.cS���|wA79( ə4g��v�n������rCUEZ�g�G�N�V�;��n8�)�ʐ��n:�7	k?/S����φ F$\���s2Uz��[���LQ
rt�%��v!v�bR/ҍX���>�˦���������
_��J�>�P�d�o�G�-�?&���%�7�d@�W�8��c&_`f�|��'��x�?��j��V�Q$���cra��B�j�g���c:��W�TD�sxM�6K���s�Fw\%,���pǄ_t֑H�ߥ��K�1\�=�T�����' 6���a!*n��+���yV37ey�٣2�$�PW�V��8!.�[d*�I��<J�B��=�my�c�p���*��vC邎3(e=0\�j���pҦ�4��V5_�S��Jg��JF�C����t3'u8��^i�+�s�h��R�Y��L	�уDhz�,��[�<�T�~��	����"d���Y 
���3Q��=�é{�����F��}=Mn��B�Q���P;G2}&��8~ \x�6k�.T����7B	���"��Z����Gn�wbѓ,� ��<ð[��}>@���ϋ�*�����O����9�X��3x�Jd&�����7-��:����8����E��#K�8)��j�Q�T3�}@���3�i�ק�M����`�����vS�|x�~;��]A�Cf�F��:�0�������\v�u��Ƴ}���������PeB���- ���8��)���t�����?;�*G'L~��CH���H�\�=؍�@aܷ��J$;̖�Y�Mk��T*�{.���\0�Y6�A�d�c'���I�l���r2ti�ǬC��+�P��4��I���y�l�ڤ*ۖM}f������T;`g������$*=���沖�+9����QG<m�ڹkw��Ơu]F��@X��4���Y��!҃��}����?"	���-@�jqE�/dY���$c�d)�2Y �ߖ�C����q���R�O����:WV^��~�J{:�q�b�J&v(�P���5YП��.�V��+��S�G��哳N��\y�"��͋�Ɓ��at��T^���.��9|���q_�nb4�b.,������x`@9d�^Pպpl�L�P���h��������f,�?;��w5�[�����5�)`щ��:#�<�s�.NTS�C[����,�S�U������:+|^��MQ�B�\�˼iSȋ����;�-����t�ѤA{�m���MգMW�D�������NE3�myܚnLl G�A��L�Wy�GePylC�< ��1Fg�0�b[���{� �V�?mm�jz�
�R��sN;�mȆ���٠�q�?�\�3�u��)E�!��EJD�a�D[�o�:���Hw��mÿ��� [�{�ձ�QU1J�{$f���\�-���6��V2$Dy/VXv�
�k^JU�nD�<�/>�|[�(��W��֩c�&��P��fMO:��E�[�}J�I6ؖL�'�6nM�[|���h�?$Z@�r7+��z�ЃVm�ZS��mF��ڂAQ?�����J�K�,	�+/y�=6��S�ŗ���,�4�O\{������!��],�tA�Ng��N����m0#�J������5)F9���k*������OdD�v[i͹���p�ez��/�~m�Zԫ(�Y/����M������U�d�ak��C
���r�����W���MVņ���r���;2}��|*�p_b=�b
$H=�\�Q)����<��2�Y�8iY�feUe ���u0��Q�@@{�1��p�޹W���Q�� X��Q�����xB��}��|��������p꣰S��+kL��w�����c9V��C������d
��6���Q����Y^�Y�PO�Mˀ��l��K1��*�