��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�����1�򸳉I�$�/�G�QQh��X7�y���x�]�C���}5=��g�)��k���:n�f�ɹ`��y���C^ڧ\������'JQ~!8���nh��F�E6Ħyc�B�~�x��Iɳ���O/�V�RP��B���ӆ��z������-3��^ڝ��Hv�������XT�d�w|P1�Y�H4�I9��zf�F�N�_���Лˍ֚kV�s�x/W��}�d6k����צ��up().�F��ŹB�iR�^�@�D|�k��_J�5�HCť��Iֲf�n�DwD\Y�c�1�<��@#Ŵo�L:ģ�N�^�80d���8�
�����c��tNL3D}e-�vt5��$�Tho����I��zy�bHt���n��6�"�6�w�)�L���Ğb�#w�LA��r��x���l�MF��^]�j�t1��C=U�a����D�� q��#I�>0���a �5O�8��8����э�^Mť���e�� h��3e\����g�I�㬱�w+�7�Eu���>�=���G��B��+��/�*N�,=
)i����P��n-�n�a��G���G�Mp�-ᾼSb3�;�}��C��S����~��������VO�E&w��j�'-�=g³J7�&��Ң��愑���X������А˭E����C�Y���y�vdPG�ƥ;�SA'�i�|�� 5+B��f�����{�d������Ɵ�2;CT�C�C}l�WbC�}��0F�3�����+3�y�A3<�eΗ�4V�D�^Y�m G����(4ŋ�hy��W}�x;e%lS�N��*�p~`Pz1�pu;V��gj莐2_���v�L��m.ݑ�aX#t��%�F��w@�l0��D�(4:�ʸ���a��"Jl��V^��	���l?^*b5�Zh��n��u��gݟ�y
:��ڎ�k��}L�xc���We�>�:%�3t�a�5|�!u+e����-�3�* �,�Ӽ��+؍7�����6��9�e�1��C|��R�!�q�[r<!�;	�G��E����GXٰ���`��.��
!�w~��̄PFS8T8����R[��u4{��`䤥���{2�'%��LN�@{�����LP��K$a�¥^�=��e３!P)}0�p�2��O%�ؗ�T���F5�$��rH���Y�~ު�f�mA�>5}n
(Į��5�BDn����U�^�,d&V�&K��S�-�������7mL%�\"Dz	`�q�=�c��0�S�� Q�ڶ�%G�8��Th�W������N�F�;�J��Z����?M�P�g���ܤj�u.�P�vhxX&�w�#Y�;Љv�[�Y�;a�����D;�G�[��B�rw���dV$˔�p����͋�<!V
�y�>X�j i���A����f�������I#��\�qC6�6����q�_2r�/܎^������k�+O/�n�~����)@�j����,\�M5��������R�N80gtL���آ�Xye���F{��;0�8��U��{����[2G �{���2�YĪ�|&4�a� ����dF���A��i����lЇ����A$��b�E��y^�e��g��@�zv�"qc�"W�X����5i��V&�Yz��۲*�U!0Un>%C�:��9�B��\�a�gFԥ^���OvRK�wCT�x0-�y��78]oo�C�ƾ���R]8$���h�;Td��Ԇ����[3pG��z��,,j��<�	�WCP��b��AH5�S��=X�%�_<?��l�C
�����9(y�~:�Z��2ћ<CIyhaF�[�zu4��������0�Z�%�jr)8M��c�}*I�$���O.+I�? PdB��g�����$�����S�.Ek+�ƀ���O\e���'\g���ѵ1�ZQjX�G�:�wS r �1.B^�d�8._6G�U'�q����/Z��rk�V�A)��[t�B� �S�D7-c�)i��c����O�o*��D�������:��N!��5�,��Y�����h��F�$�&��Xy�E��,���&�[ǡ_q�uE<�,�g�?�:(��Hh<�U�1w��p�J���m~��ګ����D��j轕C�;��-Z,�xB��'<iQ��+��6��c�v3n�����; $�2vmu;k���-[ �U��̨K$�����YS��CX�p����8��P6&���f�A�eN�E�K�1��O"�>����A����TN��g5����)�wP�T%*��l��YIh�"yj��#�y�~��{X�3�آ���c�e�{�nC�"��e�7���i/B���V�DD	�}����re���Ιf>B	?k`�ҋ��	0�D�70	uS_����S���ȸ����%�F�x!�r�Z��<ncy���������5��������ǟ��m7��6�9�� �ANs�ns�*��C|���	_.ڑYz�`��1D*0���B���ɭ^C������C�eJ������}�� p��iz;fZUM���a�DT����Px����-��-B���l*g6�u�p�a�N�y�:^���镟���ձ�G)1ܬ7�Ѹ~���~�N�\9��ȗ?+��gS3��x��Y�hG+�w+6a�|#�L�'n��}ݐ������w�� PM��?ȹl���[����6�Y���%\J��9�C�G[�k�=�@ �릒�d
�q'ސFS��$����2yi���C�s�P����B���v��� ��!��-儅��wh4&�w9-i-����V����I��2��0o�_Zj`�n�d�]G�(�JlQ^`Wi����[#�,�9�+��D�� dʹ�1�1��`�;HX}����[��G��=<�;��`�S�P`�@t�_���!�#�)a��`��zïV�?����z�G�6*�,�[~T�mm:`TF�[kڶ�*=���T��fϿ8` t�m@��[c�"�[�
&�q�@�A���iN��2a^D���l[ l����.�X�Ġ��I���9������:*��co�*�,��%M������u�p��8 M�c��^w���[��$�f��Ao|�#�8��e��b V=ꯕ�#�5C��v�B����m���z�<WR���	�����ă��<���K;	v����t���\�vm,���"�7���b��Q��6,v�_U��t�_�z�+�g���`M$��z�Z�}�R5Ka-��O�@�]�CVJ�J�lG_%jDbý�� Dx�5��s�5�x�8|&�dmW�*����֏v|���Vc`Cw8b���gĜzԸ�#_�m�J�n�D�6=ܢ�,���V�;r��Д`� 䞁J�)�^�� �<Y����a|
�"ݣ�
��:\�=DH"�H�)��'rxe�>�
[�R(0|�w�eĸvM=������bcw�{�7�1�c�D���
H����$�� ��	{*�;�o_-,,�!�m��=9wlL�b��ʰ�T��ث2��E��a��h�����������vq9E���fʣ}U"߬����%Z\�'
�e�}D��d}
j�C��W5'9�u���5ܡ�w���54P�=$\�VJ���D#u7�k�"U�.lG�<ӗ�m�H
����V*� ;^��#krNg�����y��[)�B͌�$�W�`��(�N�b�cBT������� �̗`1�M@�rh������G���)�`�G�B��ق%b���V��?���[ё��>�gh9�T+e4�t�S����B�H�����߉�ﰥ���&6։Ǡ_��VE(\)�҃�Y����L�����e��a����oJ"I���y�(�rΌ$�vz�v%�J|����'��)[���6]��0�̃�K�4��.��d�����;X�E-�����/��W'OD@u%����Y49�_��׹����щA��W�o@X>�̧t�L{�J�����Q�`���{Q���7�b�dJy�M�[��ʙ�_NԼ�L�m��K-�4*��_n�!��	k{��y�� ު�}��zG��T�9���Iz��ӧ���.�.�fZ��?��.�r���t�W�dĵ ��Q>�ɰ���C�j�h�M@���n�9ŰrU�%��v>,���܂�#�g�ý��Nh�'F�$�d)MP���;�C<�	X���3`�f^M@D(�H�r"��T�t�WhU��x�l}2� �e:�Bݔ�4��,��{T�E_��N	M	&�,�#;?�lV�����B|[��#� �t $A�ގ��;�E(�&�oX�]��_GV5��sl�bF��뜿|��^l�	�/th��c�X��-S�H��؝E��.���D��}���s0f��!1����o^�4���0&��;�(tbR�~2������ ��Df�z�e*���J�&�^�G�p��ݿ�	�l�M��WL��Ȏ����d�d���hPw���\�Z.�w7�G4�1����Q���
�*���Ph��s	V����W%�Ig��"ڢ:c��"�d�"��
��~�yA��=�� c���3�p�l4���K�l��� V�a��EA��sn�i_^k�PI���t�٠s����΢C�c�zב��	�4����XLqq�t���z�M����g�tz�Ea�3XٟZ٪L�a��p�n�0�i� �^���!2=�S��A��V%C\yt@J�J�G�}�OrG.&���f��9ts!��,��0�~�ټ5�D"�����x�R�{��[�~�({��(����nP���:%�Wq��&m8"7����9��c~�Dag��y Q�f���G�6�)�aKp�ׁ�l�\M�D�KĞe���Jv��$q��,hV��A#����@�'�WABM���4���>p{n%��w U;T/�HH�;��-Ṍ������2�g�0���Kqb�P�C�6��3\�����hͅ+L�ه���v犝�:*��.�>F�����4Q��WG���`�j6�C%�r�h�5�a�v#�
a[��X��ƫ�R�}?7 �:GL'�o��#&e��b��9R�rRL�*�0��$L��l�1L[�������}���F}�QG�2U$���`�~���"�Ў?��sG��Q�ꔣ�ɟ�ۻ��I�ƻ^��w+��Nk�*�S�'�����r�L�%Z���=�c8�Uz��&"��χ�q�ʫ��z��*��L�l>e#JV���S����k��2��U�_�iR�EE�'z�5�"���=�',��Ƒ��;�G	�M<�o�&����y�6��Y��\$$|����H�ឋ�#P�#��=���?�G�g��$�4n���C��ٍ�˘���	k���1J���u�'GIÐ(�O}+K���*����	#�!�L��i[oun�qEV�&�Y.Z}G�+�����q�\ܱרif)����dg����Ҫ��WQ~|<��o����dϊ��|`�f�;C��?i<��FU���k�K63]H^'h�g[��b���m�Zb�S�N<��Xc4#�0p
n�g�$����d�K�(t��499�����Wxl���y������,ښ��(]O�Os�7����1J�ێ+�J�L����=�LH~�Wrn���.>���}��4�;1�j)��bt<��~�$>+��Uq8��'!�$���F@^�Q�tcUF}����3N{F��<d!#
˃����߀T_�l�|��+����}P7�Arq�O��3{'e��AEkk{" Hc� ��E����w�O�-EJ�*5�E~�Ť��7)j��Q�;|Āu���7Q�g���ΦІ �M�O�7����r�Q���3�MW��KG��y�y8�W|��o��F�6� Ij�V��&�z��uࢻ��4�S7�c����?��1R���D����8��{���zG=��]e
���4V�/	�����%Ȣ��2��M\8}�^���5����+�z�����$(�����	N�I�vBZ���7���Q���z��@�����nLǮR�:��i16���c��srk�]q���M�gS��P9S�[rh�;�w$�T��N�H�6�\!�>���n���]��U��g�`z�)�j&$�?Rٛ����t����T�'�,3֬�߰K3��|����N
��Xi�WV���[�,���n�֖a������Rk��?�Z�m����X���	����-���8���}��3�}���0b�
K�
�<Ȧx_�I�
j!��>}���d�J�Qs�N��_�攓&D%.+"	�9�O�fdӳ�YB)���Lew+�`���{�8HWH����sȬG��\E=�ȝCw%jN	���O⌤�Z:�6���I�=B�`�H8E6�s�9�F�Ӌ�s(	�r�O\�5�B��W���2�p�'�W�rgw1d5'=�fs��s�'���s7� @jdr�q"��[���vl�"�+d7�H|t)0O�_�|_f�M�� �G�A~�yE>Y�j	�`��(���3 :^��z���_N��`=��J��.8��軘���
#�&�]�,���O�x���gQhQ.-j�@U3Zx}�@�ƙ�-���T����Y�D�|=��O�d�P�fQ,�Aހ>kn9ڰ�C����O&�@$0��W&�-SW!P\JW�ʥw$խ܏�ҋ��\�����ޛ�1<�I��,�>�!'19q���c���יB���rB��#U
v&պ�#�!+̍�{y�U��\,��d�w1-�x���*�w[�2��k3���:���h��i�� �1��v������'[Ƿ�Á�߂�lw�V	��x)��o.�����o�O�rC;ޏ�nu~�t�Mn�Lf�iw��N��i^5 ܧ:&����om7�J"4��&������\6�ɗ'�S�Fȉe�_���0�������f@�\;�G�6�?�<0A��5�����d���ȟ�`���*��,��׍=�4��Vޘ�]{�Cu=��Wp<�� j_gf,�x7��J�˩WH���g��(��]xz�^�BL3�ӻg����%�3�vVm�dX�Ř����~�m�&|�M)�mM ���]W�,���`+wή��'�?y��d�SЭ쉑�.Z<�/��:ֱ	�[�<Z|���f�C�$_r�-�.'Qд����Ŧ�w����F�O�����Ud꿂�=g<0�� �R��IY��è?�e_i_�*�ҁ�8�m���L$42�q}b%˨�ܟd&���"��C���~&+��H~��=�N��C���
ɚ�;��#rO�7S�ܭ�Gn$F��V�=w�$jրE���2Ԭ���Y�)�Hw(O�u�C��.��?�,�Y�PR��Z�[g�T�Z:@|8x�^��y�����@�:���aA�(_g3&UQ��q>��B��0�)��OL�S�Ғ�������;�1����qw�5�`a��Q)9[�(sB��g�ܠg▞U�Ú�<��_��x]�5����qu.�%9�T�d�M�U�iNQ,�ó�Q`�i��P��`{�sP��Dh��12���s�1e\�Y/�Z��8��bZ��:X-Б�����@5��]t-�)�Y�6e(�HS�&����ߨ����-���#O�\�N��2^YTD���M)aRd��Mͬ�Ic��b:���1�u[v�D��	\Ni�N�Y�<���O���P�����}�e$\+�7OodEdx�+Y�4��5��èZ��~i/^��:R���k��<�Ǿ�/�-�1)::���|�6qԩ���?+�`AQ���jG�Y������xH����U»D&���o6�W1|D)n����W��y.hy�l���3���&����x?ɗ�f�@%�/���*���`��Q�e���:�!/�hծ�р��������?G��]�Z��8{�6�����Kp���{q>~���^�O+���#�¬8�HڡAn(�4$�O��k��[ܷ]KkPFd�_�X<J�.V�'M���4\���דH�\�(� �S���'�:���FZ(�6&��_%�WN�ĸ�v���
�8�	U�/���t}r*��t{��й\8E��;�Ҙ�d�
X�q�~���Sh�\�y��Čf�q5 ��BS>F�y1�7�[�L���m�����/�� ��X��KS���l��[��QL@܀a�8}��;BZ��3+"�X
�x?����QWu�68�\�VǗ��[�M���T��0��o0��/�?�̧П���G<D53cORl���_�9��9N�b�Y�^!�`�~��h���ĺ��~���\#I�y�ǭVA�Bŭ�g."�`�����҂s�~
Pl�jG�&8�Jk/vpV	O��J!AQ&nA�#�������t��l�X餅��m�j��t˱2־������Vx;�}��\	�F�m8�����6��n�O���V�c����b$~�nY0P��N��/ �E���̈���E�j,Do�m~5ʹ=�F_����l�F�А���6��f� �S'@(�I��,Y��������Zփ�ŢZOvCe��%D1|�����)[^����Nt+�_a��s���&�Y��l�S�E{Q�&���o�&��kE�o�*�D�q�x�2|��!f>QH�� �]s������;�n���"תW�N�ՙ����0D5�措��.s5s� �'��9X��y0T�L|_I<�HWq�i�����|Yq|[ic�^<&�p�C������˿c�^�qh�Zł�n��l8���i�|�n` 3e�fI�>#�3��>k�|���˳�$�.ت����M�S��T��"1��I�U�DjLhe���H�G_�^h�"�.��h���b�xa���'�Tt��)4���U6��Ut�J5��آ��� nx~��w&�	3?!m�g���_��#�IY֘nˇ۳	Uǖۏ!K=� ��2�R��xL�&	v�����E�#M���īY�M�����?vU�%)�WcYza�^9_�xR��K��7�S&O�u
E�j�3i�^�x_��S7�S_Xt;�J¾Z�R�����<��BNiO�߂��bqm�yE�G?®KC�-��8��U�AJN�F?��K�_��H���A-��M��
5&>�&�K���)�).4,���|..*bN�p�I�0�?F����RF��>��?�{�Jk�V0��]!��o��J��6�6�*�y�YH��B$<uU9d�HZ~d��[#
`�YS#��y�j�<�<��9l��?#6��J7o������u�`�(�6J�M��`��>��>�����̡'b0qP�=��:�ws;�x╰��Hh� ��Ь4yiUP��	�2���-&W r�e��n��Qs-0��<xa�!������X�� ���K�@�a��>s,����ʍCO��A�����M��n�P��L|rF�bw���I�)�7�E	��gZ�
V���(s��+`-9C!��M��a?Z}:cg�)_���̀'?�4�lT�*���O7��ò�y�a�~�{"w�=,	��vZ�K��i����a��P��˙K
#��M�X�8N��X�46�Nm�|��M�C���$\VHG�zd�x<�L�w�tC ���&e��qKs��Eu�ļ�7I�u���*չ�c����n��&I�� ݑ~�8� Y�M�m1���\�s�8ro&�>S���VE�i�4t�c�r�,���w�:5B���-�ݨ���Kr�y�R��0�m:m��o�.�Or��I{ƈ���.�k�L53%@sO�5qW���������Sص���.U�`>=����B��;����)d���T�F��r����ɫkh�
������$�y�C������i��6͑T�!f�n�x�`J����z^v��3�,�z�*�%j���H�b)hx=������q�8���Ct�I��8�5~LkO&�2VI���S�U Ym���.�$oP�y�|Ϊ�Ag'K�98p�åVQ�;�t|a��F����N3����a��1�ߏ��IHK�̀����A_�����e�U]���Rmf�8�J�/v(빳����ŀwצ=�f���JB�<��_&{�b��c.JU��j���*���zx��e"V��q�ب�~���+�(k6*�����]�U�X�y���ɧ�[�R�P�����,,z@|ͽ�2�Q�7$�:�3F��ʡ�L4	:���Mg�
R`� 9�F��I�E�����<�p! Ae٧ą��4.�o�x�2�c᫺�[&f����9Q���O��Kc����.[���Z��3"�|\\G��<bֈ����{�[�Fz��oI�u��|��FđRcu��ם���(D�]j;öV����'_��v��a؃�]C`2�̻�2�_Ԡ���~u�dcF���pO��$\�,T���I��i��xqRn��4֪mqVёҼŶ6�xAx���]�H6U�KvJ���^���\�ޥ	w���͒��%|�N}j����zo��X�[qHc�)> �Z,WoL��9!R��p����j�XT�&@�B�����x8����ʪ�%Op�%h�>kJ\��1�hJ������^��
��Z������(��������� ��p���O����n��uu&gE!b���֒�?���u!�.���B%>���i|Ch��,�-
�t���<d����6D���\z�1�N�q�������E���bM���P��D�����g�}=9���${j�*�?=M��#�����>\��^�!��P���a�Pd/��0�@^��ƹgnP��v�&���q��D����������Σ.���Y�Pa�~�޸/��pJ��T�'�E��
q���RAr"25��"s|�1�5�F���8��>/�;�wDT�j��<��Y�t�ݕ�D���q]�C�Y��7�gO��]�Y�AhMt�?�f�.�� l;mh�R��Q�0�>��q�@�\�<��'������(W�m��}bR��e(ѹ	F��J瑩ⱗ��;�P'	[�D֯9��I+�bi$?����۷���@֜;В��f�`�"e�]���!*��Q�
��BҔ��5eq5O��E�D��67H��n�nU�X�B����QcF�c��:���������ۙ参�5(f�k�.��2�9������tO���}2����C!��X,Xm��� ��	tC��Sb]Dv�Al�"�ʽ�|ز��Kw�v��7J�y��ʄ\�ƛp��y����[>�0��S@n�mҺ�*�P������;����6���͑�>�
��4���4���q�a7����UPǜ�;��U�%�0h��B��8i�q�̭�~0L��@�狤��?�L2>'�d��᠗�ʗ�
֑-3�|����X�Q�Z
��w��!+U��h`�{��S1��f��y�O�6O�b9��c�-a��k�ͫ��h���� ȴo*��n�z4�d�\�)���I�������̓�ۋ\ZU�M$������Y{r$qa0M�1�~���؝����l��`�C����z�YB؉<�=g��C�!��ʈgҞ���oj��T�x@b�����Z��D_�l���*s|KS�����_�uB�O"y���#ݫ�lg�H�.ҋ.��_�%�����נy.�K����j�B�	��t*»��֭�Ԙ�G�D��2���g��oчGߊ6���H��V�n� Z`&Y뱗�կs8���[�ϱwP+dP��yW0�岈H��)�چ�]~�k]�J�uE¾$2Oը���m3�%�g�C��
~ǀ�'m�Q6��i~�m�!�/��2H{l�R[W:K�P��F���Ou��}n��A}H�Q��@��dC�#!X�s�4�\Es	����8�G����Z�E��ȶH�T��9��ج	�en�u�ðExC�8�����W�[�A�z�E-C:7b�˨o\�=~��r9�};��3q� X���~��f2�S0�I����0i���e�N�(|��ع�С�8se�0�N��O�A��JV��Ȭ"YU�j�Z����b�����j{w�W�+{��Z��T�е8#��E[�g���_��z�:���`U�L*_j�P1s��Ћ*O��N��q���0�D�����؈ ���_����U��$f��C�b���H�]p.�]�@ێIͨ��q���O�pS��h��+q@rv>�
�����Z�[ĸ �$-���K�*pC���i��i�J��}�I��9�SAdE1ࠍ=��7���T��N���0�������D;r`��Iu;9F�y(��Hv�6�fR[�N�I�Ƕ�V�I��/� V�	W0��z��j����w���j�����Iɀ}}=#�Y�`�P����E �4�c�ɿ1o6Q�i�/��3	^Y�wR�R{諒f2���I�`}�6\�^$(61R�ok^�6JP�믅_A�W��|��ż	j�7\C��	A|��ܡ&}m��$_�N�O
1���wk�]DԒJG�'�%q�^�g�-c�8˩�U��YӰU+�Ѧ��9���w}��,�s��K9Q7���nǳ��!���[KJ�B>�Q,���o>��Rem������cD�0q�,q�A�����31p��C�ɨgB^R��ͦ��#�}�E8�eÊ�}a��$4�b2�����+��?�/N��N����K���*;�.�e���-%}6͙���'�r ���
�=B=����6��ŕ�B����I��.�%�k���B�T���9���d�J�2ۜ�U�d�jd�z iw����s)�ߌ%�����c��(���:G)��vd��7��-�=cȮ��c�r���?����jΔ�!g{��m����F�8�u�r�u��%�iR �aA)Lf�ŊE�
���T�Oy�6�Bü�ˡDA/�ni$�% <D�OÒ�P�z0c[����G.��D��$V�]u/��4Gn���o0�Qp�R'��_Z\ޚ�JO|QpEk�w1Z���m̓��C���������E���%��{�`�YW�9�=�w��Ǆ��%F�'���1��������+r��@�fEd�3��sP�|>�d�Ț�1��������+�,&of���x�S6�EL
[�
P��9�D.�Ã�;�� ��N�D�;�c��p��ج�+S?o_ݲ��/w�������s�ĩ4gWh�;+����.p�.�@*]m8_������7a�L�����2�(�Z���a���.׳��P�w��:L_�-ER6����������ɻN|Z�h��bCe�p��k���n/�,O_���)45���VE-Qet�1R𔤓�B��5�=`0�Y�5OY����:*a����9M2]Iȁch�K�z�.��J����2�7$M;A�1�syi:7���-��N�����p2#��њ!��<��aP��'I���������=�d�C�-bB�als�,�H=�0�_�ſЬ,�&��
������o��ý��4`
�d�V!��� ��%�o�x�)��aJ�G���DC�<��L�]s+�P�m�I�e�d%�̠c��� �����61�]f�e%b�l��U�~/Z�ש���\��o���8�[(�.�xП�%Uq)�ZG<Oz>���C�,.��/w�oJ9	�xA��;Q�Od�??��ݐ`��~�e��c�9�;�퇚���m9���2W��:�M
�$gć��$m�C�kt��Ҡ	�=�_vh>�֝ͣ7�Q�}!��g�������G�'��^�rD(�1�}��k S���Zh��-��I�q�Xh>
�E���.7��m&�j�U��S�DrdFʖ]ա8�L�1(|e��[61+n��j%!�
h�������>W�L��������12[�s����.d�@�lD�B�UP��H�R5ڀ�xԎ&EcƋ3*�6H~���[�Z���(c+�r)1�|j
�����
Kg=f��I��oa.�I���[���*O>�X�$�;��u܋
�E�=E
�O��	EB���6��7�	����k.z[[g�s�����N��������4��Q3]�OSȁXD~@|�k> Ś�>�zF�MWF�-m�Y��*ݝqCu��Y+J$�����rvo����V��~���:4}i u1*4,^v�G�8�wǾy�j ��$͖���׊#�,�0����y鈨2�ʪB���Q���P'x���ک�=�DOɗڹeeZKR7��K9{U���;��͐�<�]`iO�*��,�)1�/=�E�#�؊H�l�ST����"��bv��6�l�s��5��՟ZO)��!#:ג�3�h|�:Mc~ %�ɠ��!��^�y-X^���t'���+c�'��h����/��V��=�/�b�~��\���S�}���ES%蝱��|<�)sͮ^�+nU��}�ݟ�����A���l:�X��[�w� !���[H��E~��p�tr�D���)k-���o�70&��+?S(w[Qw���.��8j��u���ֱ���x*u�}����-_������$�z,Nb�+�
���+T���ш��D^��]�<?b�z8�*�}� p}y����2v<��hx}��ٽx+QK�/�P��_�JP 8��i��v
߻F�%���pB�޾��Q�k_B_�j#�R��W9��#fh������Y^&�BRt�ŗ
&V��$���͎��<�dϞ[��Tw����\�;�\�#�E׏m�!�R��Sb��}d�f~3U����֬��x�p��|��� �kS�`�r�aW��
����^i_`)�W9WK�x��~mJ�}��iD��G!ԡR� �//W��O�N�V��hnϏ�< �.��ֵ��'.j��4I���]�dځ��ktFV��ΰRU�Vm!و�rO{��Ir�I����y�m�H��/�&1B�94,5����g�<�QyS�C���� �P��w.O!�|�u��O�ꠜ�-=��{Ӣ���Ӈ0�]���T`gPl��Ey$��4-�U�x
O�hH 
��$�×@��@Ȉu3�2����Z���K�����A[�{	ӥ���"��
3(x��}���L��JxиU�yM\,�8�K%4��i��/w,#VA��eG��U�.�M�J�?l���r����3��JV7M1}�;w|���'k�y|�r荦��W���/��S�R��|��\ϻ��B�Pe�82���@_���椕i�#�!5;Ф�%�×o�
l��%��P�;Z�%�Tc��"Cp��!�J���Q�Y,X5���8�?��ʴ�	V�{�gQW6aj�j�Ы;�d濹��a5��Ԙ�b���D>��ɲ�ta����zr���������=�h��F�G�]�z�݉�U�_��FO��b����)8�?(;Z��oq�[>�ӕZ|MM靄�㏊H��bo�o�|�-����4�/1��`��^�>f/�l��ɋ5�pY��~|�ﭲ�.��.U�Hާ���1�����_Y��[������S3V��i����G��U�z.g�o�_s�+�=�Ns�g����>���U���XP�^Q�K� �١�< �E!�[e��y����M�г�c�r���ҮėnoRes{�-�e����h/�+�ajh)�E��z�[����� ������2��>�~��"ެ�s�^a.�ּ�QV`���AR3.����$�1<P|�6U��X4�'D����y�<�	��}����d�[+9��9��ھ�O�.5,�����b�1��S&����m�#)�qH'����k޼�J�IO�#�!�3�Fu�d�C�h<PW�Q��-\m�_.W�X}�ux��C�c�Y�Ҕ��=�?Z���;��Kz�%��J�v�MPD�/n��2D&q����� �-�w��?�~<�F�:����1��0�q8�?A���N(�@�j"���*�N��Ā-J���zvlT&4��� �ܑ�4A�-ؖ���53��
��ж^�����*~Ǯ��A8���,4�w���z�Xr&�=�a��QJ�905�Rư��W������e��,_qj��.�A�-٘��f����U.��@|�8q�<H�.��8+��\epŠ�J�<C!?YϾi哌��"k�fR��\rh{���VZi_��7)��.�@{�"!��Se�G��F ���9~�eMǤ�%Y5A����2�I�J��I��2�u�^����Ae�@"x���؁��i�{i�~��L<%��O��,.-�f��PyhP9�O�^�*��t���N5i+��T_�6��u����g4@8�_fg3��-���$(��������N�� j�"��$|��X�ɓF��C�)�A`�V�g���l�>ڃ[����v]~�6dc5@d4cQ��jE��|>m����B�h��f�Q�nV���?��j�/�]�9�j�y���"g+k��Zw���[ڠ���q�{��z%+�j����3�^;_�y�Whk�T�#X�&ȃ"��ne%� ��%<��/�`ely]iGy��*���é:�S��j�U<��� ��K��M`���x���x��������cd\G@�&��z#=�� � �_�o�x�P�Q�`��6�+3�|S�X4s���VNl���*�����⽶�����X	���.d����|��4�G`�� L3��[G�UҢ3?����q��v�f�+����?����a�NtDJ�a�S���j(�uP����0j8��q�����)��=ؔ�Ccd�Q�Qk1XgKS����v��=��0p1�Rv��������d@=��G�Fw%�Fz����Y.6�O~��R�a��A���G�
b�V�
l�t'.#��Ǳ.�6�+�W&�k�.q��^��=��0�D�S��Lfه��s��sћ�˖�X���w�82�N��!��}����Z�[�&gk�������v��nHD��fzC:�~?XK۫#`K��m�#d5�O(���˵��nu��}x�Պzd>���|�Cޣ��m>G�P��]�[MYI�h�,(���/��H_x`�z�-԰�m�� 9�*�%K����J����q5$��P*ߚ?yh�i���{ke5�B��Utu�=�7�v¥<"���0���,�wg��>�ǧ�np���<m�$���xX�q����T��Ⲯ�� ��Z�3٢$Qe婳���ܹ�[��N��Ib��Je�"t��ل��F��	ی���dAKc���C{*������Ѧ�z*prΫ_&�N{�=.bX{�~@��&��#�Ҝ�y���YtU~A��.���S���߂�b��l��b.��X'1)�b3������l�����o��e^� �̞Z�fAȸ�T"����)���G��s=m�Z��`WU|���T�V��s�����7��O�v��"�g%#{Y��?�mvPXʝ�I�_��u���D��A-�[ҹ�&�",�,�DV<[�O9��m�^�n�tKgR��(�Y�" o����W�C>�3\�{@�K�9���1�妏�a-�`�Y�m�V5Iț|;�r�3j	՞:��4��,��#&��Z���	��L�Y���ÚI��P(�}?K�QZYH��/�����-���\T`5�=�"�C�� ��!��3���������p;ݭ�-[,՞D�S�8,��>�ƃ07J��呉���TU�'�ƮU_~�i��X��S�d��\�z�6��,���9/%?؀TFdg��w��o�+��qTkY@i��#�����"q|E�gK���y�� ��fBx
��9��j�=�gZ��i�Z��◁[��U-i����L���%1�<��/w��L���)ĕ�M��B�,ё�V�_��]ͣ)B7ڮ}��{���2�����vb٩Hhޏ��/?9�[B����j8�:>{�m2�vB`��E~��wN�~�.xY�\��e��[4ؚw�b����s�J����;��##�Ag�j��]-�����m��fv��p��R!�Z�;݈扭~@�U��Z3J:��X
�V]`�~�<ty����ވR�.;�nY��sh�7���u���Ue�³ޙ�!��9`���	�oϨco�i�#�zE��ƏpI|�t�y0�T�Q0J,]����a��(F��J]�]v���z�a;;1;������ա�咖Պ���:�|F��5	����h..���E�(���4��3���4�� �Pd�|�U^|L=� ќ+������C�3��xW��;0R��ԓu��1jw~#9m�9쓄��.<�����w
s���ˮ��阀巟����I�p����>#��ʪǀA�B����9�[�=�������a���H6��Ϧʚ��({���;��7\d���5�_��d��/E�VV%u��2	��ue�XeN]�x2Q>��J�$��W���`��j��k���N�����b����B��NP�G��}���h�B0�4}�m����&�q7�$D���C,%m��ӻ=�'�`�,��Ch���+�M��M�bM�
t(%&�<\Mu�H��ڦ5�H8��z"y{�52�NV�C� ����iǢD|_�<�O&+����q��-S=��Ǭ�tV$c�+���<��7��E9 �:� >[k6Q*��i�@�P܂����,�u�{~<Z��J\Rd<�a�v���y�����։3�y��Evɵ$��������RНg��j2LV�vsP'�Z!1����cJ���2~2�����������d?Cmh�^.��e��lmE\-���O�Y�1a�*
	��R+��^����f�h��2�NU`c���{�QBL\�~�Ş����}٥����\��F*8���)<�6֢*�y=��vn�;�+U�R���:���_��\2�nv��
�oE�|����t�(F>� "����w�����xA7�Oa�>k��A�H�% frY�̱�0��l�.,������]���Q���8�bQe�Wpތ���50/y�?��a%�VQQ½,�F�;���}��W^4ș��u4�zl�a�ˡċ������ yl����i�Y�w(]�M{��l�sx�?��EN�-{7�gx����oOUY+���[�"w�T0ͬA�"(F�g�-�o�Ԃd����aEe/���Lxo�O�z{�s&B����^P[S�a=UY�b ����Zh��O-G��|�]�L��o�zŸ;����%1�E�k>T Ȕ�`ˋ�bD���o�P���k��,c����rb�j۝��݆".��!�kdS�&-�1s�cx�R�=��U���?������C���E(�2-nR-V#�<����XȑsXg�`�+xկ˃Wψ��}5��e)Y����'���"���#0����֠[^+9ffJI탦[M4�TL�ZT�Ӌ��{n	I�	�Ъ�����e��U���,T��9W����J��Z�7W�֙���Ŭ����Y@���XDm���^4l��]`�%�D�;
�&���/c_��8m6����NXV�� u�xQ|x��>P�BA�hqUq7v%<QFm�N~���[�u�HEˌ�"x .�]4��3M�$���\���g������~���8�����E�k��;[ʛQg���q�B����4�k�1F;HH�j����Q��`�S��"t�[�+��.Ѓ��>��
z���2P;P�9�fw8��U$!,�':�]�٨�!.{�g���(J���82�-���[e�G쀭��F(������d�8�N��F�E[섲p����J)���(�'U���m7��Pea�۩ͱ��n��@�c�k+�5s
�Q�%��G�Ё���tVV�]s�u��!��/bֵ���?�	/{��8��� _
�n�X`����ds��de�L|�B��8-�}ء;z�M{�S�I�\$�-F�N	ۉ��Ԫ�4�i3�=�뵧}�o���R�B6�$����U��y�"|�<q�n߰إ�[�ֹw�	����l�[���,l���� RqC�v8�l�ܳ_�X���Ҳ��^H`X�6S�o����?a�2��j��(1<��������ڮ��η�Q�����e��G�D�����j{ĳ���8e<�[h�MA'��݉� �{6�7k�BG�9Ջր��/�����'� ��U����X� o�N�*�:x��_[p�)��^��n�J�q��hy�<�,Ϗ������u�5�����%LV�].ǯ�(��/?��O�/����ڥ�]�|iQ��>�)��%g�!�^�6�D"��U�������Ћ����ߍ�@Ո�\����u�
�J��qnc,,@LY,�����X�Rw/��Fͪ�%>ƅ��hpoD�����Q������>��w����f��r{S-+ݒ#��M9�WiL�Wx�[YŠ�[RlY
{�~�0U��5�v�:����VgbLFS�ΡX������|N�8Ke��k�HM�'R�D�Ud`l��O���WP�MX��=����?+m�͢��]C�Lqg̭�Ȑ{� ͤ8v����}H����'B_<�mDW�+�	�v��c�u/-���J�4_��I?�U����
��0*.�ΨP��D�댵%h0aR�gn�^����{���Z[��00���f>��Q3W[��������@O��B�*YEZ�1�=^\:<��q�-��6�m��)����
�IKs7޴<K�:���hb�Ix� ���EKj�WȰ�I��P��7iDn�	?gf��9�g������ڰ]m7>!?,K�+n� k5�ڌ�ھ��kH&`��������x]�lƪ��^J�a� ��^��Jg$X���x�w��%4� nUX.�w�Sm{M"i�F
e��I���})��CuP@��4L���q��/QJW�i3}"\wY�������둕v/qA��~��%�c��D��e�~iؼt�"H!0</�%-� >�l�v��"�����p����gJ�3>�X����NKiRzkZB�V�|X�:(I0ȷ~���x�I0=�-4��9�O{ع�ֺ��À�����ԯ��Gt;R�.���͝��O~D4�.��ƈW+�"#�d[ݎ�XB𥫒��s�	��Ҍ�2cqv���1:�o��	�Oe���'���S������ޔ��}�kr���MYK�q��FNG���B�N�k�J$%�|�'��]��DxV0�wN�t�=�d���ߵA�P������y��ݛ2cXHU ��%}��q��`�Ǝ�4���&]a� Q�bW��V*j�s8c�gT�\h���%�b[�ŕ:	���E_�7O�0�){νLh�V�-�o�iO;[P��"X���+1�0���
+�s�w3�NCF|�b|�={�1��d��7�ЕbZ��PU����N���e%H?���\�M���J��R��?1���c��ڵn��T�M��A߹�{L�?���
\DMT�\�����w��25!"�6��/��GH��~;pl�
D���)Po(��CD�8?6����+{��i�ï�"�>,<��_��h9��>S��ø�gU>�:gB�$��0����0Ge�B�A���*��A�qH��o��m��鲘B�ZJ_[�o�V����3�����5�	[�}��ķ�U��hi�D=�8�	���yP�i�33sw�jB䭛��"�b.d�a�јa�?5+t���j_�_i�
H��ˏ����]qk�ʙd�%�q��y"�u`�Od�D_^�	[&>S~�,]����f�t�'�t�g�\���4���q&���伷+��o�FJ0��t�*�R
4���b�X^%�,oɖX����(L��*�h)W�������[퉞V�Vezoju�Rk�ʜf�qC�����B@���L�pE�%�*B��?B�6o�`���|����:����e"�/FN `��t@�c���Q��aJ�Z�ik�?�' i�0��=��(�ë&�l��&��"}��x���[¹	xص�v��Ƭ�qܺߢ޳�Β~�]�ီߖqcE���SP`jȻ}_�D��a.�	q����&'�/�}�:�7 _��|,ng+5���6	2e��e�L����ϕ���	��W�����T[���']ٻx4s�W���+3lp{�vS�&e�_3;6�Cf6%�t���Lw��5������¶��������v�n"�}G���E��AS٢�}����ߧ�4h�I]
Vxt��;,���Z8�R���O�\a�%�єŝeȠ~�0#��2�UxVa8XTNm��?Rd���&����b�_�-�Ը���S�ljT3�������meC0�$d6����\�Y�:��[G|I�o�I����H�C��ƾ��\j��Q�SƮ0��C���;��4v�l��{�4s�:$�V��㼃	��~:�#0Bg������v�R��l�q�8X7��?���:�"o�L��zh�Ë��*qE.�Eh�͔+��W8�Hz.��a5/�C�C�x��]kg.���¸ީ@��9���H�q5O���:�)q̏o����n�Ruu�M�։���|Ն�E<cݒ�J*����=p��qXՋ��h�� �Оb�E�m���2�1B�B� f�'�C�S(ZF�'Z*�w�$_��
��B��JQ�m��WҰ�ʡ�&Uې^񌪒�@�;�5��g�����$KM7J�n�÷��1]���42 u���i??�w�fsѥ��Q��Z�`|+��»��b@e�h�:���$!�m"+��5E���I�P�#j�7��4����E����A��P/,vt�#yg����'���/��8�NP�C���Wy	�G4���ߝ�V
�.,fPʇ����������z�f��G ����t�0`x���$����W���"-yg �2�|��s�O,EO8��$�O�a�������O�1��^�8�
%%)���Y_]��{P�\��>96m�$��J����-۫/���Mj^wO���}��O�J�ҡ�e蜁Xܙ�[_F�	)�0;�w��1B>��$e2�!8UȮLNb�+<�� �*EJ(�G��i�.b%�D���ɏ>:3���cOi�g;����Zv:���t�}P"Da���vV6�Y��"�r�=Z�$��� �7tx�hخ�>	�6)$]��ۍ�^	?��ώ��.�ž��[{ܦ������B�ĕD��h~ �a�޻��~dFm@l�hg��~&�T�����笪�3$xᏴ���V>��{�( $ܛ�غ+�����飦�i�U�Xv��'�yV�mK=�r�̿�bg�8@�r��NT{�s��(���2N4�ʙȹ0sq��2����'�_7�����]��9�Y��?��P�%T�U�Mk�	����@�m�Rd}&M
X����xT��SG�҂��e@���#a[Ms*$��#7��4�3�iI�בֿ���K`���_{)&�ח�QY"�ڧ�j2iQ����������6��|�/�$A6/}�}wE|�Ia��:|��6��gF��kY�1��يT٭�z`�'�vƩMa�y�c�+��c��Z5��HSI*�B�#������E~C~�D�'¹��վ%�
�r]0c���]N����I&��@#ٵ�5��p|����ϔ� �O��9�Բ[��m,t?����1����ɘ"���<�IYl�1�,$Jja���F�<�� �F�6�J�v��P�_X��c�ٷ��!��������oя�"��[�J-���&Bվ�F)ЧՀ�� VW�^>۽��Q/��6{��K �W�����o|�O�3ڌ	�Z��p8#����	�pS����r�Ǯ�����ꀸк��$(J��oy���р,�j#��uӰ8A�����*h}��O;�A���ƚ*�*�s��g��RS���Gk��;AS�=�o������d`��c�*��o�/=J�J��2����)c>��2�$�IO�X���m�4��"U�.ނ��ɔ=,j�)�aJ{b��"q�e\u?s,}��/�������h��jR�������1�6i8��ژ���O�A=i�E�Zr�γ;�T���jWwM%��Ϸ����>Ľ�8�P�	� h���z�V�����hSs>��d9m��F�f���� ěH�5�/͆1#�*��/�����i��X���k�m��[U�uG*���ZO) ����A��gB�Lp�C-���Aq�߇���YB�f���j(��'kM����v್������DqN�%M�0���o�0�u��2�����g���N)Z����G�3���U7�����S⑨BҨ����Hx�����~F��T;�|��D3����P��������AV���3F'g�o�8�G6z��n�%����6\�+WVb�XG��qxM�S�)�)jjMx�y����jƋ���l�F�
�����X"�ް��ؖ��]��4Q�����Jcva��G��`�j/��zC�{3��\��3��v��	���^�W?׸�c�A]C�c_���(���lXO���M%Y�cVr+7��Ƅ���m./N����b�5b�Hԇ�'�_$j��G���Զ�uR!Z�w�	���x�T�ل��a!6�-����P�,�6�y��D���_�΄x)A_��e,+�x�*;U��Oc�+�%F�F5��)���R#{Xl��|���9P_p�� R��<cC;E\�M��ǕB�p�Zc]�M�.v0D� ��gbi9� ���#��Xj<%�8���w���*F<[��I���=�y$x�4Rq��_BXg���9�N -4z�T}wMkau�e��l�}���sڀĪ��{^�I�u4#��҉o��~Olx�,�TOo��ŝ,�z"���%d���=Z��V��?����5��.nE���2�:(zO @7M���ޝ)�x���6~,`�F�9�i�|����KY�H0> !���0������[��� ��ݓ�w��A���``��B�T[Wm�I���H�H�~�a�!�AvЧ�QE"a��u�O1�d����c�Ԫ����T�>�flC�KV�����K�EPU��Q����)P�����֨`'+`V���A}MO��:8�@��@��O�yyp<���SK׳ I����:H����Y(�e�C��W�Ɣ1�FE�0;ya�d��U@ ]*����gɈC���$�=���Z����9��7p���R�Ĩ��6��ZFGf~x�F�$͒/ZW������2� )����P�Э�%��M,��f�b����FV����Q�+-8��
1� �qӂ����I	�>�S���P�9���(҂��!z3��ύ���q�|Ie :_�?�ۢ?�[YD��_��-҄�N�/�ݸ��n����AѴ񬀌��o�����(��1�a�o\=*k k�B�Wٔ����]( �63��i�_^y�Ě�u�(��x��˗��޲����3�k��[� h�I���4{�%O14R<��z �C�$D���N�XJ.䁙î8LS� |̟�y�R�/�P��`�*-:� ,��u:{�s��3���Y����*4?�׋
 ����BQ�bݼ��i�@�윫g��30U�`uL��z%_|O����&��ǅ�ۈ���rt�V|M�"Gx�ԝ���%��>K^\�!�������H��4����zx�,$4�x5�m�.��x��[)�(�H`i/�`SK1�ݟ�"O]�1B��p�����>'a���m�(�}ٔ@��$�w��
�:M�Ƌ-�#S�QG�vV�˿t�"m�_&����]�B�b�����Դ�Z}��w�ߓ��$�#ao�����օN{���ޠej�U�����!%اF�-:g�䅒���鏪c��6׫��<t�я����d��3���:mQa<��lW"x��fO�2�;ۃ�ڦ�G')0�kr�!��Y��<�J��1�u�-�S@�^v�91�"ٿ�T(Ji�1Fk���\7�pa\��IX�֦�Ỷ�.A���]�B�g�R��_�J�3�����&ӂ�r�}
��zJ��B/�gg����(�$%��j�V]��Û[*^?��M��²�:弛�o�D���Z�;���tM����e��	��p�mx:�9KADk^5�cu�+u���90C�Q��7��W&?��D�:��+��"��G�*�����B*j��0�����Xy�J�M�ާL<0�,~�$�lt�&�K�e�V�����|O�6�A
Qi���4�[(�nt��`�M��d�o��:���Vg7U���F8_�u�D[a��0G�0���oGr���~/*#���ؖX)��vGC�;D�uD�I�/f���*�9�:����#>��i;�1�%���3]��G���*b��FYB࿾=��)	�a�}06�<��a��#eX�*�����s5G�G �Ѓ�ǀ8^��Z����kz�r/ͣ�,���R�)n��,�c���D7��ɮk�2�h� w���=�u����M7E	�����9����5-�w�1S܂c�q�s�P�X>��֖�)��8`&p䫑J%���3T]��s���U!��u�:Ol�`0�Su'/�t.3ƻ^�Q�:�d+T�����S^��)��#v	��W�wl��ҫ�����MS���,Sn`�l��}�s^=M됈H�)�E�,�3�s.l����$�F6�z��A�^o�l�b��:�1-� �g>:���x�$�����eT3}�<�H����Sӣ103G��Qzx�M|�2l��v�0p����ߺ@�t>IZӫ"��C)k� �k���PBu��Z{@Eڲ{Et�O3��*�K���23�B�~M.�C)���W��SC'�('�yafm�7�%zj�!��u����$Q�Um-.$�M/�
8A3���a���a$�#ˊ�r/m���)?�pa��)���uJ�3l�(�f��q�gCdαѿ��=?]�$TL0�4< 8�:��T�b��3��p��d���0g�Ң�{4I��:X�n Y��F�ӵ���G7MVC��,���r�^D�K,��BH���O*�!@Eޯ�R08�#��a�gs��_���,�yRa��ޙ2*�7�S��?W�D�:����_��A��&P�yf�V��s�h���_��[|ǁQ��w��sB�ǉ�����{��ܳ(^S)���E����X�l	�����tF�֏�B��������A�����%��l1� u���oĐ1{ li�V[A�Փ�Z�{t��
��)2o�K�R�>+��N�\!�5�ߪ�}{1�(��8���^���6�Gޏm�n�����b"?�_�]�E�b�H�	� c|=�Чk��c�S%x%�
��+{���])y��-�)e�D�ZǍ��s�\��oG?�c�������	��ҬߜC�� p�8�W����� PBD@�p�*�������P���� g��Ni��E�y2��Rog���[��ܽ���<�H�Ү<�"��D�rD���'S��;:_�MA<t�q����\p}}��lM0� L�\Y'�bx��	����s�@V��<f�d�m�����wQ�g��z���;�j�EzI, ����W�j;A�Qt.h`E�俲�3MxC2��2� ��+Le"�0�-�ބ[B�|�����y�I�9���:�G/n�����cC����K	A�_ф���; y˜4�w>]6g�",��3��tG���j5�YB�kD��f�#�����禓�+���^�	j�A�g�v{t�;��(��Lwuw�s�3A�2zD)�o��]Q���(�/�Ci�I3;�U�/�[#��cͩ����	ǷFp��n�6H4Pi�t`��Mn�h8�^��P+�>;?�llpGov�)4wy���T�&[�c���)T�lL]��XC��Hi�_4�}g�I���n��7���ʼ X��4l���N��_������}��c�J\ʄ�t��F8!<�T�WV��lR#�}0�YͭшN�.T��4�:�xb�걿<�1ʔ�H�ϴ���!2�֏��,t��~�i!�ZG�)(��8�D�)�����+z��u��XVκ+���Hf��`�$C�ń#:�b��������b ��Nqm[o$tqr7��:l%R韥�n�c�x1H���e]��}�߅��quy�g�vv���G@��]����N0��]�r-��Nۤ.��Lol�4�	����m{K�Iq:�v�L����p���i�b��`�l�w�~r3��VRĨn�B?��ń���{[��
��D@�Do��&�a��0=��1Zβ�@��*�Ž�zs�Y�� �Q�}�B�6du���7冞T�_�ǃ��4J��D���{G��&��NvB�C太���THPih�M��+�ȵX�n��� �5\�n�	��M��a�i)0��Of���\���ui����at��f8p��2IP����C��C_�7EE�e~hG��	��G��2�a�S�e������T|�
E��w��L���2���ݺ�D	ך�?��`��� �}�8��ҀJ���i�.���(B�a9*�ÐX�5�W=5/,�19����n��R�Ln4x�^!4�.��f�眑��g��zT��lX��6J;�c���6��,��:�'`����+��J *��f�}9�B�(y3t�, �&^�B}�"7 =G���E�)&�p��o��8(�G�ʰ�Z�>.1bt0~s#}��(�{$��;� W=��4w�}��BF��ԅ�
sv:��,�`��̗չhw��t��l��0
�S����<��$�|Qh@����i��/4DH��ۀ����stX�5b��rT:B���oc��]�^��:��,�;����)j�K$��p���~�C��=c�3�~H��SB��*0��ϛ��OCɱ�A��o�^9��'�B�������E��j*Ivh���/��x���R���@���<�"�XQظ�;�^�bzI��m�0��9/��j���=��V:�����z�Q�U5�^-�p�a���ć��Nڬw����[�m ����|*,����!�� [������o�1�CA���b�/x��`z��0g���,3��Zj����p�+'
�{(,&\������	|ێ�0��}q)#�!�/�jl�t��yF�xk9��tP��Y�Y�Y��wG���#'��@���۔�c�0ɵ�MZx���
�2H�6�x��
���# k���A��|��!�ܹ�Y]���w�~�[�f7n X�Ȓl��ٷ�C��>���*h��\?�/ҕz�[��ld��S���+܀{|��=Z߲��������Ō�=X�>�߇�ʻo߶��JЪ����tݴ�fՈ-�aG��Э��i�[h���P�	m&|����ϥ�g��&���kn�uo�e����M/rRP�b(Y��&wmP"�jR��-Y�l"��Փ���e��ξC� ��\p3���V=Ő唠]�iP��?�)�����c�Xb�����~���*��֌n٫�:2F�ոl�<'Zzk&<[c�^'4c�����5W7^f8�g�"�McT2���K���?߅���s�Z��z'j���q��}��i<xw��y �t�zSZ��B@�~)�:jڇa��V��i�,�WD�ˈt ����e#�z���nei������E��\bN+��d!�R�\�T�j��'x��[)e�WZw� xɬ�O�M����u[���6h�Ӌ�߆���\��f<�Qԓ�Ԃ1�hI3���F_S��KU7�n{�Ş�zf�c,�}~:��Sf�oK��Qު�� ��k��Ƙ����-�)"񠮿����Wx$�r%�,��}���X�
U��w.��a�W����v��'q�ŉK���Qѽ�"9�c֣y㏤<ڦVFl����w�)��Y����i�5lq|j�Rp}���
T�B�+����J��Fr�6<�	,��Q���Gw#��,W��]������d��)�F���ޔ�k��bA�cw��-(����Kh�;ROW��+>K���J�+��<y�ñG
G���rW2�����b�֔R)�%�/��q��]]��G�'�p�7O��U��Փ~���bbEn�j5��-�N��Ь������0
N����Omo�-����ђ�I|TO��&Aj�:���
%szL��$������f��R��f��`��བྷ9���bE�x�s˓��Ė�H��7��>7�і�쓩ϸ��3��3.B�A|^E�
G��"Y�X�Uy^��� ���8�'[o�A�; TC�1��:�K6�\�	Ǽ����+�"�MļOѨN��@B�d����*�b ����O0�}?�
��(-l����As�	}�۱T��y�~��b��SQ2�+��߬��zZ<�6��ʃ]#e��}��.���_�+-1�s�q���_�Jd�̑�h���-/��zx��zP�G�� {Rz�sF@�l�F�}^�ȏ��m��UN&P1���3�t�E�Eï���x{/�T�h:�R�����#��څ��%��o�;��Q=NCo�<Z�N T�t �3������Bx2խ?�w(�@r54�������ǫ+ J�,�m��KC)�q�k�ؕ�(��ؒ_���(�~���x74�h}��TG�.�Y���و@������OjvtQ9�E��;�h.�ߧ>��IsZ ����^�Φ���b2X|DW�=L%�ΐ���c��J��Z�gׂ��;(#`����%�W��'+Zc��y|RB��� R�YT�?F�`#��
�0��\/2/c�X��I-�'��`L�r��S �'���p�$R��-E��,v��r��3u]V��c�I�	�<��DC�]��
b��j��(��:y�8|��dnKF�'�ߧ�6� OF(Z�7���f
��N���hl��tR�&x&��h��j���k#M��S݇
��'���q��oV�]�\��׻�)	��h�^X�[����� _ 
��-#��Mi���bURD2.m�Ù2'�$uV�8�N��";.䲈ji�eCO�7��s�(�K9���QWk��
MH6k�*��J��5����>�nQr��ߋ���a�V�έ���'��}�A�d� ��O%׿������|Z��)g����Ql��$�F끛�22�Ո�@)]��u���5�-S�e�x6s������7�x���z�B��y\e�TUv�R�gڑ�=^峪Q�N���p�#j��0�%^�N����R�˺z��WD���
��*�6Ie}�
���nC#3�]x��h�*����V3ϝ�J�<�dyI�U���_�P؏~����o�e���;ד��t?/�τʎ��c���t�r��V���Aө����r������.+�pqNb"����y4Հ&B>�%e��$�:rjf�����xt�)��1Y�9�0����\�$�4mhYY䛠��!p^�g�S;ф�]n��=�p24��EU��O+��%�?/&/�T�Pz*55��!cXm�I�(n4��:f:��I	z1$���c��� �$��ٿ�{�����fր���{K ���-���9A�-��zZ�=�6L{�����Y�(;c�nD�����Af��f�gҴ�Zk�W@e̯.��n��7u;�<��=�uG斥���؋:�A��;���s�l[.�*�_�Hj��W�Fr���u��%+dğ�?�x4�E��,E.�蔡?n�g;�.�Ob}�G�:����K]9^�n�l�**�����`��1o�N޻z�g�(���!�ܱ��
@�9��{م�C�����8�HlS��YV������ɄN��t�e�S�e�k�/�M#�o��x��1��V�O���� ���lT�3:x$�.�Û��=�$'_�8�
�U�����X��R��z�ީ��F�`´E�c��c���'� +���ޅ@��:�>-@PIɺqMS��C&�c�@�yP_�&DQ�/$���X���� �Qֻ��@u��|R���^$~��K.��Mќ��5�5���( s��wsq��ęYW�R9��OY_�aF	yY�&H�[�S=0
���l�HoM���߁����M`�3V��ib��S�B[B�yQ�[������ɧj	�mEz y���8Ka�`����к�ޡcmtd��I*]x��B�
�����!�6��G\A��D�(|����B���H`}��G��j�%�D]Ъ}��So;��!�%�E�q�/g�X�swb��P��[��L�wq�;�J�G�fL<J�#AB�ϰA�ޛ�_J�7k�({��!wyF���:w�u�[J��Ȕ���6�,���P�F��������"����&8)���	^��+�<9���k�.d��˓�@I���\FQ ؘuٚ�#������@|�� ���c>%A���Iq�Gt����fAV��u�tcC��>�^�$��Q��W��M���ekL]�7�j*t�N$�-��n[P���Nc����("���x $�Sm�L��7�iX	]:��k��[K�-��c(R�6�l�5�Ӱ�A���`V0<�R-�����[!���,X�����վ���[�O	J��I��EgyLđK��v�i���K������9�� yv��n@K
$6"[�p%J1��+D�C�K�x~+rm���?��q�%k�~�ߚ8�x��v*���$g�,����x�\قL�w6�K���l�M����ē���W��R��%7C��Ik=�~���8U� ˾s�{��dB-�B�%��ѽ�z��V��3�xB�*�i:�D\f,A3�Z�����ND=��J�.(Hi���:0���Z9~bÛ�"V���¿��SB7���=������Y��δ�j�2\��V��{����Ec�&�MD�a�~��(�J�43=z<,u1T�`���7��q�(���p�r��Ȏ��/��0`{S��	����ڼh_|���< V��W��wL���+Hq����
|������Z	ڂ^��n�ۥ�75h����Iy00
�`K�$�h��B�h�_��lu&��-v⸎ߪ����g�i���xp��-���43F����恷�2�R颓���:��A� � �S`��N(��(�G����ҢSt>k=�ۧc�$��>�]Ւ�#�����h��i�"A4�B�\"���G���M6�u���ŭ0��O&0�;"�=ֱ���&U5�ֳ&�����gd�K�ʨS��q�,'B��'� J�������b��l*K��+"JE2F�4� 17e#k�Xi%^u�E��#r	�'��R�/}Źq���7:)>�Xfj}�6`z�=,��{7:Os�k�|}8���5�P8��6��K��!��l��h�$A�.�7|����H���F��[?>)T@�7�ƚ2�ڒ���إ��8��:؀��r��*9IU+"A�y;0���ǘ-�}���3��>u�ҏɑKt�/N�>�>ڂ�C��2�a�C���
w�hZݎ�{cFLs�G����d5Ϗ)2��?^�!���P6]��7	�A`�E�,�`x��%sҗQ�w72�"��c�e�j���8H)���ߧ�c���/X��-�Җ�	���V�E,��Z�~�tWI/�*��q�#�z\�US�r,�,��>j1�0+���KQ=��웢�L�������)��*��j�X����'@T��=��HO�B8�K� � � ��]ͩ��F3��5����0��+D�Cky=�����ftg'�yl9�☨�@�����[��|C_�|r��..��ʡ�$�]�I���x����o�(�#���vq	AJ@^CXî��:OYL%�G��B��,T��K�K:o��D�%/��O��J�׶������c����ͺw
��"��,X��j��[��ī�$��fBɠ�y���:p?������oi+���+1�Gt������d>+�ȋ�N��c��;�N�O�l;��e@��|�5a
_��}��x�a��X��w�<�%�W��t�6��/o�ԭ7����H cN�_��u6a��:Y�e���W�q�*$O�Yb|ڒ~f�췶x����8B�$3��~�$'��}�U�:=7܎��6\��=�s��,��[�o��S�5sчDZ(�k�L����tH�?�3�&O Ń�R��7�y��յ�'�yySe�/�@X'��C�]���
kS�OG8����a���O��P:<�"����[��q�*
���g@��JN��������g`��d4h��'qX�?�ϟ	�����h-A��:�*��6�t�Ԃ��a��a�'�Q��ױ�*x��"�3���
��e�)AB���G&��pz��k�:��kVpȮm�?wj�|�V��Ú��28�m��f�PO��_�
j4�)���V>[$UKQ�Ʒ���a���� rΗ��.� [��
O6�L`�OKA���,_|���!P��rE��;�8(�� @,���*j��5��{�=s���A3r�܎�G�m1���ԇ�D�����_�^��R;�f6p����mb��!��	��+���v�Hw�QD��
��NQ`H��\�5�B{Ͼ�[���K����_m��@Ru����l�.�CM��j���%�Bv1]�=���f{q��l&�
_|�����}$>m&B�qFMO���s��<�.����(�'���2��ߦ�ӕ��	��w�s���oɜ� |9�<�rP$y�F�Ɏ�W��ل@�ʹ��(s��|�~�K��?�F�~�����I!n��J�@��F��x�������z
ƀ-d=ӽp�X,�F���d�{h���#�1g�Q���!�?�����W��	@�qќ
�#�{xW�i�军V��Je$��$-RjA�EY�N���2Ebot�����"��F��}7����lOf���4Y���?�]\�	֐����7��zc#������D\���ra*��L_�W7}F�7̏Ii�N����a{\���N&3�#�Jل]�G�����O�ɲb_�r�)7e-����*M'yV6К��J��w�_頡�Zۖ�A����`�59~v�L�;7�z�w�ץ�Bq�+�O����w�=�`.n�Q���^TP��;Rr���X3�ВT����/���?J�Eg�f���OE�d��Хv��R�צ4 >>/&�|�.qn�;������f��zM��f�aM_��V�Un�C�p;��Y�́�y$r�*3��-_�#]F��w*DEI��Q϶+��?/6X��6摜^zQ�%.@.��~S�=�)�ŭY�++��b�ˎ`�o���E7���?�2+��2,N�FK�,�XۙS�@7H�+&	�.�+��{�����s�q�mφS�\^���LI�h:�����~Q7�����V$:�J[�<�<��M�X�dD���gl���:`Y��\��h��g�N���Gz���:�ʬ���%���
x@o�_�a�zy-�� E[�7�
�N�tt0�)W��fm1���=d"��g�PU������w/��(�I��H$��[�i� 5���E`���%/h���@���p�Eg���4�~3f���}$����7����D���r�b�1���a���\���~�M)�8�� ��5���,$��#R	2]�-3���#�xo�)��ꤚ#�����;��E��NY~᳙�^if�6�L��J�~�D=�%r�H���8�+m�Q*s��u�Md ?�ݫ$�@R&��	8�&�-E��9���i�c�tɅG�����$�*��D��e�����@��Q�H����܁a؂�w [�f�o�Beu�d� -�z�|4�}r�H�9�U�=�V5gu�p�@?��n6 ���y恍`�͖�)ہ���	�dLe���%���f႟ߚ�*�]y?&�o�6	��>1�g��'�cz�%��&�����0,�����,�S��0�s�ol�J��ţ���K�v��d۽\;PXp�i���$T�.Ie+ZΗv8�K��t'�U�И�����a���X��Z4ϟ	#�8���(C�>�s��uF��R1��xnv&P� �A:)��^��hf��[����+2�����'����L�![o2��sH HEi���r<p$�z/m�y���"���~C=�3�[@M����8�X-�Pa=:��Ӽ�}����O9�
¨�h���~0G�3Xfq{}5�{q��\ƺ;��RaSH��9���-�Z�!��'��7�ݚ�_69?&�B!�KDe�j����`��`b���k�뮢6�� t�f�jѱٟ��i5��Z��w�>b��y��GWfCY���\b��x�p��C�&�M %qT^6�t�������2�S�=A�*m]�a'*��K�*�c�ץ�YsE�n�⡌7$D������刭qj!?��N�c6>����Q��_�����*�a|;sr�b���CAw��!�t������5t�.ŷF�-��s��x1����b��<JR��J�����)����s 9�.��۫�\{x�4� :���Ɓe���:'Qe�ص1)����/j\L^֪P����̀`�, sl�np�M�g�D�7��g�mr&��夝��!�jRF�$�ҟelZR+�x�>���"���i�^���|Aw��R�/_K�Hঙ�^W����^|��]�U�U�p������h��K`�V�x_4,����).��Nf�b}���>�P[C�в�]�����M�r�c:�䂈��0!;.X��(w�����LE����Fƿ޲�apP'j.�r��cR�l��8�@-�~�z���nAg�(Ġ;��Ggmƙů��x�$-3f����|��c�I���k���]���ʪƠ���;pRT��7��$�n��R��g�#�mO��"EI��{U�::VD	�r/������1^����C�BeP�qG�ZV{
��{$���Z�$J��*_���������SI�z�?���r���L�iS=@�U�}�ф�<V4�R�\�L�g�����4VJ��"�����_\)9�72̰��rt�� zK?wlVO���غ�M#��>��8���}��l���T[6��"\�/?f��ю�/ܡ�~���}��Λq��҅4�]7ޏ���[
��������8*���g2��szN��-9�)L���lӐ�]�� ��:$~�;kk"p�`�TD9�7Ύ�I�8��Jy�d���3���Xn�N�����
T����Ӄ[�5B��qe�bpnJ8����M�,b��3h�{2ֆ�"�u�^��B�c'��,K5�Ϋ�*�3�x����	�nG�aG!�D_(�a�� 0zx������klrZZ�WT.^D(�,bk[������"��f�w
��9Sl
˞~��c�%W�v�Y�ޓ.P%����� FF��B{��4w��S�^�H������8/��2�ѳ.�<t ����[h�q��U��&�I�C�o��ou͇�`�=r�Ò�Lď�u��B��V�ƨD*u���H�A�Z ���O_K�jg���J+����D0�hy��<�wH��/�aM��tGP6�$zlq�ŷ�A���G�v@G1g~A�������M�=Ol0l!7 ��^��댜��'��J���ӱ��0C�PM�|���I-W&\9s��˺��s���,�K����L�hmg�݁��K)�� ��v��
%u�jB�6�,�־��m���H��.��;̨��`�*N&�];�h�_s�(S�)��������!�E������<��N ���(��gt�?^�3�����Y~�)ϡ��ٕ	��o5[������GG�Ե]EF���㖣y�4�$ZK����f��6����H��D`ɿ/�a`��sI���Ї���kժ���[�y�'�&���;��q#
�J��pn�9ji���\sS���G��[?��+@���!����]ѝKú�	G�QV�-��]����ˠ�pz��;0����di���X�G��"�1�rs�_)����gɚ�PR�o��)`�j�7�/N��! ����3V����$�A���aޯ�ѯW�Z�l�5d����h �,1�u�^��ߐVM.����"eLQ@���-����*�=o��_/6!���Q����M�7X���C�P
�2��^H[$^���x*p&;G������?F<�>���X�=�}�I��Ʀ\A�������	\��k�$�| ǜ�Ы�}���:�]눅����M�*�$!+]�E�8L�3�"5�VI)ԗ	�V�c� ĖX
���Ss\ܤ�Qݫ1M<�����21
*f ��/=��ݝ��6���^��
���F��a��n�&w�?����>)�0H�ɍ"�G��#t�&
�M�?�e?��n��6����68����M�f`�B�/^=R5���0��3N=F��T�mK��{>`!��&�[�2����n��߫��$�d�(����6 ;n1c��چb���R�?(�6Bȏ��̫�J?�v��`�G{�CE��ź���X����l�?�D�@�@;�ra� �6uz�0�!����I�+���6-H�1-[�4�OP�f����(i��T]"��v��,�O����U� *����:�Ƃ�1�=f�%������љ~�
w��,61cb��(��]���.�~�M@����*�i.I���,�H�!��q��c�݉Ɖ���{�"�������7+*�L�?����W��;�؀ɳ6��5��@[�Gu��ƛY�D�L�}� z�M���Ƀ�����p?����@��F�!����ym��hc�b(9!��嵱PR� �1wE��+�ɀ����r�.��A�t�-��%R!0).�I���^��a������C�*�
�8u��Ǜ<��U�����̷8��ÃZ�A�"��ط����fJ
��a5��zk)8�<�ΘB��g� ��(<���'�w�L���M���zx�B���OV�{'�e��=��c�μ�݁��ȁ�o�B�Lî�ѵ�݉�ěʺ
q��jTl��La��v����S�ۣJ�?��-9�A�zX����|,u:vU�O~Q�F��B���D�Wn0��w��T��ē�H�j̏��v�S׳"�H`�k��#��~v�np�(�"��'�B=�����qW/����}�X}�Z����t{��8���}���r���2�,�%�Z�Qh-�S��k�  ���,Ԝo�]�;R�
�7k�LK3��޾�1��d�ډ̒�"u����*F,^g��%�� %�.n����E8�������Ճ�+�x|��U��ۤR�G�]�u��E�
7��w}���yU@/&��m�}�!I�'���{wx�?���;2����lH��њU[~\�ԫ���Lo�>�@����@���\�S�������V�Ҩ���i�Ǻ�#���'1oC�Иa�٦�?؟���0��)�?c|�������Y��c�"\��^��"�r�p���3Xo�0�s�����,�	�x�/��O��[=dm4�]����V�mŐrx�3@p�M$�ȝ6�o��a�ܒ�*�����՗ī�^H/���,!�I
^�gWQa��M��6��~�7ނtw�Z�X<I0�U6�!7���4 fE~�R1�UU�
��C���V���Q���xPX�/q�
y#�����J?)���(�s;�\ݣ�t�9���c¶��<��d�k"�?��ٙ�R�U�<�(����	?��u��hĩ��<>e�1#���9ګ��5��^d't
�N�����=�5�U�!�?e�8���g�E�->�[�@F�'�`ό��t)�cy� ��jz�[�P��F�Xl��VߌAL��j�ĽTY[��x��]`���KZ�α��9���d1��l�����e��{[x�[�,�Ke�lT5�#���B�2�ќq뱈�j�bO�H�7���a���\4�H���H�kK��yPE!�H'�\^;ITH( B_[�m]���~���N�%�=�]�A��i��z����*:z��=���Yz*����J���-�ˠ�G%�8A��Kw�s6�WR�h��S�g]��#���O�/� �ɷA3�uub�iyg��Wu��cZ��G�B/����,<3���@�;�P���Kq�2ۍoȟ�}l2ر3i�.�(��Q��2���s]�1��8[C^�zז-3IJ� ]x��b�z��2�'	��(�S�e+�F���S�����`-�,��2���n�9o�����|����$%��W~����%�O"�>���W85��s4���)'���f�����P�L���	�-���iJiM����X/�p��#;�҄��u��O�<z"R�c
O�������+��J���YZ�4��VMvq������6إ.J]6��N��oi����2�u���5�1$�A�,O�,9~�J��/��$ީ�C*q�0N2+��ؚ�EM<�Ee��F@,�$�6�Μ!Ó�#�fX��c�Gfv��6,S�`��m$���v-e":�,L��es^�ZNɪ@�&{�\����΃h��q#����L�j�ݴK)k�͘8ֲ�r�?/^��{'��Ś��4r�"֝� �ǐÛ%�LX|��w��D�[֤1X�T�s)j�*�hy�!��C��UDQG�"�hB4�c��VƧ����$��F��^j���O�W��"oH�qZ�e�����Ʌ���~��+�ut�/9��s�����T�ܢ��W;��o����M%1^>3�(q�r#"t�Ck�o�����g�%�V���n����0[�n�&�4p��c��{���\�Z3�!�����|���P-���mkl%W�I��mȯ�m�z��nMx6Zn�s�
xh�"[VE�d0Tф�1��m��AuJ�a	���|�C6��)�C��[C���\7*��`y`cj�Q7j�F�ɋ�t���4]s_Y�Z��,\��g�(<�G�d��d��s�5N3��<��mӄ&�����:���������e;���Ep߉a�T;z4��sݕ�V�W�.�x�/o\���\$���lM�ç���0��#���>Z�q�D��ݝ�Ma-&��f�exs8�s�u�O�[���2���?KǴ*��7����2���)�8^24"��ܳ5U�x�'��ܡ�l��%SF����M��%�u��\�Tj�&�<d�=,��^�g���a�w���;)�8:uh�ă_~�E|��{3_o0k���p+��#=)�S/q�{�k����-�m�(q9���K�-��G�i$��B�����me�Jj�R6��x�:/>�`K�Ly�;�i�}<C���O���J�Hv������/ϥ���\$Iȧ��]�'QE�I��x�*���:X��[c��<����o�m6�޺�s*`6��X��Oñ��D�"�D�"j������]%\0�*(e�:�|Y3˯DY��있��5Y�z��O .�8��D�fz���:��aM��%U2�B�k��!�w��׷�<��S�����"���J�ue�W��v�����~�"D��F��K�	bU[T˲	M�� �(P�޷��B����Hz�)�:7B9;�J*����]�Yp�6,�)���1ȷ�+0�E���ShL��f�g���8���8sf5�LI�n���N��}b���?ř|*n��j-7��|�쭴!�e�鼵P(��Z��b�`i��Ϸ�+���C�L3s��i%��'l4wKkൈMiW"�ն��nХ���hF�]�����05�!c��3�g���Xe���mt!�Ȅ�^_x�e �)����I8y*�t#��ɤ;���\L�"�i.���d�j.Y�^7k��������Q��?EӾ��=�r��]��Y�a�]ۓy��@9����j�25���K붆�x�@Bq�q�o�7Kjo���%���r�;!C�0�*ܚf4�aq�}� �nLSt���t*y��.4煯8<7��JVVf��g6Eo��� w�[=��C���� _��s�6!���R�� ]�Ҩ��{��6�S����F��(�,�ob~��مDd�I��*ty�i�ɺQAU.X��s\2E��B�뷍�61\���+_3�U�b�ᦥ~O7o�.Y�ַ=�c7��HKX����#w��+	�t��_"3�a���E�%u��uO_t�`�dhp�}�5�A�?f�N<鷕Tl�����נ��S����!�c'1"��P�����Eїy'/n��L��X67�z?	���ڊ�@*%�~�o�
sI����X! �B�,�&���o�olŲ9R����ʞ%�R��KPZ�:��0���_Ї�D��3V������5��ݸe9Q_�����[` �Wb@�V�̞�����[ZJY��Ha��Q͡I�3h�B���.��	��%�����j�%7���֤d�r�[�����ą�* &$��">���x�������ҹ	�,�-ͥQ� ���!�N�G���-�9���B���Y��`�+B��#2Qz�e�L���t͛?3�8E��Z���3�?�g`��� ="@��a����O��J���BW��Bʺ�>3s�9U������@�z��"���r|���&���8~ߘ��S��V0���H�	5LQd����'��7jpEf��9��X�NwX�uhm=*���S�{q|�4��	������0^1��O��b���Y��j1J�o�5�P.��h10���:tc�w�2!|No;lc�:9]�{o�5���
�O7F��5Ʈ���,ȳA�2�!�~���Y��	�H.k�&��9^7է�Y�'w	����ݸ�_K�e�x���6�6�&[��F|I�c�az�ē������3.�1(�1��;�RNxG��8,.�Ց>2�����v���2���{`��Z+y��ν�=�\$֚�%"I:�P!�
e�Qa J�I�ͬo�P��:��$��:P�>��+W������:}d2-�K���"9��Ģ�b��#��A�P�W?-͊�Z��$%HL��.�xt�d������.�ܨߔ���ê�M�k^#NEz$m�+�d4���o�����[T���3���s�����A1��{x�}�S�`��)��ɥ*'��p��j��N�M�ah�K���P�ݚ}ˍ	\�-�Jj�@���y�ם}v"���k���\�&��d8O�Ùx'��}���a͓d-l���/� � �x*�"�P��bۍ��68ҩ�)��`?$��r��7#Hw�B�;+�R�f���f:��r��:lB�hh�S�tΑ��_��Rbw�`0��ے$�ع�D�*v�q�A{��"~������HIl��
!y_[ö6��#C�{tW����Z�Dʀx�9;n��L+�)���+c�
��']Qz�±�UK!�f�A���o��Î�I2J9�hd�3Zl˸�s<:Y�?�F��0!��ޖ�S��$�qx�@��\�<R�̟Ґ� ���C,t��v]��W��(�>�!V��;��;H9���v�AT�����ޙ/	���#�1�k����@�`5���k�?Df�V�=&4�JS�̧\z��L�/�X���s�;�d����4d��l-�
/��ا�K�,Pl�s��}'y^�zrS�ğT8��[�܈�ʈ��li��B�1!T�=#9��QN�0���\�jojr�	�#ᦺ�B¾��Ip���T�~�]��䮺���{���myd}�3��l�h�=U���4�j��8��a%�EI�
��r�2���!�E?tM&�����&k���L�QS�;2������~�Hm�.Fg�Έ�yّd=&p#� �m�`���ǭ)�|kCw�0m���΍E~��g#�O=���s5�uM(�K�vѱ&���AVg�O#��u;Ӡݪ�P�`��ER��S�b����`wJ_t9���X�I��ı����膓P�%c��0(	�̹� a&��4��Ăl�:���t>C7y$ߥd��P<����?�3PEJc���#��F�N���~՘�!�ԝ�9�픂������p���(�k���Y�V��@�̴��ap�3��5�|�t�b�C�qzг�j�t�,ڿ��N*��kh���m������u�=���r��� �;3���g��ׅ��4D,l�;� +��
�4��O.S��)��� �Q�#�d�VJ~џ�PfΊ` [�$1W�rm@�oT��$�?��c�Ϣ��������	*�I; XOF	M�����e�>#���&��_�:�t�����hj��݁��`�ӝ-x3����Y]|Ln�z{pr��(a�u�e,L�S�d�ޢ���o��]K��[vʉ��5A����g��vI���ㆶ�2��s�3D�)�Պ������'���a�{�
�����'�����R�Iz���	��Lv�+K��_!��T�Ö��������x��?H��cTB*v ��A.�<H!����I��%�6��@zB�I���Q�i�sc�h
T�a�T�uqYWp��RF�ļ�L`"��D�
%K^��|t����Xp�J�Uz���B6Je�_���E����Z��_1�)A>�߻�T�T2�Ѽ`d4�'�X4�s�ϰ������W�7�jjgʻJ�L��H�$Gl�k�X�rU����1j��gO� I���7&�A���}�	�����	��Ph����l�-�4P9�G��'0�z�	�ӂ��]�՜m�iݎ��o�^]mz��=O��|}��	Ɓb!�¤>�������tlIp���!�}d�d�?X�3�
�����z���k-Y���$o��'��-.�}��`n��  O����A-w*�g�gcwO�{��OӋE�_=�ǯ0@�v z�N���-��8N�nm$,[T�N��4�}����c_��� ��78v�{	��꡶�AmQ�N��toT�@��ٚ�ň� ��6͚&�a{�.�Z�C�.������*U'�2w���e����y{�ŝ�5/:����R�լK�?��+N�%5$m��+R��
����&6�Sd��8e|���-Կj�y�T$
y���ܬ��y�Xx�c-�d@��}��S먈�6��'Ǉ�`O��k��5nP�7�\�\�|�0XF%�/��z�F��2�6s������I�%��L`��7�>j���tG��3|�;v����%xVj��_l���yZ��`Y�4�Wy�@�G��#ޟ���k�W�*�4C�^0)���Wo�"\EH���`���WƏ;��C� �D�0��&��]>$׏^��g�A�%,��@#=����������{��T,�*8CUR�jQ�n�Y�%����_ź��iq�'������y�^�E�sQB���pU�Q%��[N�P�t�)*��J�އ�b��sj�{]8%�|�H�&�!p�������\��,X��y�)����S�P{��HF��M;����w�3�o�}HF\s��_���m��/&ې	`;ϣ1�VG�����a�搘�G�ST����2`=�1a"�yWg���4�3��:>U!C7���g����{�Ёh���������$?�= ~	V{_����Kml�zW+�8�X�0&��Ǹ�[��A� ?�1�6�z������1(��F5���.N�J�C��8E��te�2
h���a+n�Y`��o��|Q��>���`�]�$H��Hj�M��ĎǿW)�r��;z�#-\�e��$G�~�Z07 &�⭦j�O����$�)���ŕp�~ش�*�:E�~�_�y�H�>����l\8�z���=��K�wġ�B����0��yǖی2K�<5C��Ƙ��&"��{}w�*w�j]����B6IS�p
r��C���,�S�ViHf�Za���Z8�]���{X	&���YK4�4����{l��?�T��h�W�H���'4BO��k��Ɲ	�qV�ѝh%T�Su\m?��W�jW�n��q%n�H6�G|EY��������� ����s$e���J	��o_7�d�ex01�6��V]vk�[Ip��ƣO;F�J]mۍ5�>f(��吏�mf%G�Ӎ̃�S���_��vE��11�)������N��x�N%�o����6�� en+�v/j�:����s�4�S������ц�/q�b��q��W�\T�p4�ů��4�n���?��K����)����(���I�<�Uy�?,�-Ï�<�ۂӰ-���?U�h��lj�a���U�2��P;�-��58k�c�m(��ڏٹgzo�9.UPox��n�MRe�|�wSYG�!�Ɛs�0Y)x���j�a�v�r�F�HM��,�~"�STV�w��pf�dⷼ���i`V֞PǞ}U�`Cծ��)ɦ��ǗK�͹fV��Ք	*9�@�h�}o���k켕"vP�sm�f1"չ�0�ġi��'��k_��]tI�=�:�3E�I���,,� 7����p(3k����}mlB�:�QİcJm��9ַ�6u���Ƭz��+��f�$���6߹�U�����9k���h4� �ζº
>���+��;(c~	'y��|a��ٻ � .*�+�����mO ;�22h'b՗RCn����w�s�I��(��B�x9g٪���-#LKIzG*,������i��d�IA$9�HX��k��Eúɒ�cy�^����6Y��q�솪8�e�_���v��0 Q�	�^xߐ�Q�z�,�K�Tln�aԝ�W���d���R̚�����(�#>GA��K1�O�̳<רmQZ�'�bXJx��g&�Ŀs
�C-|ھ�6A�f���\�&_�kwm7�9^ȋ��70Ml��8�2$Lk�)��*{)oh��	W<��"�Z�������1�4j�RIJ�(����N*0a�S�UK5��3�jT ~(!����07b�S���xN�ut��RPc��z"�8�i���_�V��dUm�Q��
�{�T���/��Th/�L��S��b��$A�4�Ʉ����m��U�%���kT�zo�`o�WN�]��D���8�d0	��x�>��������>��6�r�")�?�5��~yX�r� �X	��S��zo4����4����Ia"�y��¬>Р0�w�T?��e%(���}����I��V޾(vC=�&?(\{�k��T�_0"�c�%�O�k�M�f �
Ia�5�M»(�.�+#t��nZ�g���L~l��	��t	�S�b�r�*~���S��wt�O�ͳ�g�`�yAv���Q�c$���4y��|S�)����LɺY��J܅�FU�N"��]��¥�R�[�hî>����a�	��z�{f�pj[3����+�2�.�N-�v� ��X�����R�Y�?.�+��i�i�p�	�y��oK`΋��\���+�TD���#5Ҕ��w3[J;2:x����	���Ci������w��Ȕܡq	�&3Mam��bg��	n�*��Chǹb�>=����ƧW�����:�)�S1�>iK���j����E�Ln��aZ>㣚�j�$��y�!�+�ܯX.�s_aSw��I ID%	C-2��;�^cyi�
�>I�⏟����u"&8�$��z��&ť�}(��2i�� ��'�R�wr=����IxꏁF��1p�N�o(��5 �5�&_��A�}
`C��"��E�_o�A�'��#��|�]�ӵ��2����ў��^2ϐ��ꬥ��G֯A�Y���+���6F�b�-[!�"����3��=j�y�"Q�3o&�Yxo� ����.E9S��h[{�3ͷ#�L��&|D�Aeٞ\���w�k�9�m3�;��Y��~���ET$Ю��X���B����k��K�+������Q W_�2k�~�և	8⏖w��s S����������N*�����f|/��iln�{k]�;��7!�I���5T�Uq�c
0�	�D-��/BO4*{�#B��D}Aցn�L�+�'߀=2$��煫��i��v��z7Vi&=.O ���>g<�� Ŗ1f0W�����g�>x���h(���L�W˙^v�s}r~�i��31=��˯�-�i&|���U6�0P�mt�(oe{�{�q	�d ¸�kb���9k�F����SX�kƷ�Eؿr�>�P$����'���~G��L�۩�+?Σ��҄d�Wz�����Jظ�	���Ĵ�-�c� ,B۶�4�8�*� � K(�3���۠���a
�������84�Z14S���8�j�_�=;��f��$]�� ��%�EM��w�l=�5��}�<"�
X���R�|l�zn���EqĀ�è"�I�f�,O��{�&grO�v���U�� �ie�j�-��(L뼘"SKi�8���֛���c0�t59�x�$��P�
6O��ԕ1Rb��6@���@�c�ez~f��3�e��@���3V~lizd���J��V@���yn�h^��W���U�Oq5[�D[{�KYtL���{i�&I���>b�$�F�B}]�;?�E�&@AI�h^�G��%������F�3��_dE[��v���$�h�a#�
�]#�G�⋐UJ���g�>(�G���Q��`�p��!O_Χ����}���؟��d� ��TC'��O�b�r[���/K�$��Z=+ϳ����~��R�8�P<5�Z���B�M@}��9Ǡ��a_A�Ɠ��L�9*�Y-L�[A���8���2I����|,c�����7��_�nz`��,͋{�K�F� 8��YS��\��2�=�D�!�������q�I�o�����%��kz��v,A3"��/�^4h�4:������tw��m@i��$���zE2���>�DV��a��x� g�MK���1���|4)80r�� 3�h��MPR*����\����kğ�m~��g-���:ė�����j�R;�t<�$ٱ8��Y��y�K��ш'��&
C�������>F�x�k
`Ĳ���o�����k�~K585���+Rp�\?)j�b��P<z|]���^�RD��Y�z��X�oiyK���R�"{�Qnjj����!�T�#;���wd|��v) |����/o����G�.��0�qfS&���ܤ�̍+1��ȺZ^��x��ޒZ�
�(ѝ�D�e��f�_Fb���k�`������V]?P�C�q^�i���gG��M�&铷LM;���DrIL�.����e�݁�)���Q�\v�bհw�G��d�XN$gf9��`��`�1��zu��r>������9��L����{�>i����#hn�-�![K�^	��{E+N�7D�I��{K�`��@��4B�<�E�N�sf��1�+���H3��ES�a].OY#��|{���AUv�r�xߏ�rӏ��
vS�ߗ�q��n:1Z�[=�)U�-Q�D]���ޗ����>�l�d86�%���-S�{W�n&���eBB��@N����؜�M�	+��#�/�oٍ�V�1Ձ8��7F�x� [EWŔj�ݚF��;�;�U�y�I���?szخoN⭗Ƞ~�[�_�e��ĻR+B�o|��{��M�������w��69i�`������"���J�WfE�`�¼6�ϙ|�s�!{��		D���a�t�HN���3�
����v8����j�8�3n�a&�\b�t��l��>��7e���(��WW6ޣRYV~�5�&�V�s~ೝS{3&Uǹ�}�AF(^�=�&����s>[�j��'6C�I��4���o�e�=���^t�|�k���`̊g\%�U|e��P�c]67�^��6�cǼ�t+B�W����/s���p��<�E��K�Cǩ�*��g�#�~�P3u@q~����ߚLe�F��-Sߝ��0�_#����Bz5BQ=�R� �l���!Ygq�n�7���	�H?xL,����� c��=�Zc��(���F7Idq1ڸ�&[z^=��I%t�oxp�2Ex����3��e� �c�$7�i��8��#��J�������e%�OPב��<��A�����7i�[U�~+����L� Y J>~�$Y�G�]�_;��>��LR)��0!���W@ߑ���w�m��˗����U��f�]ڌ���pbΚ�����0���.��B���j�꛲�r��D[g�K]e�W.�jn���񧚊����_[����o�t�&�.�Ƕׇ8:��A>)����c��&������e\~���� ���N�N�d�w��%	���jc�G�!�tt����R�&�b�ƾn��L�b�}��E�͕K{��URP���oig��N�z�d�D4��m.n��]�+�B��J	(�)8�Q!�k伍�]˓�>���h�t
2w��Q�e��d�?p�jt�p�ҿ8�)���n�`��6���>�Mkx���H��ޠ�?5����,Jgn�Z� ��|&�Q�ʀ蘘sUƳz���^�hҀG� �-P�C�3�����V����"!%}���
� ��D9�*+F����>�}p����[Y��M��UL�հ<U9;�L��]�Cyp�����/!����Y�<-�u	�d5D�'A8װh9�^��_\�wأ���i�����飑��qK�*��4�AO���3�_c�>�C7��t;j�o��c`s�JT��J�^�odt�eQ>�ܨ2B��$�> 4�^x�YD�2��$�$�m�	��MW����_�9�uln�o����k�_�0��:�;�B�P��1�a��� 9�'��37n@��)�	)�cIو�������F�)c`�2��dQם��N��	Gl�g���c�?X��4�O_�ѽFzR��4��вj��x��yP�O���K��/ag�6�_�:�P�˷�$�MJ£BL�ځ߫���_��A(����U�q���sj�����5���J���~r��V�Q�YfNy�r*��ө�̺kH�R~��+_ߎ7���,�������/V����E��Ҥ~��Cx�ыTm�eWoBږs�M@>S�j_o�8��`;�}h.�ɶv��4Ic�x�[��71�C���U�S�K�%���Rkx��ދ?,v<���O�t��Z�<��	B�#�p*`���XR%}���'و�L�r�P�S d�Bz��/GS6��R&-�}@-�܍�/9/�v�Z�S�g\�����D���A�6 ��LGcR2n�AtF6"����$�x;G�,�oe؃�n�pck K����7-Jzz�C��4��f�o�<��W�B�>�]�����J�A�\.�b�U����ky0W����k{�#��\T3Q��t���%��kH�ۦ[�
�W�Z!�Ύ��g#���]L^�"�#d��%c'ę́,{�3���/9ZV<��#|s�pL���m�OCE��*�6������CGT�p�~&�^zvk��+���V�8�=��s��V儆q��$ɨ�ڡ��̦a � 8�AA6���CY���,�l���zG2�)��ek~j$U���>+�X�MJm��j6��x��@�C�!������(��ٻ��e���e�,H����H~�ȶ]4ug�������.�P�^`�%�'������S�8��� ũM��-��E(eMY��pݜ����=�jI_R��y�)c�����ēv���f���d�L��g(b����@��R�j���ke��Ĵc]�������ғ��h>�4�%M^L�94�X���g�B��{��}������_�}�&y�e_]v���F`��$�.��1˾fo��?Tp�yڧ��NM��c
�kH��aM,�aE�R�C����0.�gp�dR$U(ͪ[�\o�:��cwe=����<����x���� �?u񬏍��
�p�G�~�u�?u/\w'n�W���Dd�(�
0M��i1�(�A�[�]��W؀�o��:D|��5����P�Gl���d:,e8�n;�{y���uo|��H���D9B�v~���N/��^��x��[b�r7Q|c���/Q{���W��F@��"����{8]���zKW��zA�y߷�c�N-�e=�&�cy �-�w{�?����> �|��I������j~@�0��ۄ���:����Z�����JK��Qpi��c��0/ ё"�������F��6��A�|[����Sry@N���~6x��@G���H}Se�R�����31 /1N�9�@�t�T�:$�3~����!���W*O�B��"v??0{y���(�Ӯ�O�-?��pj]>����A�v������%�DT���d����r�a"��p��J�Q��z�x�Ku�TR�6���O.���	ԧ�>\|KM>	��'��~u�Fż �@.��Ǵ��R�t@�=/��|�М�\iŰڒ����E��H��:�d�[⦯Z��,g��@ya������T2Jf7��.�~�9ô�FIbi��z�v��-ش���K��5@+D����� p&��	����5'hWo�&�������ʒ9�,�)�(��� 9i�v�<��o�u�U4 ���$߻�E	��>P�X��l�;��]a�>,�F 	�ć��(I��"�=�|�U~y����s�WM��9�݂`��)�5��]�Q9�Wk�)$�%j"��ƕ��F�pMɶA �bäL �b���gݭE`�^�,{t��M��9}�S�qK�������(�K���c\�Ĳ�1�ٳU�^�;w�c�Oa�,d�8�ϤGp;(��ܪm�0)���=מndy�k��^������[���-P[�n�a��V.�j�"�
x�vtS;[dʧ��_�Xs��ѐ�����OMc�JK�j�bҨP��T���ѓ{���Q��u�ȃ�J����s`��*!C�B%=m�&����� ���ZO����?+��D��/ȵ8H�v��N�K��_w+��;�t��=��.��3,�r�������'a^���������y���~����?��I�068V�a)������Njݻ��Xh�?y��	Z:hb�M��:Pf�&f�����u#�̯��발�ߍ�:R�e���".\6��v��	�=jU/!����-u�"]�$��a�|�����z]ّWV������_,�8�6K�1��w�}R��m�d�%��γ)�>�;
1��I��-�)��#v^���L?�����AS�
����z�M{��6�(Զ7h?6/m"!������Sz5�ئ��@:T��(S!7�ߥⰞ+�\��n���.~`؉,5L�Y�yL�yT��x\��	Ȥ����<�q!.Y�LBi��W�#aL�&Z��K�ޖ� O��:��o��a�u�z�+��
E5e�$�����=���;�j��WFԄV�y��r��ֲ�&�|F�60����O�QHbc��.5�M���%H�����������t@W�c݅�l�3��'��VV~���ޫ�c�����{	��[.����@�����TTZ�jd�TȀ'fa�D�v��-�Jr�ێh:�o7��գB|9�N���7rVay�H��C��q�2��o������;i��6:m����_'��\��vR�<Oޭ+��LEQ�����B����W�1d "�t���s�f��1�T�W��J�W#Ѣl�↕�����	���j�
�Jء��Ͽ*e��DþTt,3{]B�4�a>�[�9�3�S�����P�42�P�!�y��7��C����O�	��u�\��A	���3����H� (\Ľw��Ax�C$����3Fb�q��2 ���S����(I���'E��k�J_��"d�������_��@!q��.3���Fu�4ƍvwh�G����~���V?%C�q��lɿP�e��
��#pZ���GkaU`Ø��ɪ}CoeB�6����`F�=&�栯hWi�*O�{��7�O�A�
�A�0�7G����r#�p>����S��PH����J�l���*]�"����������
"i��<����Plݮ�h��כK��p���l�g\�`_G�ZD�aI�f*��J�آ����D�ʥ�}�d�
.r���3�%4�r"#�9ɴ��:{�Ǔ���[��;�5��N@)��=���=���j�T��<'��,��,K��~�B�CUr��A�,k�g%�-=�#5�aF��袧����*_5�y�#�iJ/%d#{�Y	��$>����0S���.���ɕT+�dU�	^�|��Z��R}���ڐ��{}�2L��x�N/�_`�������M�4P����_�q�J�]�~�9f-�m`ki`���#[�_��_n8|+����U+�pj��h��0�襹��	�L^+X���3�h��t�A��p��6���Sh��PPN��:=�F?󼼴�r�u�^�>:�+�6�e��2�5����:�I��4V&�&��J���Y' �k�%:�g�Y��Y�H4�}��~#��$���L?��-��GL�yHFT��7�>,��u*����<Y�eq�UA���@��j�q��z/�q(c�����@r��|�'��3"<;Vmf
_D��]xL�3P�q\b~�o�9���ʟɢ?��we}]�n>K�i0�x�.�֖�0'�LM�|�y���d	T/gmr���x[i�+���2�(��`����_�9g'�M�L+ѐ�Y�.��v�����U�%"c25�i�n�X8�"p��j
=��v�K޽�C���e��/�v'��.�B7��z�j�r5��2��
�:�UQ�0�O�>� ����b��_�Ȫ��J��V�;A���ȍ�us���l9&@�vSy�����ۇ�Ǳ%}M0�'͊��2��s
wY�f������=EN�\� 6�s�/K@=.1%1�"z$(\<�%�RW����=�����Oң7\{�l��jr�51�_��UY�,���de9Y`�J+�Q|����J%�[����,~χ�m���f%)���Wר��?��_�N��g=d����uj�aB�o�K=���г{�"v'3�,SkB9sT:t��/�mam��h?51d��(��#R���N�y��]�	�ݮl¡T��T�'Ŋ�¦��������.���P�7�9�U��@M��P�8f繎 "���.���uRN�L ���Ix.I[�|oy(�l��,�.&{��:��r5��z����A\t�h��ҥE�cy%�W�N
��h��GRa<UB�j�Lv�b��z}�����`w�mm���JNy�]��_���u$J�Y�{(_��05�X�FtC���Fa;I1�Y�j��x���V�n��S��5�V
��V@]�Bz�]r#3�^'�� .���}7雋�K����1S���
��1���&^^Q匨��g�ǧ5c��\��G0W7c�i��)PPZ��N�J���`t�����c�Q���L��a����֪���zÎZ��	���q��_<vXrŋ7���ư��~�lO ��Qu�o�ۮ���,�F��L��,
�SZ��ž�Q�w���m��o����{G�;�޽���2�4�(�U���us����	�5���_���dF{�إ�x����G!�R	U��><�H��$�x�� _��F �^:�y��1ܹ��>Գ<�����/��/*�&mòr�s2I��_'��`A���36�$h�&P�gs�0�^_���Z8~�ZU56!�"0�c�/'��.YE|��L�Yu~Y�0��)\�c��:a���j !�#�n"��=��7�ԹS�Ϡ��B77k����gr�e��&���ϟf"��44
 ���P���8��jg��%p"���Z(�da����@7����'Lu*�E:���MX�P��bU����L��r(�������Y!��0e��nb�͡�|�f�����ox�/o�.v��K��@X�O��{LN�q�Y%��~g47-�Ʊ&kj�U�	 Lqu0o�i��(�뚪��q\_q/�.��&p�=�)1�[�_q��X2:�YH!��7)���h��(	PK�_��ԟP��:=Q�E��[W�q����s��MO������m���iu����M��]h� dx@#����}�aɶ{���Ў̟�����N�"���re��i������JCp�sezG�go}]�ӂo�߹&y����h'�7��Ik���G�@�Q�O�1*uQ�*~E��IȜ�f�����w"��>���+j�*���Ӳ��w]%ψh,v��*��}�P����?v	��/
� ʞ	�M+�0�m�W:'�9OD��`(�4����W'{�cs9�[T��~�T"��+u��{]�o-�|� ���+�_�F2�w1;��}s���U�3�L/0EGHzr-Ȇ�R0�i{	~�j!��e��JV#�s��@e��$�8i�/̑��u��?-��:z��i`_��X�������H��[��p^y3��
�s+�ğ�F�'M��R���EM���yӅ֒�5�K�������_]�f�5�`��-�|]ԣP��d,Jl3�xuv>+����"����|η�UZ8B��Z������iv�
��`�!�3�똳�D��EA٫�{�v��Y�r2.[�ԠNI,H�Z�t�:�܀�l�Ѥ�J'/C����Vi�����9Ǥ9�%OT����lg
�~<��k������Ũ��Z���0ӎ'������#�>6��~�C��F?A�/[����e#G�#���4	�Q��y��3��o�4����K���#���嫝J���%[R8���s�c������d���Xsץ���K&�0�Ëx��'�!j�O���S��1 ̬�^khvd�`.��w�y�8��(N|E?N�p��N� �ui�O�J3sf�BF���Ӗ�:���P�� "!-0tAt�Mq��o�E��*�d1�r<�g�S�Uko����)���QF�Ŗ��^p��9��QG��{7�f�eN^e	[��^����D`T�p� ���ԣW�`[����|��A}U�#S� Be�,v��cN�N�M��?eL��`Y@��oE�r�|-�~�vh�"��	��oӀ��w����/�m��8����5[˟�4���S*��{��8�M�Q
��|�n %�ĉ�z-�`�����"�������G����\Ƀ���J�|O���'�xpBZ9���-tYnJ�m��d�����ĖM��V`:��aD*`����{�Z�%14��E�0[�d�Ƹ�SJ0F �^Ku-��	*��M����&�a���g��@�nm���y �C�Kk���j�={f\HOF�q_���Q�䳵}��N ���tz�iq���N�*�2�i=`�L���<��2���b���0
`� ܤ�>�cX�?�N��� (�g�Mu�p68�k��BV����n���|�J�|w�Y����	p4\��	�����X|{a	�3��K0�%�[2��׹<����rJ��cN�`�v[�4������U�XD��>r%�0h��~}�:�-�`�B�y
H��n.r{�DX��]ґ{��!0�~��z~��Da!W"��ô��|���~4t�Be����!�v�'e �!�S����4dj�Vj5�Gs{$��ل��s��8�È�Bcڂ�Fr�}�Y1��Z�����8
���ξ���#��Y�ϙS<F�P�E�Lz
�C�:�n��ȝ��(���8miZ�"��
�PYɂ���[���0\l��{�O��/;����l����O�{�tB�"�����|#�����+�����eX,��S[ǋ�y�"-�W�w_/%��7�*4P?�[$#C溲
>��8��i���f��+���|"G�등���!+�?�F�+����7�.��D)G����/:�@�!�N�%񝛻tg-�����1��.*eM�t�`��޴"�F��x��qp�#� o�����+cS��O,�938^RNIiq��ѻmM ���Ԅ�(	ل�䝱���Kx4��cvR~��-g�Zx���ԩ�����.�D�f�`��/��e��0(ך��(B[���a�p�%sS�#���:,G�+���]�a�Z�k�%���;5>ʼouJ�-�_�>}��{���kâ�N���}$@^�����)M�Y�_��a�\37W�EV"��[ ��"sÐ�PWL	c^�5�Z����O������[�!2*'�JЊ�q���q��gI��P�Z�Q��~�����SQ�+"E�6D�+�x��J���h�w����Sᦩ�A��Ǽ#B̃]]؁$��!Z����*�퍵���X����"';X�/�IW�́ϲ�Y}�=�ɪo��O�U�I�0��QG<�g���{���؞8� ���$]Z��l>������ը�~Ez�څE.�Z�ݯ��y��x����r8�CGq��OpW�?�$�g�
w��H;���&��(>iQb*.�PY�j�+�6Z�1��|�=\xP޾}���I�=�wT�QX0���)o�!!�������H`�2w��.�P|�Ӟ�u���Rz ?�Vk��ǮŨYޢ��|���J�d�7��R�"�@��R�|�C���K�����)��.��kb��A��^/۾\=9*���;^_�.�,j�(eoY>��7�g�����WTEj�O4˽���g~��כ1cL�^�9c�D9n��L(�.��X_���K�X@�&��/;�Vm��x1�. ]� S��`����0Z��c9��3�_��Ҹ��S�zF1ܑ�h{D���QY�=������+G���dr����]��������M�RN�>=�b������/K ���#�f��f!�`��RY�(!�� n�²f��u�ҵ�m���?�?7�P��D�H60���'1Z��
�%��b�˧ØEq<Lr�5��Y��:$[���|/"Ō��B�0���k+'��,9����̓L/�,�NڷVB*�'�R��ב%�[<7,�I����L����������6XⒼ+�q��[��_G2�i��K�gR��N� ����-�K��;�Eɭ��!���	��*0y_k�ۿ�y�-+�k2����o�j*)�������ܒ#>3��������ֈ�=	7��qm�gLa�O.����@:1{m�hO^�y�y��PE���g��Oi�9�x�z�b��������	�v@�:���0���V�R��������f��(��ߜ`d"��x��2��|0a�-G�����dI,���0��:}s��ҳx���GVY)g+�*� I���S��\T���5s�O�=�wJԑ�3���5�
����ɡ���	S���c��Ft��P��3��	���V�3�o��bM��8����o���wP^$E�1�8���Kx�����*���w��JO�Ux�쯜�o�RB>�������I���:�l&�c����YЄ3�5������$�8��U_#�H�;�2Y��8�#��f�	���r��IT�B�JƲDNE�x����9�"8��[�Q7�&�i��� �!Pr@%^2�u�K$ m}[�4�j�a�Z]��h�a^�������$Ca����Y\�����a�������)� � ]��p����n����&J�>�*�J�3�c���E�gT���cby�m�nC��aaO-�.����.�a��3�������d�E.�@���B��\jU8Oc�X�q��Ţ͇5��9����;[����=Ŧ0��X�β��N\��G�]qRQI6e�^��#[a���N��[g�c�ꍝ%����c���.a8 -{��N�5[�����QS�P��o9��+��/�2�J/�!�@���a�Vj�@(31}��@>�x1��|ON8��T���.�2�$3
�tN�̈́d�sâ�8)�\*?���~��-�1$���2;l���:�}F��.E�m�B7�0���ԻWE�Yk��
4#�'�a�^R�z�ʺ���kU�]�%�)p�t�,5jԙ�Z?J0%R�C�s�g�Fd�YtI��U�̦M6� ���8��'�t�ď���'^�!��Mu_�,Ri)���$�Z�9�؎�w���H�����}Ci��u�,%��K(S;�?��Jd17ⱼ��54��"E�Õ�Hw�r?E��Ǜ���y����r0����m��k���Ý�5e�oA�o��@�`F�5f�����[�;������In-��ڿ��Ny��lm�C&ES��H\<�AA�JV�Mt��7?�s'�U���hHey�o<v{c�=�S��{�;^�R��T�u�Ud����^�q\�&��N�#�>�bƙG��pB�������$�?>�"d˯��R��t����'� 
s��5�J��b��f^�o�Gﳡ�@�qC:ۻ�����>��$����:\�x^sL^4��C]���d�^�}�~�
�-�W@d��[���E��q���_z��Uвs���<K�Ν�tx,B��?��87�	B,g-����o���(�z���%���L_�360cn�i $���:0¯=�Q��H�ȯF���kg� �5�F�Q�tG0*/�)��1(l���lh`9��n����=����Z �xd����̭��F E�������G�����T�as���^v�1l��x��Wbu+�'6��Fi-�H4�Ӑ}�U���a;8ٽ/�PBɸX�A4D0ds��/��d�ɣ�\�g�(~bWu-ұ��967WP�yiL'������\Z1ȤI�aGÜH�q4+���>����*@�QS&P-k�sr�S{��X��!_~e�+��2�տ�+V���6P����:y9u1;����̧3ru���Z2~Ig
F�O�x^�F�L+�U>v�5�:q��qz�}�:�� ڰU���@C��La�}�	B�Ud��x��f|���H�{�O�x!l�o��BOn� ���S�32L�y�0c�/����:�M�;��fK�o3G �I��7�&��pz��R�qtՐ��zK�iU�K�/Qm9��?Y�zJ�Q?Qm?�ehB���-�������`P�l)¿�g��ST�f�N~LmU��r:2��&ʭ�E���Cs�k�N�~ݺ��2��C92���0˛&�fCUn��Z�w����֤U߁[
�����k
H6	"��ہ5����
3��^��a�/�2|lM��^�x=9&e�%<�[��1s[�Lt��Q�:���Ð*Xu�T ��IO�߂���3*�5_�W� 7�E� �[�7�ፒ��Q��3.�������H���sU)s���<[T�:q�z#چV��Y�����2y�� ��1�&�l�����$�����gǻ��t]#?9_k7i�~������`!CV��Gl�aAS�J;�����u�+�a�wW�{׎�B:��{�&[5�*!h�L5�pDc�:�qG����V�[�د?�!%���6D�S-�7�q-q���D4��v�_������H`����`��؟SQH��S��8'��G�����f(��K��+�L�睾[8�ӡ���^f*���@�����q�;��o�Ut�+�*�Y��xA\:�+��b&��������^�"�N|���֔��ΓWf��g���
9x+��"{������N��2Ȼ����<���:m�.�!pF�C���J�R+��Jߩ��q��š�����H��|e���I�J,��b�_�W����?M�q;ǘ~
v�I�`�0���YX�cBD��u�a�����(U�I��"�F�N-��Ʈ+��,9�s���V�|�\*f^��q�.����G����z_��*���a��o�q���P"��u{�@� sd6�Y^�M31�[8z�xĀ���CDZ�+_�T��rҠ�=S��O�<��s�i%7�Eu���ȷ�6��8�c���A�	���(��3�V6�.�Y%u��,F��D� 8F��T�q�RJ\��X����Dx��N�#����DF�������o��YXc��&�݅������S"Ț\���6�e��2My�,�X��F������,�>��nN��Ѿ@����q�����M��6���u�����С"\U2�t��y�A8��W�i�?U�+�C�Z������LL/ُ���	0g�K��ҡ��r�(�/P?����$Ղ��f�ok���;��He|d+�;���ܜBV�qQ��� �<u���ې�����&d�4yd��Ч%e�X�:� �	^έ��u%�.����$��afg�`;�chP��ek���w�3j�tЭ��~���V��&���L���Ɲ�`D}�����Y��?���<)b0b��r�9d�?U-�ikR>���ۆߏ�Mn<an��B�4��������L�ʁ��h~��q������L2����~b�#tCu�'��캨�ѱ�%?��,Ƅ�%E>p��;���'\75��a{b��1�!�t���r�נ��%?�}���QI0���d.��l�v��"���P�r瀮	�L$w8�!a��{�P�����㮿�|�N7�'ݽVVx��ʪn�5���3��;�噩y:�Ch�{���ĺ���#MP���Z�e��C�D<���SY9m�a�+g��ۖ�8�9���[��~=����w-��)�[���|x��L^�n)�po�a߬�B�g��Gٯ��v�H*>I�5����� �ýL��U���*�:ā�*�=�r��'q�P���1G`�2J�['�pmp#�E��at�.��ʵj-� >��[i��l�a`ዜau2-� ���=缦�T@����UuK��P�v��:�0!6+��^��|_�#�?AO�	�n�Q;�=��I�y�x����*%���E)8��<ˡ�A�=yn��]C	��A8#Efb�,�h�
K�kO>*��89q�XE�`�ȈP8��i�Q��٦4�������+N�����e���E��� =#�W�aMC�XI�0f<����rAxh����?a��>)���l��nd���?��|��a��r��l���)vt�
�Z���/�C��������i7�mv��r�;1uH��5���$��ص�}j��6�B#0�}y��\&��N'�f���Ӳ���/�L�(��TdA�w�7�IT�/ep�6�+�^����Q!�5�R�w�.�Չ`�19o˨n0p��p5=��"H�訌@}�����g,V�/��e��NuAf��%u�厔T��3�ch��̲ �Y|1�(�(ZC��ĸ$�e�p�q�q�4�@�n��l���_�k� �4�c�w�yCJs����Jw��UQ�;[���L�#e���ligm
����&X�i���-#���&X���qЁ&��L��Ĳ;AŠ$Y:��`\tOb�#��T3��7��{����bP,�ey-��(���D_����z�+½�h:?3�t=����uE:��gcj�,����b�$G���w�x8���
0��b���S�Gi��A�$Ʌ�1#K�w<g���n%S���FV�AF��S�ʸϳ��vC�V����_����d�}��c������W$�M�~?��������
İ3���Kp���\䯜#��JkurЦ�n5�/���̅�!�[�vA��������~�PF)�'p�	��4�?r����8�wi�{�p��Ȥ�f_���d�X�j����a�������ߡة'��;���/㐵VC�S���?n�(���T)w�T�OC�����P�\�A'欚�"0�7���l�S`}ՔP��\��G��b��>��_��0DS��{�{�R�h���ޙ�,��{��u�H.��O֠��%=��"4U%�K\6��r:(�bg?��U��г��df��x�r̬�|��5{ܗ�,p����.[ "RŨ���6޼{��i&�ҋ��h!��П�2U^˄�X���G`�ъH�a����yn����%��R��4U!��� sĖ����s�5&O8����Z��ڨ&�,c��+�޴Uu}X�\m��ǩJ7��V_g��3�0�i4���5�C�J��R��U�Q&X��P4W�</hֱ��x	�ʂE=�f�҆���Hd簇'��YfY���a��"��`�ȐPv�L0��<��Ge�7�(Kt9��U�����!�7Y�T:g��\Y�~#�RHÔ�QU��1u��Ɗ��|Bԙ��&�;(�P\-.���Le�� F�IL��+' jL�;��`*lJ��ZD�_︥��6�{��#����F)�����-��f�=���!u�%�p嚯
���	׫����mW�j� ���ޥ�V����	�	�;KlҤ!
�N���FJ�4���S3K�̨o���y����<������'嵤à���Q�#߷Z̴K�}R{h�p�j觏$�� ����O�����][q|�#��}���j)*��F�r�,�7��w�K��Y����\�h� )�v�Ic�$a�T��������'W��I��)X��m7��2B���b�R2�8�h��z<����o`���}FF����k	�T��rĘ�>�Č1��:��Fr7v*�x�8�\Lָ�cu��sz�9��0/8wj����c�M/��'�ƛ��^{�/;s�F�6�I.ŷd�h䜼�:]�����\̳ۢt�ֆ�9��0���ZZ�Qv����b�(nCʠ�/V�m�7�����9
gil|��G(���שsV����W��Ǻ�g:	� �^8�ۆȘJTY��[�Ws����_�~��;�.��	nm�ɬJ��5z��T5��W���d��q�����U�������:
��,���+�qc�;��!�?ƭ�8jS}�u��`�`s{Da� N��AS�3S��3�z����4���),G7LZ����	���+;K!%Y�<��}���Ic���G���m��sT�Q>%��m��5ql�2�ץ�\�KHް��	S����bm{�A	�x�=q雚IZLz1Z�#m����Dd��b:S�u�Yi��_L�� q\��������$��/�����7=dY�k�'v���4߲ ϴw��4/��07�(�>s5�#h�g���L��5�9;:�~��Uy]�u1Fm��0�.�����ͬ���O��w]�4�����>7�:7x�2��֘R�}3��ygʉ7��!��U�x_#(R�!nAd�0����eڨ|�&�p:q9qYG��:K���(��T?
˚�k��a��q�*�;c؃٣�חH LUjg����:��
��\$U�!�Lp+�U2M	WB�V���!��*k��
�� O����7�7}<�%$��@ÎEYr���~mǧ���sG�;Wͭ����o-Ӣ��[�(�G�B�b�r\�D~�m��JU������L7����7��eB�gu �)�8�q����e������7�.@`�ET�P�4|m�_�s�h��:�WoADaX96�X�	ؚ]G�Lk%�)>�(���43�N��z��i�,ko�s{J}��zH���}#3��gȷ��[R0�`e��b���3�5S2�#�SG��;I\�N��d��w��恘�$1�lA����h��a�ܺ���u[���X<q���$zU�{��m���Wқ���ܗ�U���z���m�Y���Z#�a�8'+�� Y(��p��Ō~fK��S���~�B�O,P��Hǚ=8��H4��z�h �����*B��P��ڎc`��j��5W�MA�HP�3�*��f��E��dW@?*��g�X���Ϝ�����(�D�Ղ��J��7�L0��z��Ŧ0X$ig;f.p���=������2A��YB��zs�1���,�i�F���IG�jcgi���x��t{�B,Vz�\�Q�> 
Q�oW�טeF^r()S�D�	�����F�9�)`~����fՁ����ښ�Y��A��ȣ	�E�;��1[ꬮ�Q��\� �c��;a�ީ��!������R��A%Ш���e������VHo�s|���a��́p$M�T����Z۷tYs�e}��1Xa¨٭ѥ�#:Ԍ�������T����[�=Utd���fZ�]��dr�����YKw;kkޓ�o�p�������}z�j&G���Sm�~o'�������EE��k9b΋���b�&HE;M`M�2H�Vm���	���>?&j6H�� �#�;�^��N(�c�E,�˲������~�K���9��9�W6}�/��t��W\vO<\h�#��I`kf��3�������w��v)�@>m��}Z�>�3��,�p��lR����/Q`cᮻm�X�2��]������8{��sG��\�tQ���R��(�h�~XX���[�U�b���Gv'*.n����h*G�J��?��{*�(`���S����>`pRi
�ؙ��_Sgi��2���e��/���9�Q/խ(���K�A\#�L��۽����]]k��Z��ЗR�i�Ѻ�7Mm����� 8���}�&�G:E,��ow78��FP�&��h�ר����1�y�k��|�h��xP������'K��߅.�;ȅ`�>��0&}vH�0JW�5�U�HTYbY,��
�u�u�(�Ae>�a��ˮ׿n�&�q[U��%�c��V~�umֿ��U�3�Uf��Q�����kyͶ�׵��I�-��j��T��B��;��݊��m��_yF���7�.����ţ�8��yn��]�X��6��M��|�rM�e �m�~�I�"[M�)ρצ0�c��l~�d�(#dS;`���9�/7:�73�NM|:7�8�:����s5d,ν�Ň��J�p>V)gn��P��Δs�0�ВT����:p�o�_U�e�Km��>OlD�Z�Zs�Km�çYu����Y��ZS�i}\w��r&�;�}�X�u���W�A�S��ax�Xn'�F^�bt?�d��7��s<7x�x7�s�R|��ܮAP�ނ�S���� ���M+��*�:>K��Pz�{]D��2��q<��O`�'��
A��3��:$t&��XKl%\�N;T�dg�(��"O܇��� �u��b����?l�V<���-3����E2�lF���C*�/���}�A��F�5����gR�'���w�dI8�f8��?r%��ß���u�V���,I�r��Ċ�4f�E�m�F���e[�� >|���V&~y��׫c�)�N˛L�*���w-b��=����p��6�5!1���j�K5�+k2���}!&$��PhDx?+�6�&�y�~]E�t�N��[��OCv�9���\�Yp�TMh����h�`�%?�sJrZ��-�ֽ~�G_� i�l���Հ9k.��qZ�b���$Mfo$�Қ���d�ފN�=�r���=����98 �4�#T��	cJމ=���[���n�|����������i�{�6D*��i����U�����jGh�&W��ז��t�5�3�q��$Y깺ʍN�{�%��3zF@?O�z#�\n���u��d{���9�K$�v���Q���ˬP�P;���ܮ���.�A�4�_�C�֋�5
IH���-$�e��V�K�(��"� ���j���9���G��$����Bo�ɹ���H[>QT��'�O6wLׇ��͋��W,��{%GK�وN;y��<JB���Q#諾���g�����iMee��s]�tv���`��9(X��]�놗��&wk(�k��7C���"���jKϵ7��E�&��k ���l�����i�5�Y �eU��|V��T�<)�u#�p�p�t҃B.!['<Q{�3!��$=Qd�OҜ�a�o{��e��]<)�Q��j�
�l�����F����gϚ���OK2��F�E�X��;qE��RAEO�e�hLgq	K�/�!��~��`����S��'R�$�n��\�I|���4��{-V�#
����z��k�XY���8?ϳ(I˛Ñpo�" %쎼�HN��n2�pk�o��)f��[p� �Ss{����}����̪�]��A:�� O�"S�&!�K'�O� ̐�.�V3�мu&W��RDT�U��'�� ����:��h��jH� �}W�q�~K��8t�оR�?Zwe���}��H��q�4��Z�[\n_&ɼ��ițE$�8��[�j�|�����bc���CRɆTb*�A�$��)Gj�`����6�j�uxd�K��	��aٙ��Ϫ+�ޏ��j���ʢ���Ϳx�#]�P�}��o�Ds�2gT��g��P5�^�^��͒m�{�J�?}�ɣzv�����t>��o��Ρ�BК���}�5%�4Bx�G��(:2�������7 �Æ�3M��"��O�)�r�����w�/�<�-��>L=���b�y4�p^G�U[�r� �qy��=�YAp��f�b$��`h(�p��Z�>�W|�9�fn�Oi�W������K�g�$礚^nW	)MsL���x�i`�"l��G8��N��B��j������?�9�Lb������L��[-�44����oLQ���y\f���l�
���Y���s������"[T��ǧ�J��%��
������{S4p�x4����a�AZ�P��a�Ӑ>�X-��Q��-�;0+{=� �N�uy�g��]S��8@S�""��~��d�>����E��@��Cj�ǈ�F? i
��M%!��1�.9��Q렺��-�.v?�@X�y�;_y�G�}5h��S�_\C���+Y-�_�f*e�,,DlC)�rT�`���y��28��Im��'& �8�(�O�����F���1��)��4v/e�s~���ݣ<�ppy:���ed�q�OH#�T\"�`A��� �@S�SpN���[�I�K�����#wϧ���UVw�[�D�?N#0M�H�h��vE%���q��h@	� Tk��QZJE#}MJF�W����	)2�}Uq|.����<��c vyb�|:�_��#�%\����U� Y���F�f���,�J�/1/�=&�5���!�
eő�r�i�x�p!�wJ}����ed� T�+c`�k\�Tg�`*�&]|�}~rO��פ�'fm��B�>�;�"[@�������~èu#/���h!}����xi�b5H`��8@�� I�X�e_J?6���o�B��/'BУZ�-�Bڥ����8]i�B�tlP��=��x�z*���Xd�~� K���OZ4s\W�O��(�Ł�#�ˡRLA�cc?3k�L���f�	��V��+G���@�,�?Lڍ��n&�<>^�}��RStM$�Z���_�zTgtwt�C��L�b�m�B%}�v�� t��$j �o�8R+X����b�, Ҡ�����S0E�:��[����Qs5�����7���V/ԁ����u�y��z��k���r �fp��G��'�k8�W��'�0!c�C�#SA���;�^�|g�ʩ��xV�A�rrN������~vm�T�$��'�^�paً����k��ǯ��Hx���j|�����8W��!U,��E��s4׋�2Bi�������ҁ�[�a�����dՃ����w����t�}��9�$�M��u�ӵ���zg��>�!e�����
���1�/�OI6&0�\�T)�_�ibY��y� rF>����}(9;	V��N���{0�+&g�d�nO5����g5�3�ϔ(���b�EU��Q�j�_{�ӔN݈d��
��w1�KLZAgj��%���	vcG����%ڿ�ԍ�h�E�v��

���S~�E�E�J�U�(.%��[�!C݇�b�Wn�Ez�_�շ�#Z}����c�j�-�	�b�M�� ,����-�.�/r��сD77�:��<�1�y%�?o��첰�0[�2�3J&80f&H�x\֤J|��ّ�"*c>�69d�j4�VT&���x���愐�_ /0�˄�OI�Ő"o� ��@��~4���	�#���`��V*@�>�.��VC�V��,�?V�<!E�lA�A�7�yi��Uj��m�M���2����(����&G&G��V�I��|B�<º���%?�K��+Ȧl�t'�kM�Z�J閗|����h�bb���"�g\Y�*z�K{N�����!��x{R������J��Lp�7	��C��r�S��)�<m?�fK�k@��_F�X_���/�g-����vO�Ds���'��sg��W��������ȉHL�N�3�i�}'�S?�.)j�����Z9�3�:��"��q����5�^=�����f���줧@�Egם�xݭ�Tu%�U6�e�*J�SeÛR$����/�dD���|�mZ��mH�_b���ԫ>*�H�{S??�ͳ$7����ƻ�En�����ܰ��&�����z�q��u�e��ì��c��4)��״M���ۗ��Ql�=�pMi��zȆ��1���5���.�yh;[,� }��+QV�Rn1a΁�pL�U������PG�<���&'L�b�y'�����VK����4�Hw��_p c���B����$��H��R��&��8�4�˖��x-�1w���G��>q��"����tl�r�=�7'�'Fc�RI祯ח�*�Ǯ��H�aէ©pZ����ON�r���~aVy,'8 X��@�d �z� 3�f�1`�!��	�l�:�*�&ĵΝ�L�%�ƚ0�C�p���2��x��Hy �s7����(�Oe1���%���=�AW\$����J�[� ŗ�R�MNu'�#��J�K4*s�*X�eыQh�Z���}%�5.-:=�"F���$UAx&�fj���eX���5E'�_?ȳU �^���7�쳆G�%��*Z0�yq��_\������!R�0�yV�3��R5m��Mx�27��jׄ덪М��F@x�����D����敺�:� ��gN�_Y�Fg�)J�!����qK�`�d�Xǰ��\9�~5�uD�D�d�j�C�7�nOb��U��ΰ�朶M�F�B�B�b�=��xB�AC���X�z�~�?Fa�6&]�1�C�P����?��˱!��yH���ۖ:E�nV�$��������5Ye��~o~��7	g"zp��V���[���5��|�Tӑ�Zj^L�1��6�7�*^Z�#��{���#%Ǎ��N#��Eʦ�F�~b,Eٕ��JUsx	nȕ�v���wI
\�V��VOP��ɀ�ï�ȁ[QB�	=6U�AϮ{�W��)�Ǜ�>�ٓJ����핀_O0�'�>�!>���U��9��O	7#��ܲ�"F}�GB%O}-�A�w��3-͓����:���׀h]��b�/�1�"*���#� �J��ɴ���n�PC���8;B��01�Iú�K�9^&?>�O�r��/�䢧P��:d�q���7r@$
���E�VoTm0��4��ݖB���/��e�?�ߒ۲3���C��_�׶�QM�팮)6�=�\l^�R�H3��i��������Oa�.�e�W��?đ]�.��Hu[��J�
���l.UɄ�G��>����g��z�2D���2�E�5�W!��۶��5�n
-eC������o�ğ<z�8zWu�T�ԧ#�-���n@U�9� �sV����<�9hB���H���/1����������ܓa��G�"�������=�!*�6uބ��PY�ύm	l��|*�M����D/\g�a-��F�n�y�ѽ�eM�v�11)�>P��<e
�nW����� ;$ƌxݰJ$�N<��l�g��}=��~��H<�	�(P�˳[�#I�ȳ|Y�@��aݫ�!+���Ԉ33��s"�[a�հ�Jq(�{�ڑ�9~C:�t��5�J���V(,P�Zz�f)��{^��G<;ԋ�1���'�c����S;}3�����V��@��yv��5J>i�Øl�|Fg��!JE�C��y��,�;%I�����|ˢ�i]`������>��[i��0�@^˲j ��a�J�3�+��i���|�rt-F|�z�.9�!�_�P��z�BL����3u�s�.r�T �4��*������kp7Ć������ r���|vݞ�Ӎ����-e�5NP��2�()�WN�1�c8�Q%�:t�eB��*��-Kn|�u=��/c��9�jЛi2���#I��ꕫ�o���j�V�hl��A���h�o�}|�O_)�.�8�q۠@�d2^�c��po��Z���o~8*Y�a$p�)��J���m�R�=_�U���T�eZ�{���xn�xD�o#Vd��R�7lU6i�xaE�1ߐm����ҽ�)����'� �+[$��J�OL��)��Eĥ�>���q���Hk���N� ��0\�Z�����d�ͅ���p!�Ҝ9Q}'r�BYs� qd���C6�}\�Y3ہ�}}���S��~���rt��OA��-�<U�| ��I�RϬ"/�4l�L<}^�;�V��.h�8�սw+� L����I'���j��w\�0FM8������b���7��D�sT�.�z�1w�=�bO��F��ȯc�	?�"i{OǴ�$�ڎ,��(�ڀv��=p�& �UI��uq����Ӑ�D1z�6��-�"�!M�T��e�=�<j��Ao@�i����1�7�d�i��Iu���g�!�@��s��%�|�Bb��1P�~�N�-��V�9J�A_XCY���zM'�Z�Ȩ���z��� ����ֶ��s���Ր�T7������4k�F-� fR&���Zd�U
�aP���^�����q�Ʌ���?|�,5�m��pB�y�01�T=�s�+-XbUw�����\{�,��0�+ӥ*�'�H,�b���� �� �$��Y����cHm�� u�),,_O��Ջ��m�y:��P�?c�����Ō�,��#l>,�{T����j�}�1^v�������3�J!�B���-
���\n^� �׷D��T6Ă���e+���`[=��w�4�xI޼֋���6x���HcEL�6�Fڐ�o`�1��uo�:>�>LUB��i��$�� �4d���tml�	Z���ԭ(S{9U�]�Z<��&�1�\���+�~�%�C��L��|���:�����I�D�Ob�sk����?6��2cn�oHS�Ĉ@H�	0F�x(^��m�"�w��s�%	h��&�R�ݫY���=	Dyr)c���:W<�*�.X��WE٤�?b�ߐ�{��5԰�<�Y������Bvѷx�7����������9J���M�Y}+�"d�nU��A{oLBp�^�1�<�	�cf�`o��.���/�)^�UZ�7#��moI7�f ��5�b%�߱Բ�W��qa
��8�k,Qd �}WLY{��:���Ȇ��~8x���
�'�C�\�5f�Q[n���t@\3<�>n��wU}6RI���x�����g��1�~�+Bi�+NE�jVc敃��ށ����T���A�d�n,�t�����1���?d"z2��c�&��b9�<�_��oh�L6t��I0�����1�2���Xm)�6�R(�ax�ͦq 'K�:aF�6d�	7�!����:�����~xxF�J=��Wϧ���^�x��F�-['�h �Cqi�J���/�K)�҇R����'��XrЅ�0�� /?�+���F�f���V>/���73r�~ �^G�l���>�Ht��U#��	ā�>�#�u w|`ܵ�΃h�A?�=u)���)����a��Ȑ �D��������J2ӦX����jM_�~��� V�R��1�s+�A�lu����K��<��*����݂d�<����ë1���LR-#z��Fǀ[��0�c�j$�0A \bߙ�Yhy
���v{KzH���vCE�/�#_� Ư���Vm�Yq(�!����t�aJ~�\����z���v��t�����qG[���ڦo��M2��H��1��V�����3]��@��&>ئ�К�Y;��K��h�ځU������[��<��D���ѶB2l�	��%�f`!�7%W�9�F�������kF"ʘ��5���K���V��"h?$]�M��8K�8��	���bZ&�?֠b�!̱Nv��$�	�����/�E�ُ��P�����U�O�-��!Zӧ�=&�d]�c	.����Z���3Cs�E���Js��'H��$���о	�!�3�jǵE}bw�r������Ó^n!���g@�".j|��c�^6i�58F6����b��ƂOS�j�UvRi��i�����2�a��1���F��04��&�������Ie�=�q!���y�}r����=�B�~�D�;!��Z}���$_����~���UO��K	�XҌ[moe�`�2��l���H�`�
��HZG̜�E�p'����\*{o�aIKl�Ļ�	���Y�s9�͹}Sw�����ʦ7����di`Q�fG�j��皮0�f�=r0E}��V�c��#�M�J[�� ���Z�9®V�����6@R��E���M�fZ2��6��ڛ@�>-,���π����K����k	"���4/G����oB���K��z�*�K5��'�/趒�޻ �T�c����}�`��e׬�q��0a���U_����ߌ���e��ҭ*r�P����哩j�Iv���RDq_2��cdD<$���˙b�3�ٜH��L�|��
k����U�n[�kب��4������1[�q�U��u��A��xҳUÖ��L�������/����<&����kԐ���7	�?��8ǋf�YL�i
��*D�YT�jhm�6�s�CL��+H3��!�m*�3��g�ߖ��!́�h�큌�[�t�X���ф�!�{�T~�}5���ī�?~�z��	��{$�ҏ�0�?(+��Ez�݀)�%"� �.n��\�L�q��&�qT���i'�^	��K�g����9��D�0\�U���HTL��ns��{Ip�Z����e�^j-�q�7ۺ<V�q�8M=2xA���9�
7ˇA�។7|�te4�d�t4���o��p��8|$J�/©��3�mas�&�7�P�2��Ύ���n{1�#�Q�.��v�#�k�O����� O{�KpD���6>�v�T��s���#Z�5,���+	g��:4B^�Ɗ� �<�~�+DEȿ�%h%�u����vB��9]7�tɧA'q�AjP�Î�3�+��|���?0��X�M\b.�{\#�/�X�9�X ^�'�i�Xw��ցz�X�[ah��� ��Ab��$e�F����q�B���T����{B�"|'� ��#0������#���j��d^P%\���g�:	���$1�P�������g P�@D9��&�AU�;�z�*�T��A��6��ܧ~��{���r��/ ﵐ-�@M�8I�=����R��/���BaA�>%@U���=-�HJt���X�v�Ƚ��dCh�V��8�Y�Kyńjt�kY:��|���Oi�Vzj��q��G�;i��5*�5�0��Y?��jbB�MrD��K���j�����t��e����k�!f�e�Qy�&U(T���&��O���ʈRK��N�u�yf�(�����=a��yS�Ѯծ#�oG.�t���*�p�~p׌��/ξ!-�c��P��ۀF �]�|"�84	 ?��q>���NO���1/r�5:nV�� T�*���;�U=}Hޜ@ ��bB��-]đ��ʥGb"�Є�M��NV��*~���1������sf�1�����ZS	��Z ��D����	˜����f7�E�U,���ZM{a�->B��T���
1�+�+,[Z�y��~�����v8�z!�\�E��󽕗){)d5j����Ε�Ǣ�QJ?BU	2�@7i Wˍ�B���� �1��d�4b[��f-����k}G�H#�D� s?�_�r���	��Ǯ�P���@��>�V���$K��mw{g}��Z�ޯ؋��Pz�`%?C��u�9��|���]#x���p�)�O�z�D-�����)�Ϸ�-��I�4�$KA%lE�IB��1����%w��Db!��b�uĉN�d��<�h^�H*��Q�<��"���`������G���� �P~�5뺇}B�{[�f���n�t��Ѩ�����n'ɚ��"i���?ʪX"vR�Ga#�?����@V(B�38��Z��jt�in�xk%l�`-�oشf{�Mmbt���B���M�L��h��B8�[�;މd-�]�J�]�'�3:Q��\�$�t᫟�< ����^�Ϛ�f��x��+]���
�9y��Id�f�00��ѣ�ȭ��YՁ�.�G@�(�����Z��!Nk�a��)�k�,���I��2/��S���)��J=�����������w�sy�#*ֵ����%c��B��Z�p�A�ۆs�D�w�����v+k�~�^������K>��g�E�
�F�s1ą���(
��u��$@s�Fצߓ����	9���V����Ջ㈻�)�N��ۦ����CBEU��#+[EN\ƾyB�; [8���3A>Q��e)����k3���G�S��%����j��u̧z�z=t�w��'�e\ z`��t�"�v��l>3Q�kXCͿ�,1y�=�#J/D��X��H�%2�
�h�WX�H�e�g*�[�4�BrE��]�A5� ��C�-�IP�	m���E����hXD�,>����jb�l���Q�B����?E��#�R||�J;�E-&�bI
b�U"��uU;�	�~�w<�n!����0Ƽ@�����1��-.M=��,�1Ԟ($-�:��4ނ�[(���s���]q0A�͈I*a�r�k��v	�˸]F�O���f۞��[����Bڊ2+~���5��qP��3p0�M���? �f�����vH4:�U9j/!�Z<
��I8�����d5��c
!T�J��U<����-�-�F�7��׀��i�B6���i�|���0=׬�\H%�0�xDD'��������#<�/�(L��g0#6I%{�O�;>h����`���^���N�%P_n�߸U��)�t��~��q�0k&�'�W�hQ�Ot����u}�zǬ����P��^ف�\�)�|�1�H�v_)����Oݼ/y2bL�Q��&,���M��
����e"���?�A�;37��HbmK�.y~��&T9�f���Nb�=a��"�<���9aQ����]�$X�P�����%�[��ܫ�����`Ĳ����ZY:A�D���B����q�v�M�=�:\�`:���Ij��؛�F��V��<���NiO�Nȏ΢�<niz��`#�L}��@�Ǳ��������@���²�Ua���H/�}.�(G/s���W�i�ЈS�49�a&�cM��x���6NS@�m��3��|~�6(������㼘;�N���iz�Yu��t+X��ͫ��U����<	�cIZ�H�UK�!�����(-�p����HY	b�������(2�G�l�Z���	n���IJp��Xejߚ��7��˹�r7����Yt{Jxq��Ǉm�-�;Ґw� C:�_{/�u2�����=�o\�*pv4�Ce;�H6��
���9mϻj�=��J������f���Ϭ<�^@��oM������7�c�^����[n�����PG � .Q]O�
�s��P�{i�@�<���q_�H�Z?d��߮j�eDB�k�W��>@XT6	=���N�$��=G�rC����o]��z}��mj
4���qL�YY��	��=�g�D�\�ڻ����c�nװ�lݖ⴪j�JM���OK��AI��I�/ �]�*�S%���6>�l6?�55xA�O��F�bי���m 6�^@�M���Ƶ�h����?*�?P>�����B�[6WT�d����E��u�y�}Lˮ� p�Qx����,�v��E�W1҄��į��V�W3�l��` ��P*;E�J�'0!xVα~Lm�4�^�ui��h}��o���#����S�Q&���}=���:Kn���QN�:�02P7����႙�����a�u��^H=-�p��
��|>[1�Z�Y���.`9v]ǩ���������/Ѐ�����^�D�u��P���V�gK���&yCW%�@3��Ƀ]F���$#rDf��IL���[XR��.�1�v��өf>�x/�`,6��5�=N֞��'��@��W��S�����U��4���o?�Raf�A�-�r��C �nU�
�6�ٝ���i�,J�ɱk�Qg�myqJ0h�Q�jfq�=Lm���O$u���G�i����Ķ�s;��j��OJ�d[�]��W��O�Y�Ki�5�l�qZl�>��|�b�
z�aS�cȉ��0�F��&4���弦���V��|��?��}��z�A^����2��.��a�(�X�0ԖН��Tx�7�)PL��M@�ĐVc���J�r�<w��C[1Ӿ�W�- v쀴
$u{�Z@���aJ��KH��
��M7����e����JS.*v�LK.�=E�\�[#sc�/��,Kh�H�b�Mǣ"gO��_�l� r���(���r�A_Je��>��Q!R�1B%gj$�b� {B<d���I��s�H�L���ޥe22�-�8l�,[M�h,�IFM�=��r��k٣Ӌ���Y�Z�ل�WA|����w��w����!���c��Y��lh��u�;�m�┸���P˻{*�����b&1l67�7:��g��G@Q������7�i��l������K`��t����R�������^5����haj�]yi��u鬐0?Wv����k���x�X&����u�B�4G����j�J��G����[8bA�u�ү�U��l� O��*�T��O�����/X<���,f=��.|��T�vxD�-u��GFBYmD��Ko[�[@��	XB	C�"ZPD��xs�DF�~G�����-�@� ��&1����w�|P���ɞXw�"�6���ąk���a����	2[^�
���ךY5�^�����	����r�Һ�y��>�S��Q��rj�j8]�2M��Gh����(5`D�|?�>�����=�fCq�UyD�������ߵ&k��NeaJ�k���)Y���F|$�l���n�����9Yet-�#��þ�g�l����Ҟ
���ڶQ��XD��%��WtJ�S�S�֗�V7�ό?�6^��u,�~�4
B_�qőm;o܅	�Eqxx��w�6
4�����g)��e�bk�����BH��=�Oe%�
�:�Sם�o��>�Ur�_GF��y�"꺤ҝs	p�%M��7����m+��z��c"�l����e;gleW����>k��ݶR�<7A�������#d�ߍ��d�}��ϔØ��[�<��d�{*�v���#J����� ��p��^^jSm��!�ƇZ�G�#�q�s6���	Q��ȓ`���� ��G��>c:t;uLv�S�$Y�_�fԷ�w�h��\��泬�_�����= 鬙��3 ���`	��N����v���o"c�0�jȬ�wk�P�HB�/��Aݞ�ÁZ��y�����=����颤Y�*U����g^�?@N��W�HJj8~�)�<8z>�ɤ�V­M���{�U�J��u+U\.O0͹�,��V< t;P�� K�L�|�=�+�r���;�76�{��S��B�&ST���x_���:������&c�0�B|e������Ʀ���b}7�����k�1JН\�Q��t?�̛���E ���@V�1�C>�|����_�It�8����ǃ��^J�}%Xo��}]a�+@F�}�;�\�2��P�Om $�/}eY���ȟ��Cg)��we�7cJ�0�kq�W?V�)����I�a3��j��yC��6Df�W��PIw@֤�SN�}i~wz9,-BV�Z��6�ѕ�P::e�p�O�v�ũ
�y�Uf-��᫵��Z�O�|ݶ�5=�͛�?7K3P\�(9둭�y�!��^��pV8D��qs��u|�I���$ �U{�����h�1��DP�)4��I̡���P��z��!d����T��O�E\����Y���k�v! K��^D�>D�0��eH�C��R���H]~���M���(2//�Ƴ!S�~�����\�0��^�s�"�"}�*�'}h̑,�FY ۷�=q4S�F�{#��'F��Ʉ�iq�mC�(l�VN��XrfI[�{��oj��n?��Dnw��P���*��l��v:
=���/ڜ����^�<qk@~Ly��S���`���ݏ-��{�;`G�m&�<�p�=Kʸ&�������P7x�5QAWB��\�&�v>� ��	�縕�&v#ǋ��Am$|x�g��͐¬�
4��1�9�vFG�bm:�e[���>:�n��֪��OV�䋝�(Al���a7�d!"�:���c��I��y�'�3�R�*�o��6(�Э�-�<7l�6����L����dH���gQ@��� ��Uo�!�&���Q�)�7x���V!���)�qUP��6/��5˨��xA �#�y�K>��{�;Dҩ�M�l���y��B��x�E�-�g�C��I�+[b?Y���%,��:�C���i�A�UF���P�J�9����ڳ�?��{�u���a���
�,hbs�a3���.��!@�1����X����n�^U�u����mڃ-��R9xu�æ֧��(�:%<8���v�&���v��3��J��ҹ�YE�p��xG΃��}�q��s�Ns��G���'�@g�{Ԇ�夔$kY�u�EB�ƞ+S��Ih @����Б�h�~�%�*s�����e2Io��_���Q�z�����o�,4vB�!��"��rS�<�=����Q	�ho��婔�	�?�ĝ��S/���OI��x"͹��¹�ֱ�m��kG�M�	jP]݀� ���G���< '/Fm�����b�����ߌ�"bv	��C��iKNN5��9T�k��qg`Y�.�}���bM7S"I	�-f//;~�no�Ӷ���w?@[�V�!�3���W���q %�F���i��ш���ʾv�ś
e�X���l��,��7?Ig��lɶ�N�zob�o����}�U�n��XtY�Lg~�����\/^k�rf���@��v�#+�	2n���m�J��YNl�u��_"(�S�EB��`&mF�����e���x�K��t��&m�`@Z�r1�ڭ<.���,����7���/P��@K�C��՜�uE���9�.-�#���l��m��{�1���u�翤���7Z�r����
�^�ZC��� �)��P��v�*ߨ]yi�0> �wo6eOӅ�S*�v�Tj8���$���������mɢәw��zg�`&櫘Y.Q��x�v37̹�����\�({��$;vE@��	�Js!SS�?�{?�]��JߌH@7%����۹�bv�j1\�A(�/��q�!e[��hC��ׁ�?�F!Kx�lE %�u"�KȎ\���Y��-�����/j�D�I8������/Ѐ�V��`S_q��wg�)e?ј�L��oI�;_�M��t�;��a��!�T^_�A�y:��tQnS�Jx�@ 6U���UX��g��T%�X�Z���>>��qd����cu=s1ӎ�45�K��*�-+���}GQ��0�j��^{����=q:Q��FiE_��
����9-n�矤ͶV	����̔�@P ���\���]���
�$x��Eh�=���g?���+��d+:%�� /(e����q����9��.D0�+�vj=<�I�V����dSj�!�����nu�L�-�ZYp��<�-]y������Rٿ'��A!� 	rD�h9��mѪ�x��3�:j���.�J��Ӑ��ޭ�fu�~r��Y�-�'C1����!�_�i(&	f��t�i���:}moЮ�K�Pkx��LPNB��ts�gU�4$�SF00?����J��� �Ү��S���6$�R�+i���+�;��0�Ι�������f��fK ���phA���6�k��� ��#)K�a�B4/WjT�$���؍4��������s?Lm���$�^�H#/��E
;���J�ҽm�^�F����_Ү���5#H��
�$�l4Z7��8g�>�fVH#�bUb�ݴ�����r�]{r������le�P�tԔ8���V0����!]�g�N>(���$u�,�����i�
(��������%>@��j��B�:��S�"��oc�U�������8?��m@�C3����N"������u�4()��Ȏ����'�
������O�%����R�g�A���?7$���F������뎖pk�떅z�>�����_����B�Tu�f�*R�n#;��H������ݾ��Mb��5�\N,Ӭ�o��z v�ߏ�������h�e\�הL��<{�}���Z�sP��(%����~p���D.�G���Ki'�J����]l2+P�]Zx��z_T+�ӹ���]=���:��sW��1W=��R�O����\@V;M�[A��)�g1�=EA=|�:>����p|�m�#o�}L-�[F/��G��}��`�Db�/�J��I[�Hc���ǽ��{�/F��� ��~��u�͵~gj�b#�d�#����Qm�`�A�$!K�S)�r
���h�m��m�)�<�	ʸ�).�ݓE�W׉օ���^	�yy��lgsw��XH��|��vv"E���P��,p�=�T����(TTI#|z_�(LP��"�H�wWd�[3ak�cs�0�N����� =R��}�aA�rUNR��~ݰ\YJ�@�qB�Mg�MW?��+g?���9¢�m�TF�5�&(6�*_V�%�p��r�p�q��=�q��lNg�r��b��1�?*�N��r��Z@jUZ�5؋n���J�����%�m�P��ձr![!����@#���<Ӭ�hE�D��x
��g����P�pkr������<RMf^������o��ۑ�7��¦��dhf����Ȋۿ�V]b��Q����}�q?��.l��>�}2Nf��E�IT�\f�T��l��O�>��U�^�U�9�m?O#�Џ�7�Kl�78���V����2��0|H�6:�pk�Kj��Wr�w	�D2�~�)r�g�S��L�L�4�:>g��?�|2��yF�r��=�RW��?y�J��Uk,�O�����2�2b5QF�Dѐ���q�Ft�ֱ�+�=tъtbO��}�qÚ�~y��!��u�C hH�lcD�8i�(��$��K��I�t)��US�LN�K��SB4AÏ�u�ؒ��_��?_������eP3}���;�"��}��ݽ~:@���ĘOφ�g��=�N�tH+�E�R N����4� ��
P�L�ڰ5��(M��u.�r�gh��
��6Άeg�<}��G�d��	-�+�(�H�"�L+	���-���;�xO�$�y@�#�
���O=ś�ήn�P+S<Q�
-e��5d8羵V�?}�E��o�=�\�<R+��ٯ�(a�/�Fd�WŪlP>-f�G�p��v�'�\N��fΔ��z��1��,����ABc�+��v�	"�YU5.f�	�t�DB�����Ȱ�\�Zڬ�ɼ�)���
����#��-��(�S^;[?u�\>�^5)c<ǲ���rV�+�y��,W:�Λ9����Bm5�8�d0!b��p4}�<�J�hw?�yዺd^�H����s���_*xx����:�B��k���������{]�����K��e�z��k<e���`���l����9'�J��$�낀�)�<��넼Z��x,hdDs��;������#;�E:!�����hO�7�ȥ�/�c$�Z�ř:��)/�KV�i�U�O��*'�d�D���c[��̽왪�Vf�z:'6b���]Y*})-�O��(�耟c9��|+Sa�#j���B>
L�b���Jv/1x1�oqҐm��L�[T����[�67��WM�f��J�er@t\f�M>��C�H�590ٯNW*bM�h�V�����Ii:��Ծ���m"G��x�'���ݣJ1
eS����JU��8}{�%��4W��_���<m�.���+'��G�Y:J�!b�n���s0�d����߃m!ʺ�[�qf�L�Y�2i�6���_��5OH\�l6B��������V��KM1����|p{����t���
V�'(�P ��<��F����a���+��#*,+ ��Y��_Tp)9�xt�q�>n����4��ol����/L9O9��c�C�W�%#��M3o���dz%��E�:D�՛��m�T���#��K ��i�<�`�Nr[羔b��u^z���P�R�����vqc�݅�y�s�wr�Oź�����~mngD��|����fp0���|�+�\jAo�6n���U�ע4����Q5����(��+}n�%lϱ�6��g��F��/��nR��ʾ*��b��]�)��>��y�ύ���l�je�-#7I�ՠ(��t}�&���f��Cd�Sݧ�}ιq7��%�u�\��է��D[�����^�iʥ%��G|Q��;Q�r�tn7�E�5s������>��8��9�J����ǡ�%����`�i������!ח+pЦp�<K`�x�Da*Ti
����ba���(�J�~O�%�l`��v�\�%��pm8��%�p[
6�N��χ4F���p���C\堔񽻇��Ep	�Jɪ�f��-[f�|�AI�uOo�)=��0z@�p<�0=�_�nC�u�@l�a2q	YP�q�kP�s�����H�!�G��t�w�b��KB=��kC��N���z������ر
9Q�t���zr �h�p��ǌ}��.�v]����u+]u��]�B��ӗ���Գ�D�����Q�ϡ�!�>����7���'�h�;�ӻ��Fi��o~�"�N�	w7�C��[댔{�U��wӗK_D��G��rb�8Z_}8]�p��M�IPj~<��t�#���`byi���vQӟ4ėђ|d`m&���n���2vwCgO��v��������'���O���i�z"�f�p����&��U !}N�Ǵ���7-��9d:W��#�C��IXCkƿE���<��H(�>	���T
R<�?�T��ST̏���{EF�������o]�h��<M6.�r��R�p��@UP�4
��]��F�L���?���8�D�}�0�.PZ.q�������_#C��KP��8�6Q�G}��i6���Rm�,��gٮmN��'��ϲ�kK
>�k�u"M�w�+���<DM�����ձ��.,�*L�=K�b:�ߣ�Okp;S������_&�u!���P�fǂ2��-�!�6�"46Ryg�Ԇ ������h�^o� f≀v��=�KN�/4�~�`���!���1SK����b�G��wD�8�倯��|�����ѿ�NW��V�i�r��tlgf�ul�Pt���=8A�r���P�@�G�F>N���`�e�^��X��(��y3�y���PZ�����SF`�CB�+1O��*������T������a8,��~ح�e.5�O����)f�F'!�q:!S�j������C�h~G#kK���1MO����M���W���d�l��ţ#]vaA�I�'���b_e�`��F��u�$���ǜ%�����7�&�z@��E/���U�7>C�%g�?�L�"�O{4	Y�^`�ع���|��G>DMB���C?���8��w�<��<����_R��p��r����9���]�l�����4�'7A��s��Τ���(Z�zU�:�d�c��8��� ��G��)cV��>j���r(�U��hG��Mts;ܸ������dJN"�i�Zë:MH �=�kH2)tsl+��#��I��ݎ`��	�w.>���	���f�����FS}K�S7� $]��<�{�"�xa�̢���>�.����_�1ȣb�՚ȩ�H~hxa�$���]�h;�	�����A3����	�彏�[~�|�Je3���-*7��#�N��Yy�."�`���2�����5������A�]�B̘��*:r��w�Gf������*RY��D3 �I53e�0�|���q�Pe$�'|���<�tu@��h�BQYe��$�
�/!\�VI8������J��ض<���z��"�X�*�UD�NK��T��#��3�ޱ���,%�����B~S��(R�R2��n��R��8�Uc��iɲPe�[��!�7�j��	xQؙ;��~�n9F�߭DhX+*��L�O��%$I	���G9}���b3Ҧ@�W��j^,��%���%w��v��S!'/ �I�G��k��E�@��[7��a�ep����_Pb�"e:�b�v 9�a�F�(��u0R��[����z[($��5̂�u,�~�>yO�Jg֭yR�Gp��v#��Q�}%A"���R�pI%����~��k�j�X
��A�\q&��K�:6 |�<��; H���ݼ��������nva���~��m�/��l����\L+�7�� x�I���*�I��D�_��8fL�T��<}��X���Is�ꌊ
k*A��0�$w��_v;!c���Kf���V�rn� �son�f5�s�ͱ�J���4�V���?�QUJ/4��v';on��WȁX��	��x��P2�r8���z�����&.��ۄ�F�;�D�ш�}q�jꖟǏ�a=&�f�Yh�jl�K	�(�k��Rx�܁���v�T����ҎӚ��Z�'7���B���Pԃ�дc�� �f�Dе[DM���@��l>"��}��u?NP9a�{�3���7�����N��OU	�\[H�
�U2��%�g��z� ކgE��A.�V���d$�O�1�fq]<���)���(W��K'�5*oأE�*{��/>Q^w�n4��q��M;�"��Mw��@/��{�=9@24k����o��J�:��?����JT��6�8v*Bw���{��R���	 �}� ��0��=������;��M���7�0��N����mN��b���rЀ��p���٢�Ϗ�����ö��_=Ŧ�����!"SŎ �V"�AC�x 1���"b�;�\������vl���HD<�r}��ndܿ�~20'�i)N�v��棊JS����[���󒟿<��(Ё��k�	�jG�I�SU�|0Vni^��s ��d=Z�24�z{���$�X6(�j0A �l���[۲��JJɒ����_ը�֏3n��\�-ț2}QTuS���䀹J�3|���o
�Ic���t��F0���n֥����ɍ ���g�����r�:g'����%�H6�� �ĩ�]	���-[���q�z�IȾ����`��ީc}Y�8��\n��Ĳ/�"�v���'���LxYS�g�"����t5�@����z�,;8���a���U�`n����dO8j�ۘܰ��K���\��铸XP@(�?�,KPL��p��V���������!�cBr�@�,�7��;��Z�Ӻiۓ�S�s��c��.���N��;@��Q��T��� S�*碨���������W�!��=a{p��9ޛ�������f��M)Ԕ��.F��`�lvl�Ʈ�����'�}`�$�Ǫuim���o@��^	�/ݱ��z�"�i_IJ9\]D7�hי�d�#�͔z�n0��� {�� �b굲:�\�q���%M{x�2�z��#�c�>U͆�V�%l�+Pm�1�<�Aـ0L��޲���4�IRR'/@ò��,����*Zg�YI�o7K���C��X*���9�-�G%��ҙ�PC^a�q�=��Z�K�˷����	^1��}kB���c����B��[�w�Iv!2Ef{
��b=��p�����p%�Űa%�)/aI�R�k`��4=6&8r����e���n�����>Y!��n�y��nl���4��f�{Z܄�9#��T���*�P_Op�o���[�?�������+`x_^��c/�
��O�
�i�ݳw�%.��&�/�Rn�x!�0�0��L���D�BLϛ���}�8�g�0�P"O�Uo'Q��y�[Ơ�܄`w��"����T�|~��N��B}�A�y��	!:����?$�-:�X���?���Ϣ�"*�#T�����V�+����{��/@D=,pO���i͚|a�1we���Ag�-{$yN�
�:���2�9�͖��!�y�UG��u;B:�d!+��ڊ��m>�$�.b��S���9���E]�o}(�7V�/��iyb��򸰷��QMΪ!Ƈ��a�s�8�b�z�v�`��h5.}Gj2������LQ����"a��t^%��8v��!��
6xc�vΓ����v�AQ��,&*����J���	�6�u��1�v<�;/{��>�@H�ջ�2��ӑin1a�]QUd��mE{2�gs��{����\�[(�*�Lۤ��C��lt�<�9�ڳ��E,끞���En��0�W�+m�%��)����r�_wc���C�W�$�Z.񘃞He�v��Frq e�G�����S�%�_���OCZZ��6?�W=�9����֒��e�̋f�͌�� ��ś�/쯂+�^\	k��}Qe�����å����5��n��	%_ [#��נ�����E���e�6�Ipq��.���4�ĸ��6�j9����P�e��Fғ"3�!${��(B'�u��xA��ǥ�5Al��� �Ob*8f��&u�.b�U����/L��(�KB�zs������jm��Ҿ�o�'��H����ؤ�8W�,{�/��o1Ѭ7�������o�I����2N.��X��aX,|�m�4�0����qd^��76��Z߷���e����>�ξ�>�{S�~Uq�NH;@�<��9I�A��Q9��#g���p(3@<�1��:iB46�w7%�i]r���&NA��$3d���0A���0����#s��o�����1�ʩ#�d�Ğ(��A��A���>䌋i	>��|$�Q�ʶK�.�7b��	�y#g�����֧r �ԩ���Q��H��.N�]��O/xL����?�0v�l���!��]��7'��n���לݹu	��**P�=�8�&q��	P���Kփ9�?u^�C��'Ӧ�����*�5�����l7�ɕe�b� Ed�⓸(s��h��LH�2[�0��{��Η=,�tj�ӹ��
�m�Ԃ��I#��K�7[�{��(P��$�&<k��t�U�E$'�P�ۛ�$����/��J�ř�L���Hmү�2��2I���Æk�T�U��{���1��l��Xѻ}�����>!9��	3"�'�:������.�@���%�W^f1\n�$��`�������Z��z5�v��(�ѵ�D���OҖ�����z,�=���g)�C�R#���E�r`�{�rP3�*7�٤TcQ!͎�o��D%�m�<��2l��L�ز\��:GH��5z[!jL���0S�����l'����^�"J[+�~��[�߶l��67�������|I��w�a��׫$���/:P����,�Yȭ~/���k�����T-�~X-����s^T\���4�fGv!�	���M��=�1��y���$;�qi"��(J�yȵ������Jv������K~�MN#��F�w�u����PAj�
�%���d�3Q�ǫNFxb�;Knh�c>D�m�怘�����f�|׏ `�\�W�WT�ѩ%�,RB���(	Þ>�4�á3���"?��y�X��)G}�?.��#C���{��;����:5�b%�$Z9)�� :=b�v}�3n�y00Gx 繝p~ w��gK ���c-�A^D��<��&a�*^�܎�x$�����?�
*�����~vU�@be�U�����y���������%YS:��_�v�_�Om|Z 2��B;��yP�I����u��ϋ��P䰒s�"u�笩�_c
�,[R:��tz�)���8c �:	�b�lh@�]{�i���@
��9�8\잿}p�%�7�O��S��[�t����gZ8ف�A�4�-Mf�z%^W�����#:#Z���l�l��4o�o59HrW'[p4��.�$�5	�m��˹C
��6�c�aT�@�K��g���8nB�FO:Fo���)q�?L�,g����x�!��wL}L�^;�,�����<_���͏��#(=�=ᗚ��C����=��B&���y�[s�b��J��^���CF/8�S���kھ�s������L�C֬��]�$��!��%�86��y��z�R� ��1-��&lF�C�q1":X�Jt�&j7{?��M�|�*�?D\<�N�|ʛ[�� ��N��.W��LiC`��,.�A�}-X�����'ʞ���i��%:^ݘ
���W��M�[���	�$"�L��m�wϳ�f<(�
5ɋ��fi�{$|n:���݀��kd5PѠ|S�b&��M� ��� ��(��	]}wu +8�VQ�V�̆\B����Q�ϚZ�6*�l��`ۘ[fV,����_�W�%�w�/��|n�����)�2'�:"�"6�Kx�|:.Ey��N��c�qe���; 	-ƺ	�̵���á�d�x�8���I��9��2_���]��G' �>4��uJF�fy����F�D�p\�Vi+O�7=gz1�`���v�]�zr#�������ۡ����w9��9����N�����_�37��צ�y��
f��=h�&M�}���'���(��xp���� cO�Z5K�#�����*NA1_~�B��I_��V5�Y�(�et緾6ܻh�i�{%�KK����]N�7ݵ�M�Mܸ��MV����,s8�q�P&���p���NG�P�vV����7���>����&�!$6"��QkN��̉}�x>����1wHJ$����T+�1��|60�9e�8��,��vx)kZa��Zc��� j��Y��ϟ��Z���߲v�'�*9���3�t�8�:� ��5���VM��?�U>Z����!ċ -����'���� uw^��#G�R�d�4�a ��͹\���Q/!�a�}ֶ�e������E\�������%�2}�Z�v�t��������6�V�Bxsܿ��P��	x�Z����;���K�]_�|�����#�7BX������ce\�e�����m��̢�O��K�[6ogL���c��p���byȽ�C�)���R����9��"��[�p�I��j	���t1�LZ����.��u�_����-b.�Y�xP���+Dn^���X�B�q+m�G�$�^س4���]��HJ����,o:�Rۤ�.�cJByv��0o�r��� �uyj���-��Թ��|'b��@*E]iDp'bd��x�0�زq�{ǹ2�7�m��PO�7��lD��"��؟���;\E>	����.�D�ZFy�$��U����η��g!Nŷ}.ܒ-H_��R�!�7�׵M=K�`��9�3�Z]JI]�bi|�p�4�k��2��J~r:H|���n^<ڌӅ�PN�������o����?�� ���)O�yi�N�{��Zk���#,���c��>�1Xu�)z-Rݎ=|��EN�#2�-��J�sF�6� �����6��~q!"&(���e[�H·�Y`��N�]	<Fh-�a��r:�ʤK����hʬ[�x��]0sS��fA� �cD�VͲ��s���:�����Iq�i��v�'u`��SAS�ooŐ~w
p��p#v��8�#�(��Y�Ч�9���X���Z�� �N?D�U���*����F?���:�;�H��c�3,��/�pǟ�*1�$�xD-M�7�ǲ@��A�����ʨ�)r��� �T[���0ܭ5mj�i�@z�K���D��g��P߉E;�&e~��0-}Nh3�p���/�v
/މ�Hi">3��������VQ�-�SM�[}u*��Cb�yC�r��	IӨ�|�5J)
n?6�����~���@w��'mfsi���C��3�	����A8#�ز7�P�ɥ7���j��^���:�0�� �6Zf�K��5S�܅�:�������$�UG�1�09�թ�C�o�V���Y�-��99-Ƶ��6�T�.I<4Q�&�+��\�ea�o�#�-DD-s�LZ��@�:���Kk�-
�3�!�����Wa�ǯ��/�FNz��S�}���J�6�[Ú�e�eE�1��M"d�Ko���9Yn���&R�ڭa>d��w��D�u�Z=C�`|7�2T;�8��ܳ/�3Z��
-cto���Gǉ��-gĩ%fE���h-	\�#	[�R4�|����'��u3�Z�c�i{3P\G��8���n�谕�P����A�N�e)&9�֟���筕cO6���g����.������Dh��:`ysљ�a��x��PL����b����c�3�^!`[��8��VyPW�>g����'����3���~� 8�F$�;�G\{AY�x�������~�����1kB.{�њMX6C/7H�H|~�)Fp\�b��9�J�f�pa�	�߆sP�Tq�9��Z��ptť���'��O����]�s�� �An�޺�c�7"A%)M#��˽^b��h����:��"�65aK4xָ�k ��La�r�
�|�{��P��q�x���6D�������7\�U������r8�_B�m`�g��G�3�|�@&�D
�N%>O�Qp[kQ:��\�bFi,�Ⱦ�o��6P^(b>�#�ka�T����L��8*��F��Q�+
a7i�s4Qu���$4�ڠi�Ry�g� �13�L�i�Kn��V#���|f�|��D�4�R����*T��T��\��Y��&w��$�XZ�eb�C�+�qv+ݘ!�D8�����C-hic<��P�kSؤ9����V��ƃ��&}��IWTml��/	��5�S 1���X��-�4�6�~�]qB����/2A@E~��ks#��wY��;�@�H1:^/^��5Th�n�KDm.��������/9+م=
�"5�&𥤀���uI;s(��1����ޠ�"!�"�ꮀ�2I`�`ye��1�K��seY�Y�!؁"Z!�ʜQ�Q0����N'�o���7���洴�g�*|MwO�Hc~b�au�L��3�m;�3:	��v�2q]n���FN��f?�fn�B' {�����"A(����]o^��P��P4�g����I��WN�E�;�m u���]Tjbq���Z��\�1�.P$w��F,+=��ӹIq5��_�������(V4���;\y�u��.#�q*�X�4#�CgJ�7�9؝	s��[�=�B�����6�h��u��sw"Q����H���I
�k#��m�_|N�
����"�#c&�|�,r2a�N�����ȴ�(���>ۜfgbJo����3�9Q��Hl�V$Mj �k���e����\0�So�GC��)��{FX�X����IdW���"ȑ�V{�+/uqJJ��iD���t�n�!�(�������X������c9c�	Wo˲2�_4B?)[(�,1�a_��7#R4}��vHE�g�Vyma��e�h$� 
Ϡ3�8����"�@*�2����Tx)"��@Y��m%���.�<�{�mҊE�U(pP��y��G6��,xji6�%�:�ޞ��-�/Zݝ�u��]�^]�����b�� ��&K D��2eٍ�`�S���	��|�ઓ��#&`	����@9�_B�ɤ`�O�Ok������,�?u�X��6��UK�=�b&�L���˗�p��gCr�N���c�S�����G�}�>�\�z��5K�%�Dc�q��M$�w9��Vb�WKD|��������X���j��U����8�x~8;��֌p��\WY�>�I�A���В�3�t�B��X>e���"�c�S,���	˂���u�kh�a3cI��e�Rt�n�y��9�"6��I��4{�����-�H!��Z��O��~g��\�fw7E�EV�?,�(���=�-���ɺ��჻yI��l�rql>�'#�����s�,zh��|��lV���J���b{��	+��#��3P%SOX�;Bh��2?����[���8/���Rn�a;~����7F�79�B7\�^_�A�gF8�Ԝ'�W�\��C�26%m����z��U�z.t1��rd���K>�	����QV�9:C[E)\XJ��%G������ �n��r�+zu�ւ-uH����	�K���N�q�8�h ��i�ۚ���$+����z��$o�o�����	�Z�Ǒ�>1�wFz�2$�#�-��b��Y�(1�&�cE�مk�ު-��F�Zm3ܮI�n�ƫ�րg�;�˩��m^����W����7l��y���TA׽��"O��~�`�5 K�{̕�%��K�2E���w��'+K�S�Kg�%p�P/����D^jH\6�kl��銭�|w[P@��;0�����r�;���툿��	�����{��.IuT���RQBV�.��2u�΢/I��Q�����eE{���2A������
UPde�'#W�;
N<X�/��0BY
Ou_�W��[E6�J���x����8����I.�P�ߛ7S�/�=�4�l�������������I�Qh
���KҵT��ՒІ��X�����x�ѹ�$�"���{m��[��/�VUjĀ6��>��Gi�46P�2���7�ʘ����+#1����ƺ�$!��Jҥt�Hz<sA)���eK��{�^������[��
�<�S�?v�J�n���^s�����U��V3@��Ҕ�ɽr���̏Ɉ�hka�w�B3m���<�ƺY�xϡR+wa��	���lؐF�EI�3�^�xs�g��R�x��~}�h|l�pt(�-p��cc����g�P�����yT�"b��O!?L�6���B�O�,��rͱ�])*�	��0��� w�L����b ��c ' �iu{�K�7!��L��aʎl�4s�8�$�t�$^+��Y0�6�&_�Nw�%��צ�i�������[��.�,�����&3S�6�.����暣Ű���v��jJ�	������׬Q��
��{����3Z�E/��݌./������E��j�
���hk�'>�a��|�y�����V}<��D����͝񈙎�=S1�Z��4�\��좲�����ܙU":��@����>�6�}�\G�]���-�RӀD�]n�ؙE�ܳ̕vB"�l�QŬ��2H���>�r.0mI�W����q_��@v�z��\���fDv�O�OZ�tT��������^���vs;�,�pz�?�$kX�����MÐ�����fy���l]7�|E�vy��2����p��=W�2�䭄Ҁ0E��/x>Kڣ�sQEú�����>^kr���=��[B+;�����C}@8����N��|���\��a��{�q$*���a$�>��&�2˸!�%�W�R�V���P�""[Jy�sFI
5E��aߺw�D!E�7H٠����#4W�o�+}��-��$�=���?2P����m��07�/@3��!�!(,m���L� ������tp���m���m!�_	�3�pODyƚ]d]tK�����C``]�3�3oq�\�㠡��1��tH鲳Q�p#&��� ��˔�E)�܊��п�1�) ��4���c��I��J�������Q��o���S�!�t�ȸ]���ųS����ʥc�������кń���9�F�t�^&zş��+# xa�o�8�ڬ��Lg3[A�4"�l��n��������!�!ޥFH��A�xǇ6~I���<�7lJ���Z�M1�en>�I�����k�Ǫ��z�o���U<�^��f�s����9YY�v6F�o�s���7��C	��jL�G�Mi���5?����`�$u���r<h>�����_�m��9?�b�H�~T�H�l|�X弧j�� �J�>�7�
(sI��-\�zM��6�ض����Cd�g�oBw1B{-�[�hw�}���I�w^2��r
%��\�;V֏+�* =j�ש�w�*��`��}����L���dh��.Zj�;��FH�QJ$��D��݅APj�WW`%�:VsA;3}{�Z�q�u2 +N`�t8��u���=�q�)Ⱥ���U�Ċ��ԌWr��q����W:ϛ]�v?]���S�2av4S�n��|���bxT}R//�����S,��(\��TJ=+�K�W��tbЈ������Aگv�W�#^H�% �ϱ̒x�Pj]-�e����\n����{JR]з�@E!�s,�9���M}���̂��'�~?�:J9/�/D��8�����^[���~�٤a�����cU��?����
�#��۸@�׽O`�C�eЈ=AH4&�o � �Q������e�׬�Ҏ�]��;µ)e9#|{�*oX���c�O�U�b�ј5֧���&#�Os�b̰7��aV���
�N�q������0W:�qӾ�l���a�"�|`�c�T���"׵�U�6�GG/��E��Ahx��Q$���_�ֹa�	���0a��x$�ehR<������,�Ӽ4����v�PWgS�եU5�C����5�- �(!Ib1��2���E;o`��=��1m��� �[%��O)�H�X04��GA[�E�9K�=0�5����������eg��O�hC��� Ї��{������$Qm�2�����,�s6:���G=��$�[2� F ��S�c�Ե�ߋHM�b'�УX/� ��x:�T~�O~u3b�IC,G%s+MT�HR#<��FY��L�[ ��1���J�]N�Ѻnd#��!5��φ�I���&0ڲ�`�����`d��?AS,	NR����H��`�mah��Խ�4����Y�%c�Z,{H����>w��YT��"��'l���|+�Z�X��n�j�_��h�K7Z$�rK+c~ͤ1��gybU/�w\�ǯ��[aV�A^+������~�И.iMm�ȧ�H��л��b�M���-#`7U��iТ�+��O��/�I�C?D�ƀ���<��l_� �Ά������ו1��Lm��m��}�Z����j��l�/�D�*��[c��հL'S3\F59�m�򀆆��@��f����d��+�Rt�0�r�E�.:�/@�Q������c�A�K�6x�?�˘�)�	���}M�F�o��Zt��Ţ�-�}�(�<2��}'G��ȫ�BJ����o;{q���wRH��]B���?���at���DA® O�ā�������)�U%���Jr�U;�ٮ���W��R����7$��fie���̚6j���E(�9P�,���'��%��`㭖	��zH��w��4�Խ*�����y�u��V
O}����>��-lԆ�/�ES쳂�l��8� �ߨ^����@�77�*�n@v�\��H� Ռ�\��M�%��S�Sg|�������A�pd��S�7�-Y#lc�5o����p%��f�i�h,Y��QꮗF�'��B�%�:i5қ
Őj��{ZH]��Q����i�$P�t�������?�õ2fs��ZR�m�@>�v��ߊS���'�@i$D��٢�W�'�b��U�{l��T�I4���Bs����O�E���4B���c��/��KN'��)��k0�2��k���Q۬:�1��݇Q��E��q�@�{���~��3�����z�A�����-c8#�փhD�|uR��=7K�U�.il� ϯƜݧ[3���6�����x�ʯ�V���gSB��&�VD�4�i�;�,*rת#��-U����Om�םc9�t�����������S~�R�H5j!��Z��������4�-:p��BdF�� s��f�,U�̨f0y�/.�yk�b�|8�/ ى\.����"!�>%���M=�"h���R�� W�Q�+�84w�ɉUU��@�'���肱��Ù��3-�� �β�$��lN7%����Q����V��uy�'�	����~�S�[<Й�w�3��� 41k�=jv�rLV��|�V<��x^���: �ir�+�&�$�����̒���5+�w;m�W�z�uMz.����@���<,�{_ͥ=OAԻ��$���B�ǣ��jz�=e؟�-s&w۱�o��D���]��V��s�S_P��lg��N"j[�@:����_L`}�/��'�U��E��c�a�������o��rA�H�ٝa�����O2x=��0��i}����p�.V�_j�6l�k4��Y��R��N%��3%�y�[��Um�A�4�E�`�������]�<�_���!�C���͇��W�<9c�+T�y���4�\`���X���H2�\t�fo_1w~�O����� �0�	;���$��s�6��	k��X��<U�]t*����۳�1 �wD���sm�cia��ie!ҍ���R(�GF;�0j�!�L�C/���>X��&J�Ŏ盜�z��؜��ٻ3֢I�[(޽����Iex�dk0#��a;�9��m�)�����#;�sIΎ,!�"�I��E���9_�׎�#�~-�,|�&'ڐ~����B%���9+�.����e�ٮϬcw�	����gV�c��N���V0����l8�LqZ����)?f����+�%��^��P~	@G���%��&����h���,���?��c����	̂�S/���/�'=7<q�k�K����A��H���y�( "E5���ڻ|��w6u��oX�e�N斀�M���x4`3c����TMq9bߪ�!���u���uq������&��qd���m��<�4�q���6�;5���	�R�A���6$?��4���U���"�}K�X�G#�,�|c�>�Dg�^�S;�4��H14q�)��E+���/'��}��vA�|�	�FZ"8����6��C�:�g V����w���C5x,:�4<B��3.�''�df2`�˸�Z��lm������.#V�vd?�� 9���p_��	k-oz���-`:
�|q�
T���ʸvQ�����.�}�Qx�6ŗol��F���h�?
��#-%�/E!���Pw`~���W0g�#�f�'G��:H����C� XZ:x�+�z��-H��øl�R�.<��1֟8	��]Q��IO𾹥��n���+�����X�*�ٰn[ׄ]1����Yɠ ��CXJ
�i��#�zi			|V�g���m��Ɠ4V�"B��+�ei��Yd,*��8<l���կ����D��ݯ�}�z�u���Z��Cepr;�2^l�y5?WyWk���<Y��iS�GKO�1�Hfa�y.����Q�X�2X�� R�e
�h���׳�J*X%q"J�D����t�*Ҡ��i��"+��c�v�GD��!�I���%���Z�5Ѓ�Z��?/'|�����H�r� "����Af��$�-�A��g�-*wA�n����ot��0YpU%���"a%ʧ̚�q&�h��E�V|]\-�ykC"T�ȅܱz{.����WC;�����x��C4����`�;�)�Y��6�߀{��$�	a�x{�'�W7W�������Iċ�ms�[^0��r�r{d)}m`��R^E;��8-QN�g��z���s#n'�<d�,F5��������iz,����z�[a�{�F�w!Zs�a�Hd=צ���[y��%m�����Lʌf��]XWv���t{����w�?&98)Y�K-�X��D�v�� �f'py�(��*�AHM����q�Q��"���>ڳk�|�����\���m.�H
v&�z�0�J�&��_�O
1�����f8њ���O�<@��(�L��m3�ڢb�	9�.��mҥ�Ey���2*U�q�B��-Ԃ&u�S�ߩ�1�r����{Q���NL�V�jCVô�_�1M_���p|��e)����k�^�n[6���]1�,M�X��e/q�'P�:�a[q�H����8K���d̛D�-ALm�<�����R�q
n���t�\�]�a��T�|�u��Z�M{�T"T�V͛s�r�)�	v�WZ0������I.��Zv9��;�ٰ�q�Ն@�O;}7�;�w�Ɖ�
�F�W��7�n���5b�Haj�����T�Cl�nBs�2{�� �H7b�x�7QRҽ|S?�<{
�f��&%7��tu��Q��U2��Q�Z�?�y�5����Y��ױ�7P��V���%��f3��bvu�.��Y\JZJ��@�N�xe����QZ0�jR2�����^z9WA���3>���q��O�}�>�$�@˄;����y���&��E�(�������ʮ	�G.%X�z�����!'����ʍ����5��lR+S�:W��������(�V��A%M���>���1��>!. (��H]3����3��*�Y[�V �0�3Lm���>���*tt�~u���c�]����u�µ(�-F�)��!\��9�)��X� ��D���9�XZ������b�A.�uK��+Zժ���������(q�ߓ�}���@'�?	S��x.0"��xڒx�I�7��Y3h�K�']��)� ��J=[�[W��j��] �!Q�e�@� �Y�m�V�a+�O��~O8���O�]�j��8̈́Jy�S���.����?	�����x��O�">����v��|����?f'��5Z���F�d���bbn���l��|9C��2�u�8=�/��#���-m�tbr>��kxmDv�����tR-5]@����"a�]&�4�sGh��GΞ��:���ܿ����r���Ɓ���˜����rj�Z묉�ro�@`С$��L�~����	��nx�^���털N���.���L�R��)e
��B�Z���ł�(��j��,z�����4*c�K�o%�4;No}��:ܱ�C��}]P�Zx$
�
����b�;J[�Sต�5ڳδ��4�zgۯr���(i}em��96y���֠S�_Θ<ا��D�m!�f��j�{�N3��A�v{��9�������0b��H����v�$G�H"��r<'�7�)�x<�mA:�C���{�������5�@i���n���k�n���%/�I>���U?�3�v��	�@]4pW���ke�H� !4a	�(����f~�!��g�a����=�!2�^����j;ֱ�sy��n81A�B�3\V3�W<����3��r+�#)M���k�[�;ϹZ�]�DV���L�8��9�-�fg3�^�l��K����ѝ�ɗ�P��! ����eٞ�ﲿ�q-�)�I����x�E/�؋��H� ���Gl�	��z����x���n2�h�VI6.��zbF�����q\8t�T��> q/���&ڇ=��= m�Q)��/���x����?�1R�٫Ǝ{� �I���*����7#ښ�bC��G���ȿY��o�(:����u[����a��z����Q		�
��݉q��ϔ�&�?5k�} ��]Fk&� t�b*k揧��ܰ�ďr�G�˽�vܰ���aH�ኞ��yy���6�<�uB���}�~U}C�LM(c	��,}���N
H���Lk�\��I;��/�i�<b��Sn��i뿦-���֫���4�����p�5ӹq����®��������͡�/��G*g�L@d��ꖣa��Y��T�!�B�{d�zU�z�j�C���b���Q��o=x�j���4�_��12�YJ���:��M�F9��=v��$4����v� �y�yc���[��@�����J�Xjv��r�4��/ezg"h��*��q.?�{�� `+���e�5��l�׏�N�ʴs8���sR>���Ji;�x� � ��cr�����ֶ��/�>I[V8L���"�l���j>�/�����[ՏOT��;Oj��h�~���y�[K�J=��7���x���8:Є��Ш���}����Itw�h�8����â� O<d��cV�;�b� �
n�sn[G�?V�CF�,��C.J�-��o��9.�����x��Z1��TE��	LJ<P�wb�n���ǈ�]W�y &�þƚ\sL��hi<N�Hp��m�^��M��T�Μ���U��z��.O\ݡ5�|V�@4���Me�w#%r�(�+ �#��>ᇔ�v�x�L�
{1sиQ�;8�y�X}_�OY�2
*�I���/%I¢*��$,%��=`x��/^EoB��2 ��dt3���G� �l��x	C�R�|��"M�]L|[5�������	��E�
u�$ș٨���~��_���gD��{��iw/�'��M/��E�V'e#�P�}��گP�����Ѱ.� ��8z|��j�zp��UnZ�����O�4���E���Z4kS�BC�T��O��0�t{�8'����w�s�����a耭��IO$`�t׾,8�^���~լ��k/��zc���~�|�	*�(���\��H�dd����#�Cw�B�{�_����G��q��K�xrz�L��(MYl�Sd%��g��sr��p��2E�yDV���/xq<QШ�=�N�ܾ��"�aP��:���7H#4KyuS�t�G$a�O$�|Z�s��g��;4#�8a�l��Q�3:A�[#��*��i��f�J~c�3ae�lB��i@Y�c�>�8��X�Y�Z����X�=C:(;p���)� �����q��nگ�W���Xt�g޺�C9�e�pe1��|!���b���=kuI�C�Y��s���Қz>��c}#�\�����̆��.��y��*S�燨��٧|��q�D�˞�=Tm���}.�z�#M��|t��`P��f�fO���P�`|��+c���%��p�w�5Y2i�v
�u��w\TS��oo��o����m�{Я̒9�(�7������M���ΠQ�¨D�(a�p�i�A��7�ODMg���~���u�"nQpt"�u/X����e�Y���8[\�e﷎����&�<k���2�Y�G����w.��yF��g#�< ']���y�H����y�u�Nhߣc��}����"�`�ʃ)&�C`!A�K�Q����BS�3�NE��T�,�b5��Q�"��QiS�b��;lτ	+���f���ԣ�/`7´��ߊ���BP����
՞�;|v�!D�Y�� -.:0",g�P���|�C��t�ъb�k3�}?��a��D�FRB�4XL+��t}�Y��v�� ���.!�Y`��(�牬�݁]h~��{:���
C$&�we��#�?Cl��$9~����hJl�x�yBB��9�$���IB�0��,���ް$4�<I
~����Q��mT��۵*Ix�)n��EIz�)~�ӽ��"��%�M��n�M�=kΨ��mYM��u��,���a��<@%o��yOMd_v�� \u �;�3I�Mj4��c:�5�k�F�c>���
#V��� nE�@c�I%��]�7��fcO��CF����)�~c�\s�f6�:���-�CN��� �֩t>
-�8����^vq���%U���H��Kr���K�],^��$G�����@�j��E�`�.h�6�O�
�q�v���H��0��vW��X�QFP�@����/�>Oh,��e{b���3���&m��Ŋ��J�S�o�	`6���m�ڹ��0��cc���2Q���ֺ�i+b�񔒨�`�GX[vO�(���#�&�2�-���q5���B��-`���;0�vr�:Z��JO��qh����O�B
H��5k��h$���lW��$��"���:����U�%`3�m�.$�5���Ff���6k+�L�V5,�o� 7�X��5�it<a�{���Y�Pa��l[�4�[����F��h� )�GSWi���,A��!���ྌ�[�Go�t�1�>Y��N_@0`���`��m�q�xcF`����l���SI��I����-[l�Fo����&?�Sѹ�WMeƩ��.<�6�+t뒊� K�QGT�`'p���A�&>]:!��#��wK|o�|*�ҙ�0�k���I�_\p؈���W=r���e��m�B�%����'�h��LZ�O�Eil��[<����*����Ll� �蘡4ż`����~�>��~����;F���B����3[ҾZx����|kX�B���ϋ0�E�	�v����ߣ:��`����,�'ޥ��;L���`ī8��˽�3��k����Q�e����tѻ��+�]��(�����`�p+ޥ<`Whp�"+Y��4 � �ʩ O�8�>���Z0+���q&��)�j3W�ȡ��+o�z�d��|���i��;3�����Gu�~F3�)��`���$�E� �R��}-�GB"��JJC�������ޗ4l=���������zX��ڬ@"���.�u9n}q	�u��
��Y]�#1�S�H��X��^޿�}꤮\F�?����: