��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_}���l�'���(p��9��^P�ᰤ�P����LkSU������6��R�"��»0T��#���o�����ܝ���`̓���b�f�^�s��ٙ�Kq��K�=5��O6�ٽ��j��t��Z�ܾy��e���o&�3�{��P��dDm���ѭ���t�tĵ���X��>�����/� >:;��$��.Pe�{��7�2��ך�NG�օbżs�s<�8k��]n�P̐�ؓ�uO���<-ԧ�WC�
'?��a��^d�T��}�>��	��Ί���v��l���J�������o\d,�yb���N��O]&Sӂ���|ߞ;��7 +ǾA�'�.8�Wjx��F��
�|�	?%�趾/b��ט���p��q��t��6��B��˭M�z68$)��C�nf^(��TR>0
tC��8�D<���a<X7^�%#���I%/��f�����졽��P@��d [�d��<P���4۩M���~I*2�U�u{ �1@�T)��80|P��:�����b��'�)���d�opj]�Vo��=Vh����K�I�[b)�z�񺞞�JWᜁXh�n��%��G�D�'��=�@~i(��@8��Z�Qİ��kl�:d���"&k����dٍjD�³�*�o�I^:�X��Cq[%X�u{�C���~�©R&��M��]!(~<�AO/߰�0fkj��=~$�ll��
6�<��U�a)c��P��/��!��y�u���h��zSە������� }�3*U�{��V�쟳W�(NW蘁��n��&<,��L}%�$@0���i�
;����Z$&E��T�xq2�A�0���z��h/��8gD1	k�/6��?R�3e&�������(�� xD��z���o��U��KL���{�6V5�S�ec(*%���N������Ԍ؝] @�M[�W����[�)*��lq����ʧw��$���o'�<CN���(#��#)Q�'B6qy��� �`�lQ����U��e����Ex'�����_��6�;<� �xњ�g�g�%!�ӝ��+�>���z.)����t
�������g��2��0�Z����Iz�g�-IsY)`J�tZ���g�P��&����S )�~^���*�ur>Y���|���@�o��>z-�Ϊ���+C��O�voH�n�6��ѕ��{�[U�*���+��P�mq/TID�$��3��}S8w��Ɍ$�_$*�ƕ���p���m�1{�,� (�[�*�[a����o���}�������*GdP�OF�g���vKHL0�9�F2�e�
��>���Y�q��ѫE��~��Uz��B)2.�UJp���7W�2����y����a�L��d�cO�Ζ"�\a4��[��GWi�x7H$��xq��E�I�;�y�+��k'�2o�xOtC��ۃ,�$-��%e"w0E�lZ��i6?S+��l�/cl��I~G�^� U�~�,X"��qeÏ������Gg���z�HV�P�VgͅA��Ţ"x���m+��� ���.����L�����a3��}h�A��⎙���Dΐ���e�݃�pF�.�u��i�!����g�6����2�P|TP͓#�S�N�t�9M�*��k1�;�ѹ!쀲�P"O����B��zG�h�<��FV�x�<#��������> ��z;|ų�d�P��� ��W�vs8���75���c��g.`��?VI��'ͤ�X�ckôP'|�|�2e���_�u"�𮝦�&=�~H}�}kiSl�uW\��Úd�N��Xa"(�W+C��C%~T��j��<[���ѝނ���
��to��$�����K�<������0��QP�nܖ�+�=ܦ�
[i����+S��t���N<Q���
ߒ�	N6��u���m�V��5�-aCpy�	��~�l�{f����Rl��ٖ\�$"r���ǒ>[2�U�5>4�����_���ӋW1������}��P����<B=�w8�" �,ac�3����(�%w�$�t��W-�@���be�By&|����ةX[ak:<a�RH%��Uf*I_Nt,q=���F�°�*~�7S�r�_.�J���5U(~,�S�
a0U�&wܖn$�'��^5�r~�`L��.� ,��R�=��˙a�]�ؑ^�T�-�홱 �oƌ$�|�w�2�L�+�7��R�UD�;�%����A<5#��Ui%�NN�(�~Ⱦ�@*�q��SSN��ҋ�H���|~W�E�����G�@+�,��$S\,�M6
��6�(!�Y���a����;:����J�����s��k�Xwm�|��'���G������*�c'���� �P������Ǻ�4���I���吓����ϓ�U�ݮ5�ع��6��4���e}˗��!�V�G�d2�r�k�mA��f0������^J�$�0W���V/�߬;������.SzA����\<��\���E}Ce��T���[w��^0V����8_uۊ>�f���+�뒼����)"$��֤�K.S/ǎ�����+�0��BcXjm���z~�l��v����\�Ur��$h�	� K"0��?$�c,��܃�e���Q6��!���������SD���Y���*L�,�NaK��L\haYUO�n��3X�� �>g���@2�{��p�Gn��PBkZER�T�}�5�J;��S�7v�?Y��ե~��v����YWQ��w|���*�#�N~"1����5P��oVTglCaU�ޯ]�^i�h�g��22��$�O��ˢ�� �
z��
���R������ÖnO?�
c�%��M���PْV˸��y����В�#g��S�#�7�#
��4M�{�*��\_DA�t��m�K�f�U'Cl.��p��Lhq�a��1ӘҚo*2��a�}�؋T�Q��{����Ky�+ �+��N�/�ǜ�D�N㩈��y�ˢ˷����������cX�EY�U[T_��9�,pWU��%�e$6��c2��W�[-�=zB>r/�X��·8˩��84�mS���^��p%����`衆o�pn�����u�u�y�����O���"��z�}bJN;m�ױN�5T�{k�ٜ|��I��>�/X���ȐE[���֪��˅q��a�t�vX�zx{,��V	Yh0��ֲ�R�]�珨�r�]a�U�_�Q��Gz0,�7�N8iE�S~�4�>�e�i�x�B��(���<�f�p�5&�I���?Me��G�G��� 3&,`Մ���
GQy�U�(֒� �����T��?OziX��6�3{5E�"���åTdj}-��=�gap;G�caA���e-����>���=8��?�B&B����n&��7B��U�9����O���@�˛��$/=_r �0��6 b ��5�!4.Hm<ÿ
�r���w�5Fn7=���p��(��3$�K��P��- �jJ_F3�Up�V�-o��r�8�����H��k�����*�)f�Yx����-m)�`�[��gy/4�j��bXS�:$<�?�Y!��M�F_;��{@$O���P����~�T6 D�Z>"���E�$�c��|=��%��5X��Dz�$e)��_��'��	/�����oKZ��a-,w��� �[�*�/1}�~�/LԾ�f1����T������+w��)��tS��<��������Y�8O�	��;��fMeO�MF�R�����th���~W�C�|'�)87as^A��uR��%2$Zy��7-W�ND�ciq���J.��*[�)be�U �f�\���O}��@��JI���ا��h�
2$K�m:�-Qբ�G'�E�#�K�EyH�:�a+�I�Y�E;�Yf]�j�7�0 ������S"Ө��`�/���m>��ۭq�*2��'F�SD	��mM��?7����A�(g8�?|�?G2�o&�8�Mq�4�������wg���9�ί�� �F#�O�'x�XMD}�C0nQr?�4���ç�H�$�h"��ܮT��Ț�k� �C,J����<6\*���6��9�W1b'7����2�Vo��	�t���B�1� TY�*d� �C�׫F�Ov���2n^5uS��n�	k�t�YhN�UP7f��az�j�v�k�c0"�ӚS1�;8�w��-���R|Uw���C��i��V�T��V}.���EtdL&��W���Z�Nh4�W`2��Ϲ=j�)� d���p��>Y���� 艨�Ht~�/E� �97����G����#��h�`��*5b�q$�X.4�ƨ3�g|Q�@�6�SV��3H` >�r�y�:cM��pW�s���%x��և���� ����!wD���4/T�9�ro`�QqQZ%A�rd&��l�~���rk����S|�Q$�)lAs`Q����N�k��c$�[j���G�1�8&A��x��o�~Pf X�