��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_A?N��Y�jo���e�YI��#~B�t��@E����2u�@��G^��8�=�Q�Ps�t�N����ꈱX^�1��Fȑt��X���ސ�t\J���6����9*���$�L[P��#L�pfR������N�Gm�IGlr�FUx��盆(0�ܥ�!٨Im]�>��r�J������<{��	,�Y x{��a���T���9P7	����p��(p>��7YN����aD��Z�<�ѭu�W�B#�X�fn�ٿ��f����x�ڦ9B��B߳&B�24��f�����˹'qF�R��nE'��r=	���Tf0��6,p���g&O>Z���^y0�S.��RF����v�����CG<����G}J����y�'b���Q�;�K����ɘ>��سP�̫�Tہ����`J�� ]u�"��Mҧ��Mx�(�Hw�g��qV��8E!/=Н�-�9�E"M�3�n�o�b���� �P�Lc�! n���v�c�>��n�a}���D���(��G���'D�i����}�U��3��;K������Q�&�3����aLxmEQT義46��W������N`�hl���\ �ew!�L1���a���g�]��)<�cG��Ħaý��)�t2��a��_��t�D.���Q6�����̕&H#F�^�(��:��i*F�Y�n�����?������c�E�	Կ\�cb��z:��W,L8����o~��@�F��r�iAds�U	��̺���<�ʹ�m3V3=TH��n��@W	��#���B-�8C�S��nU�H���|����=�,t7s�c�f�4#U�^ :�)�C�+�2�(��a,��:Q�� ����_2�����c�2�U��zMjhHGd@f"jV��:��� �l�Rb���K�#�ƽ���"�}q�D	� ��=D���K�ߊ��3�j�����Z���:�I/s���e@i 5�0��}���Or�Z*���u待%��ia|?E�9?7���v����ƺ�A=uC�����`� 7�n��	��U$!	<D��:�vG�,..����K�.�2[o+����x�͞][�SNb?6��b��R'���w[7*����oh$���V�{��\o�'�A����em�J�ݰ�t���x��,�ͬp��D8�����Y�AP�ߋңi�e=���[�:��*gJ�
Gz�<MT_D�¬hb�qvf�qvJ���$��K�1�	�c�u7!Oa�7���o�Ҭ�L�~U��� I^�vT��8�K>�6hACWD�	�9�G�-Jzܺ$�=O>N�d!u	Y�렷�IR�h�EO+��=�-���nÒ��A��`"K|,���HM,�6ɲ�Z�ݣ�����	?�O�n�G�l�1��������!Ј�¨?�s�^nňV�s���[TK�T�S��l��zK�`�
<�1�Od�JI�l�U�AV�^oBG�jE�Gԗ���G�>�z�#�rK˟�4H�x3i��Û+ZP���	]�F�L,�J�C��߫�|s�(�ko���7O��P�~ÂT�����\�,�J��h(f�^��:2+=�����ub�z8�'�>� ��`6�8�[�@)��mwz������q�l�cry��N�^��=����}�mҋ܆�,-A��tC �W�#�0-�� �=��UG��ߵ�g���gi�|H
qV|P����ߔ�5���^�sЉ��PQZ����H$�9�Հ���/oi]�ˊU��������_�=,�+;;�Ӗ]hH���%:w�=����
5vXk��[�7��Be0��2Y�JoAy%�:�J��.������Ť�лd �B�S(�y�=�L����8�h��R���qH[R����`�V��l��:L4��1�],nH,���"{cN���W���A�6�T�C�`l)g`rН��9�0ѡ���;��e[+~1��P�F�u�1퀍��@$��֎�
(n�H�<����aZ���2����[���	1L��鬓嚋�9�-Þ^Y`��aܾ8�� k�TY��
D�^�$ f�~�E�.�س����$�6��~�T��M3;]�C(HB!��],a���(Ҵ�5]FM>e/�ì�j�ʼb���s�h�VL�~��L�4�ꍀ�	i�� ��@���Uj)K�o51�K�Ф>���Gi��R�hU~��S}�og?�)��+��{����G �:v�ޗ�Tj��k�S3?Q�''$
�&��Q������0K�a�B�׋�r`\e�����'0#�1E�Q�w\ch(���~�*a�|�Y�J㉳�z����=9,�5�_��~�~vF!קrΊہZ��ұ����p8l��.NH�t�%P�Ԍ8��X�w+�e���2b=��[ߍM�WJ�Ly
\��Y� o���45:�ƣ�+ܒ�5A�X~���A�k���hR�5B��@�o�r\�J �T"9\4�r�XWf�{˖��d}��-�[���:E�Sݶ�DŻ��=���|t���J�6����*��ș�C��6�dS�Q}���mHI$\I�4�M��M����n��.�gᨧ�'~W4+V7qC��}3�id���
�hwU�Xk���I��˒���{�����"޼�������>
�e����u����'�i�W�؉�@�DD {��w5�\d��q��]������!z;������G�O�ظ��|3��i��PY�䀎��V��	a�H���!��ք�v�_t0V����U�����F��Z���;�|����$��
D�k�6�3�ZP����v�ld���'�U4I-[.*�����|��dMΰu�$�E�h�Sѻ�Cxc���6�>!��J��{��{5p)̊b�^o�����>��y�{o�W����y������
��5��f���#Z1	'�q�ia�ыy��>�v�H1��2��� J �:��ᬀ�έ�/��S������Z�������68*Qs�%��٭�S�M����\6�fH �S�
�\�s���bX�qd"~n{�<)T�cl�u,�q�-!ޮa6�k�C��+>�uky4�	�a���h\F��s����pۅ	Ff�5,��5`�5�-�[u�_�����I�-���}&���V�Y�&�fQ�D�E�umx
���^%#��t��]�;0`X��=<�ܑ]ӷNk������	�_��fL۷�B��1��'�a�'���?1�[�!�I��w[��S]�~��6>�i�d�{f`�/�$�]@{$0Ĭo�UVX�􏏋^)֑+�u��ؚo����D{������,�MO�N�t!������F�}�Z�xl�un����a֔	��z%���%=��)�&d�b���������?�'�y�$||�
�_.>�h�ԍ�n���7R��5�g�g۫��89�t�e�_ m^�}iK�I�C��ZR�jm�u�H���<������p�����>"��9�W Fsy�{���h�z���� A��L��:~+Y*���- �a
L�y��!f,���G�^\��s��f�	�h'�>�OF� qr�lWREŎ��:0�$�FMN&(�I���n�y�Kx
��5P��Ō��5��6�\|�FE6c
��|��y�+�x��>}���'�@� ��p|�+�ETkB�F��R����ys����7��7�Ya[���,��|�N{��_V��:�
u�Oҗ�ԡ�Ό �~{iB3+H�Ϥ^2�� �VT���ŏ��o���`% �� {���c����]��	3.�E�����P?��c���@>m4��U�k�pPVc��O��,�"z�>��lw��ecT�0�!UD��k��iQ3�U�gI���\E'DA�%9��y\�%�+��oj+��� H��?�_�3�H���EN�Ps�|.�iuq�p�Țȶ���X��_S� ������
��.��`���cr���OG��c�u�/������嬙ta�J4�2�B�r\��Ct@,���smL�aYC�/*S��
Q{x�À�A>&�Q�+������7� Un��5_���x�S$IOs	s"#��^�4��9�N�zL=%Ǹ�ՇM�)ܹKѪ6oI�����<G�5�����#�����64�Y��7�9�`�=i<�HY��C���d���mC"���}L��(��=z��xK?֖}������ţӀ�v�P�(~�_jWj��x�M��0x�3{D��R0#}���i��!�]�n��#}��ܡ��c��s���!��N��}Y�Ov>�����m%��u�#5ܹ7jd��=?!i �vo�7D�(Ih��[ѱ�C�/PθTD�@��նY�)��	�|ڵ (�t�%�_F��c�
���^cp2���o�s���I�K���.�^�g�wRF��)~l���vY ���5���wۉ��A9���wQ`�V�_�%f���Bsi;���#{�88�ޣ]��2t��kD�
\���G.�2v��Y�K�P�3������w4�$�_�r��P�w�QӢR��R07=h�r�S%v8k�4��C�CSbPNם
;���V�K�!�uGy��&�1h�ꐸS��]��"���m%���'�f�����Ϻ�$�g���/y; s$�lC�#�\	��ی�����MzR)H�9P�2,�j ��O�3g��x���U���HJ8���,�`����M�Wk:E��y��S��y�]_���CB������N��xȚ�)��1�7���fϮZ5�̈��86���k�a}��!6�*Y=�(r�)�	���ȏ	�5����C��9���b���"S����߁b�'�F�[6Xг6�0������;��9T�1}|�Y3Nܥ�Y��saD��694�7�G�ϳT	諊��K�3r�ڼEFL�zs�:}�Mɘ�+k��%���v��|kNM
p�ҥ@�ik��0���õ��3���_�{�r&��)f�t�܅G���8�0��:eOj�$duo)m���c��+�ݚe�����ʦCF��q�U��V��8��;���`�������r���{�� c3?gdJ�{���� 0}�GN�Y~����@��W(P�B�k[��H1d�VS�	(﹆��枷�r�(;�&�x��+'�^�?I�䜥�.M6�}c)����!B`J�N%�Wn������D�|O �m7<�*;�Ͱ�D?*9P��`$�i��^E4����s1��n�o����L��`��Ab���h��8�h�4��ϻF��n���5#��@)L'Q�$��ȓ��� 	�*�y�Zq�d��վ��9f�!,�Ay�>$�U?�w��C�G�eX��`�E����%�	E�̲�c�8�¹��e��<�(춝�8�1�Ծ:��*)��-F��m�尶'���ݨ� -���p�2��8�nz��gYG�m;�5�=-���T${����5���M�i��i �E���6£�{�k퓮
�gR-b�j��Fޫ�έ�N��s��K�HX����s>���,E�,`�E�!^v=�i}{)	w`�:�8q�V�-�wD�c�>��2��X:yz�߽�F�AQw�3`�TUB��5e����jV��/f��O�4�I~p��I��k��Pr@a:f��l�=)���o��bh�\{�u�={��Y4k�*��q7\���KCch�૿�_g:�v��v�C�*�%�~7F���C����&�o#���E$�K_�%��u���l9�>%�Q����ae�cU��1�3��hM�֑Y���;M��G����!$;�����R��66tnBE<�m�]Y�R���sTz��q$�H2�UDI���y�ax�F��^��:H	�z"���SzH�R=o��-|V����B�047�~���guH�'B`)��Ѿ-��I���]�/��Yp������;"$�}RU1n� �Ҧ�{s��f�o�Ѭ�>��������z��
��]�)�w��4Ӿo��K�Q�����v�楘�u<'12~C�]ؿ���՜/H
ԫw�.E����4{����Dq��Z瓺��i2\,� ��Y���Y]������_�6	���*�q��  �ۜ����p|'� g�;�6�����{:�ш)X���y/���	g��pU84�-4�ů��6�U�7�8� �m������'Lo��U:�L�eT4�NF�͆�R7����H�X������:��os%T����Rұ:׋ք��������������a���[��n����xc�G�����At�>e4+R��t�I{:^;�!�1� �{�dI_�	�d��p�K9�$
�
h���T�Ck���b�X�j�Q��dS�_� =@C�y����D[:�5eE��fk�j�,g
�'�0ƈ��%ٶ�#��Z�ށ�Gp*&(���`/P؞����L�����L��f:�)x���"*�gٞ����/�Y�<�\4e�*�)���R��ݓ�j6��9��?0W	F�Ђq�q�� �߭�of�Kh�h�'q"�Arm��	hr���s�(T�g'�Q�����+���`TħN��c>wR7;fX^��%OvFLM���ܦ{.���� OuO��x�| ���������|�yn���-�I���蒾M����J��(�
g5kw;���w�]$�7���:m��JD_9	��0l��{X���!�}X6�+Ӧ߅�;{�FqrL7xik$�aH�x-��i+�<��T�<?R4[�q/*kc%�������b�摉�=/�JP�0����zx�@�?7/Z\t��^�Y:�('��q�Ct$��SnoG��_��`�ۿ����K� N�Ԇ+F�2
�r�bdG��qE+�3���m?�� �2�1:�q	:���8��&��13R.��&�����	>k g#ʨ�?�}���x��ѡ�}w�g�ʅ񛹷tb�V�W3���7�u�Г�9(gФ��^��J$�}���:�6��%M(7@^��v∑'�C��ɦ��P�[�l&ZX}$Bv<��)&�1�Wcd13����g:��!�2_Z�@�/{f�t��z )]�
��G��|U9ҁܫ8��\���O!���h�d^×�K��}�fu�R(�NJ��`��=����n��f��צ`j�9u����s:@d<�T�ڞ�$�NG�:<0���:����Q·i BPt\j��Ch�+���-C�nMC�ul\o"�%��x��9���P�}m�@��f]�;qN�<��Am:kz���ݫ��(b�o�)�6,b�D�-��UӾh�ltPz��@�>߮�yA�/}�x�Bn$azIGqs�%sC�XF�;t�C ��*�L�W3�fͿ��.��*�$����t�Ŏ�`t�A����\�4�P{	�sN~�N�^2�n���ϣ���zF�����:�D�%`�`�\�^�א�� �gY�ssY%�!\?�x"ႋS'����IombU��M_�����ߞ���Xk�U6@�G�|sǵ�5�}��ٞ�,��_(�UE��I� .-�|z֣�s@K(�'	){j-�:m��,��õiQ�Jd�L��'��tQ�3vW������j�A��P���d�K:�a�c
��~srl�	���ٍ	&��WT�|Њ�(��3�fڬ�}#�q��������!����`:R��*�O;^�o�}�fE>��@c�/z��Q��&��0�N��+�}w��O��87U4:�`�l�����(JY���+�5.T{1}�A>���[��-H��*1���u9ժm�v����!���C��yӟauSK�~����2�fM��S|`���kK��NF�����^5q"EМ����=�#��\R�Ҙ�	�M��Ǩ�붖�b��l:}}x*�G@5���o��9vq��5^� �ͳ3D��r���bao��2P��������ʜB�E�=p���p��+��G�I�{��;��Y`�-�t0D;7�T!7}� ��on�2�=n'Y-���u�)(=9�4,��V����^1ձ�A1qp{1Y{%o:t,���!Ep��|�;51"�؁���T�>���F���H�j���j�}g���ZuՑϿ�#���Ñ8^�0���8�v56�<�H�!��Ek�����?� �}Y��"DOw˯�ap�I:ܨ�����)��\_�ۂh�I�@{�uڋu5aZ���~�s�� ��駏|ێ���ݶ5�r���� ��ߏH~PI�|w~��3^�r��%�����ٳE�z��"�؀Q�%��^�K|���{�8R����qR~V D�<�d�ծ�VL��h$�@?��$$7��XYZ��4Aw�8#����ZHF	g���Y%�k��{ݜ�lԎ���d��D���m����:֌^�_Y,���~�������d(SI�k�H�'�|o&1+����֓��D�Ҹ��������0�/G�g?
:Ꮻ�/.��(m=ټǖ\��7F�ϛͧ���XϹg���;��Ԝ�A(�+xAѭ��I�^=�ח
�օ������wn�5�n�Fwr-J�D-Ș>a��Q��O��N^����Yq��S^8��Т>�
r�q8ps��Pܒ?ي�D߼�vs$��ԗ\~Gg��B|�0�B�8e�]kI�?�.h���ޟ�����E�gkM����X{��5�%�Yl��iRTѭ=��å(���WJ�Y1�W�