`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LbBTSFPZjL/CFYlyJT7KTr4L5iFAI6FD3M+34pNVxOc20oLZHikUzlGvuxiuX5Hp
RbkAEvkBbzqqp2TLbtXt/3/BRPlCasGBSafbGgZwIAVTgKlG+ZFf50OrF0x9Z/DB
9B7jrVuDRNY1Zs/O9c+wOL7fW46NLm8j7hxnJnKJRJY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11536)
NEt1Q799yXeYtS1QyC+XUKTujJyurkXBFSkHDyOqcqUWa7BxgkHCBFkMTlnyJJEs
3X50SZqSFdu9IBCRpXUj/v34jaI7Vhf3lltnMjevk/NeXFzNWMnX4ixnKJF8/Z+y
7/qmS/4yCKwqynJNpsk10bKrEGc320WcRU37rimWFksXNDeLjrrBHfKjG0dy68Zh
OQqqhKsh2ZQbE+PWbupZu0WsD7dQBrTp5x/U9pK3ozAqrGA533Z0gf6fNCoGXlOr
8OmS+laXs+7zZOHHAbsFspENcWSfRAz2Km2VgoTirppr1GLlO5q/07Y5CQzGFu2B
uAbq1SQMXbuN4bl98b3HX02yfJ1nwcTmZvJJX6dxzY9OQdmSszd3VkoqF1t7W/zz
camcT1OB4gW/4sU7c16QHkQc+vkQREnN31qNLPgEwV+S2A/pQo2Ns3qrfQq0AVEC
YFWlRCsQz21RlkccHLCmp7xlDgQMlAvuSxr69xnuuhCLK4XkRVRB1CUuD/Y6IKBr
ymKmKfzRNoCGieLrQrWcaRCLLpEzsPG6sKIg6vc9yhY1bsoRcC6HD5xUrtbmrkju
dFiURUhzOFtv/aW6xwdf7B5+ROvshuSIS2s/AbvoBpH9g6OsAFO5rCCVPTQups/5
1BPOXaWBFQ41O+2nvhYSLIwnAXAa8b3/Ftn9S+w7634ep91mQ3KWIpvuXB53DgMh
XjDjHjZ/OOBuccmcYhBci7mJx52PXd9mr1jgaWp5LPfULyOVdt4oJdNbMWk2dzzK
JLhasx6lw5knaFvcsjU3duisPpxWJ5r2tNP89MSkKlvqjrfQmwEfZQRBwfhE+kLy
fx8Sevvml+esrGiJaAbi4+yZqXNMQtKx69c3dDqe994GNzLFSzr1wKldz1Dum37E
rMoTj+Vrne9yo5EWrTqvHZISe/g7XpIgBD/u3aGHVcfIh8rtm8VuGGSl3VhzJTpc
qWCXXnVySaJFCe4A1VQn41CS6Gc5qcHLHSJyLmjWDvzTOWwj46oDKCKmtwzw1Q3Z
/vqbfxI9CkCsAKn1As8NxaIIdWTJfrinHI4Hz/CTx74qtriWgjmNyhrFSZiK25fO
nZDHE/p3H/PkhNPqlIe4Mud0JZfljxaJSTONCzWod90QVfNQaq5zNNe4HARUxVwF
tlDiYonkpQkclMYbsizPcNuff6CBMlS0hLzOA0t6jz94GvSDGJkMTEBqPwzouURd
DSdOULfepiY1+TKy8C5EVZipZghVYDd3nWyzhEOMrBYZAieRQObzCNoMNbX2XNZW
HK9sT4LkNFwHShK8x+kJN7zSbEHVxREfaaQsVdbi8Q18iAdHaNm8VddN3h33lBW/
P8bH+vL3WGk/26uGFJh5qjg3Qt9ZL7eEYxMtSzE996wJYaySV5ao/XBAExoOUjUX
AoKk2a+frBq6BdWly3MjdqDSy65f94mznsZEyZ4Kbj9DewmbVKkWSM2gCeAlFeT7
ZwrDjGpe77sdvbsldWup2HRzVGXXbfFl+Mnb2vGyr/e72fSK0Ns693fmsp+Mv3jf
Yha1wztuUFYfiwfiYa+4KMYyrTBYl3+VGXEzZgR7lUoD2ntrm1UlX0VCDIxQ8Io3
VMCXQxUBQqQ+MxEmdDlOdrZZnX/N0SjA6p1XT9rRM5Qmd7b+FsZzg0CrK3VFJlrG
cNGM6b3g4YcZEjXYsEVHkXLo19YfeaepZ/Ds2htf1+jdZCbz/q49naF+hoXsrM3y
3hQHy7NGibpfoRO5bBAViIO/BJJV089bRl1hslYVB7ld9ASQX+6OsKEBjrrLh9SH
XW43LqQHIX2oEwD95t9y/qxvNFL/xSqe5rnDfKJdV/BhW44ObOgnjTvuakxYp4CF
q6XLJlU4EZkFWS4MGG9Ca3IK0P+eM6pry5WLjYL6yFRxKG0xEmq1DbdtkmPNMGJw
d4CrBFhlpkmQt1DU+N3zY+atOkUSb3leRyiqYlBMIFYfJJZmaS+Mc932nDurD0w3
G8YMLHQdP7w5MSXb0aGw4FIrr2XOsjLeeY3iG/hoBvLc9eCPbMF2xcCe2e8AHN79
6i2cU3R6xtGiOyBWcJ4RqzDznzkSxBkKd7NFDPLsnICCnsFznYQBtpeuCP6gFqib
nHGVWMLa7FZfw8H/CSliCstblQhN47Un1JZsRUA8PZihJffvmAC1htqeFxs4A977
cmTRZ8kFVjqKXDwkGlLCWv2eFLNuwUMTj6CzCiML8NPkF/Xe3aw5filYNGUaw0VJ
6t2J0uCImheJiAf67dlVi5+eCMM9tZ5IqZ7JawV+4+TBeeUNeBioDAVpz39yFNwU
zvx2IlUfI7FrsjbN3BFlv2a7hh4moj8Y6+sPTrMB2lQh+qpJjnHyhxhtaWFiMrEv
VbHF12sXtzGDiYHud8We79OXCj34/yIl2xlppHE4N1j6DJo/nozsaA84Cg6x1Jy9
RnWDChDJ2jkj+B3Pkpt8CzT8EAoUwsOXkoLPszysMlQAJiDcC0tUv52BSPjTgd0e
lGxvUAyXe75q9NCWp1/YrBC3fEk/5hJIIgnvy7OApb9Inuzi2As5cDcHAPJx4MWU
rVuT6nJqPgMfuSrj5R+kXkHQLf5jA/AQsPjXLY8jp+9NOV8WxCRQ1aKK7Cds3IWC
+pMvVgPc6weTcb66kZ3PCqBh+Y1tDH3BBvf1grVSRw2S+B3/zJTteqm9pCVjFvX3
c2i8+cBHhgN7h2h5l4o6YpZCA1rtXm28POSIXkbTst6xoPKyVSLBLvkmoUGkUU5L
vz0ouc4tIqrpYnxh0ebSAyFuJnXjkmyHfFLIxPgzRzpolnQf2ON0oDfPuMYgBA+h
4wzNSaXlujrNNQom6kEbRqjxXM7yE0BdFMn0nf7XXrhWohEU7w/9mOfdkO2JLNIw
ucI0njw+NvDPryIhpWScc6OBznFeYUkMNyl+wNIdKnVx46ye5kOBQMxMU7XkSfo7
rXOKG9MwKQm1XHYzAyqkODLy5JJMwOOXLk7AtB9qKSRIHvYlqMRAdgH3qO0QdYQ0
5IuLERaDViYJj3O16hC7bI4BlNwwkenFI87ZMeFRZTozyIpovs+OSHRuMCJbgowg
7O4RhmZEtjnu63xkP11vQT9vSwABpfQDgGxX47jgUD2gcrj0xOApHci1uwPOzwxM
IbF/2mUkSjKczmYgNG9rHh0rxAHDfOEWVEizRHGiQhRiWVnljcHbrK1KVp9m/ZlN
ygHSRrYGAHtpoSaSG2vqRWHgX370X5yeJuZRcc2gyVJU3IFL4CCLysLd/LdeuLN1
SE2Z/2v7/IZgJfkOqrtuE29bV8O+3wuPjcxVf7xcnQmk+8Ek5cMbY6vhTzS7ZMwd
crlQbVPRlKXtQQ3kilEkZBSKtWurJzgIWNdlUGVo8hSh3Z8pRNjVlsOAzRIB6f8L
uCYIc5rO1F8yphWIzcf7KYSBXyVzJup2j2Zl26psSeFQDq9SP2gPwGMIpXBnn+1z
xOAbVeH6liNltg+YfXSjg81z57YXmBRhLyz2PZv751+PqcCnDcdEm0ZJSGKvJg3D
esIoipZW5Ef/Xl6ImK12xCVtWAcpMVqdDCucPJXgjIbSc6hBPAX0jdM5nhcnVgZi
Rqn1yuNVnd+5qyehFSA84luhKaBi0WD79mGm8D92KByNewvx5Rk5Z8niI+2TkcKE
RRohRsc8zJjw7tUqJrHwCtHk2YcoDNOnEsp5EiJBislTQigCD1dYAXctdV3cScrt
zcgUaeOYmrJ0vUzhl1StItiVQEpoGqS0yZGXUK58Rog1yfU/Zf5PmeIbdW6ha6Om
CexIoTblfos+LY6aan1JipqD0inOCh6mhNY+CheicpzcPN+7m6nbCiRGQ1iEu3C8
4jNsUXEQODqVmoHtgYHIq14Ps1RxE9gZMsVweLyaINIjd4cDCWFayBYPrwK9jtBI
OkNU0/g/c8Q6BpKjBFMuP/pKeXeHJZV94GLgURpojlA3yvI19KZe/yYkRWhBzIuS
tdFGwGkxRFp3jmH2w+01SzVjHID0Fbpw9DPlajeKNvUaUoqZT6C73WBNjKcVRKjO
1znWEsWuFkktNw0Z1Tto3NdxHcK7xxHaVtadmmjIJCMtabUfwJl/b3PyRTtOxvfg
d634wkASyVH0tya/xt6D4wEE/YdJ4j45wtr69V86kv4XjmX9d8FjrDUYf0zSK7AX
dZskrzH4aIi4kKGhoC42syzLp5YHPkRxwrf7SmszeENUno2O/sDHsWZDvQIaJDfe
qkn2dXWzw1jpoCAUtB/4V/bOKx0PPX4MPCjvpR/LtcqBaiDkH0F2QNeXEqw79PLk
tGaHN/invgKCmd0uc/2vUn5oJSs5VZzL6uGxImAmP1j8hv+1Hg6gfJ6EFxDiJ7lW
hp52y14xF8x5JTeUlCFmvxCGqFM8VpUC87Pv8hdCPZc5JOrF1XmsOyw4/pTuw/Ae
bgn2/sDRtGIC2OmSJRu48JDzEYwcKvXbGFJeRN3iuk2zXj0FNp9YqoCoLmZHW88P
OF21HX1VRfZKQSnLdSqzxGONSWBTGvsRFs37edacLTRQCya5yGER5hA3z8gnkENA
4MGhftbls4rTjoqQU8U2Z9rtVyrZ1aH09mN8iC0lD52wIdoHNxNadIbLch8EsErg
1MfWwzwDzxQ/TTq6g16TqDr7om9Jo9SAbkf/L/DfsWzxkl3GF8vm32h4BqC6sN4f
ug7CbxK8s1VV5CfTczM9pLqmV0TyCRPzFHw0LXdnbptKldi43JiFrLyGP8e4RQm4
Y6oJcaLk2jCOrnG3tFDtajlwPjf+7ksVeK6qkAEglaa6N9QktF8RD4c5BBZVUnr7
sazLVbP/Dd2Lrr+zSTncdZN5TK4eKpy7XtJjIB+QusiV6RdR0dcWuZ8PyOLlspFM
XAK+tM4FsTKssHZE2BN6UGpYqjl8/R1wwH/51MSludEtGQryoJj8cCS2BUnQSi9a
TcyfYsvjbo/nC74uIpJDpJTixckRD89kCOOR+Cu7btyrdtr8FO1q8xk1GyAgw4F+
G6OY1rFnrs85sTgvj/hliw8lnrwCvxjEiqcaNFYcAXAYzAfFQOdoARPfpzgDekgX
4pfaE0XIsxll/ZPqjY7KvNcTHbJGruhkzfF79o3UYd8zR6jplh77CleU51/oeOIh
C7GrcZDZYylntk1bNsrbzK3kHq+7UdwYdGNvh2hOernKdzhevY5Dm+NSspcTTv+t
hLJYIOL1OGxyhzNeWTiHrQ7OxVjbN+cPgmUf+Jd1/Py1u8ZY7dXShCm0Em2ub0Ct
xCkxcxAWBDkkDiQ5mZIFJ9iWbS/ZHysmr7v4ANtLFUB9eCi/dHrVyZtPqzrkY3Og
X8XqWuvttN13TpENLcfhpG4q1ZRPEJcIt1rAnD/wDxwCoG/gQxrGWorTa7oBQkjw
wBzKriJ9ffGQndM8yYM7dTHF+oB/zF5s5CVRFmCSL8m/O26bSmcbfxxetIN6WHj8
m12BetO77U5pyJd/ho1lBehcIqx433+4N5UM+D2LGt2Zug5n2sxQAUR/yAP5wqjG
f+CotaHRZ2AL0zAAWFNxirvvgeeo/Srt+3XqB4lQbw29ZDeuljiim1hCNslpc7f2
hqZnWe6E97mEVRvNw3zh4QuRr0a//IEjRuYK6hHZ3QuTSAkNxW9SDaigaRp9YEXF
bDzsiXm64ReT3170d2Afu1uaDi+zGd/F5fqIzo8fYbulVZr/iv2mdx0EV12AP3tf
+uw2snxIqMstRQJI0nXVVFL/+elmBbmokSuKJY0u1bS6QyCSMXS3aLz+qhG18DHH
Am+fRN05+/GRjRIleRes3cNGe4H+qZe6ZKHYo5q4B2TlRilA0zNy4KCkAHcs67o7
N21+wrcy8WToLqxF2/c6usXTqGPefUG1qZYHd9rVDZs3Hg1wFtSSFYmVRolHyK5b
+JTiQmLKCnXhhgtZhRLe8+15oWIPHtDVm/yArqf+RXmr5lV1Kb7R1p7Clmf9KSjk
q2Ni97YpfVJrkntCkWkSV4gIWps5MRaOrF1UmNTFKNvAHhy4nEAssGClSlPU2Wf+
Az74yhGeOw4MbNAUcdJHssEj3zZKs/gclbacnQD6Vjrb3m7fht2bTeS4FKMElV3E
glfKQomMLICTk2HceRR1WXrTYFBgJb8wv9jkLYoWJXcZLK8sj74/Nf3aGTU0UrZN
nEeLdgrZtYIsJBJxo4q2wmfgZk9NGhta0fr5Tb4VEnAKvx7rvQ+LO/4YNdKSTEOS
f5QTtTYALEFOFaju3q+HlyduZ4YMgl5PvJ7i1Au8nUAj5bLJ9MwCHr+UdWs1eUwK
FfymWJJhU0yoGUseYWP4ya2yEUX1liGUl6IB9g2uhkuhhWAA65CmFMepPvXXh95O
7p+hJiXdxH1M+BS466r5U+Rb9i9PcNJ/xiyDA5Qn9IinGKBeMUx+dsf2h8E4s0Wt
hvCuM3mKKa5NzPNIn2RjjSlVCuxItGLQ37/cSGbcWJXDiKCmnJ4dRSWFamY/wM1s
x5Dq8ldnnTxucd0fFvMLkOj3cA3n6VHSst2WnXClIPvmeRoD5NxEFZC0CppcEtg2
OmEicoMDwyKEJQbBYBi+0Zn3WTwLIdPwGj2fYoWd923pcfaK7uu9cDvfQZ7tD9PK
G0UPO0sDJDRCw77E2je6ItYDe64AalfVKDJRZcv8JG46HgKhHVA5I5fa5+eaFrL2
2aQOl6wJFQJcuIcTz51ePinT7UZ0VMkIqCq5xxl7Ed+peC2z6Lsb77dLf4lC6bUL
5J1hKAOGhqOXMri+fD4OMhydUkd2tO3Kh5S/1Db9MynLHvbKP9C89/9EtPHntpE/
4xpAWGDI+Pt9wEuJ09V9hYPyty/MaVOim9VsiD52+hRBtQaM5FR0xpGCyddisa0q
fy0qm4hTSavjDo/eS39UzimfDuticXEIpw5dUdYE79ExIE/xU2bF1D6yVHLwelUa
MT/8C0ValrvZEGCNbbKisBz6zSvtEHbR+t0onCLvgddxfV9sDMCgKaZGnd8OFE9T
3FvZB6XD7z3gpSWrS56OrVRF1NgTFjGT3RJuac+HnHu2SqF8LXeRXnfgcx7tISEf
uGQkmwDNgJbxXIohunwnwl7QHn6ORCAXTr6RG1xhfG+9uA7OQmm7hQiMbwBjv4dW
C50sxG1qcI7gcxswyAxnxg9gQjCoQp0ZxsMDHff0qRY401uyd1ptQ90a9TTpAH8R
ZXUbq2FB+mh04rj5+eBWrpFTZYllXXAztkFIA9xB1TKWELU4tA4AlwqUrJhleu9l
KWt8EnCcJgzjaYFbP122tuR1heA31fEb666hgUMWoxD5uL9xhn02h5mtp4wJwq8y
h8eKYEPsSMNkjltcX4eteWwrVC7yPpqs98Tfd1oJyhbkJ25/xITcw5rc6I2kH1Ph
gzhX/HaSCrZ6H9x3hHJ1IUio9GUiL5TsCK7kvhdpypxa8rytlyIpTan7jIq8N1l1
WLTEjv3JewB+rrqdCkQpQkgb9aREhSThanQBJZr2aXJCkeHXGVf85mtR6AUpDPZH
ACcwmD2DL+EQyTckJ4vw/avA3rgKph8X9Zv3qnxd2bmfhhHX6M1vvoca28y8MUU9
mTS9JK1MPif7tAQKH159yyDuJaLXJWf2Oz9GW5JcpavMALivxXDmCTjz3LsWrrw1
xI9WpHjOWLhNYE4OHY095UrUDjDlPRamFVaFAuXdtwQJ8g96I/TvYmcEYIlsBvBU
f2PpXHpKbOKS7zlvBiQX+fYmA6q6ECgrZu8ocfwe+O0EOJSsa7lccOqDN0xBg5HX
pytmuSUJoGHLqi51B9NZ+euQKBptdz7D2Q0yQ/tjDz7DOM3gprHlw7hSeA3+Fs5o
wqZh/Xp1RoGs0IsrhZ15ZXe1kpBryxijpjdg93AVUuKLFSTxi3fP1Whn//+zkZsN
GjfbFdp41EuJf4x+f4ZMgNc8bRP1cogCRXcE4e3MT+uYMeBjv5c/PeegJ6X8+I8z
AD/rNMoO10nBgbblazgYBCraLvGd72bq8l2Mz8ePwBwBEN9V74RQZUjsfSys0+xW
avTfFJyv5f/v4AkrvaJdaaHJeWQeTp44IvKF+iZV1vDS18KO2cLhF+F7043q8k8R
VFPQ80/tzOWCVrVZnjyMu9x8wWXIhIy5Rw0SrbIN5r17DFzEgyx84gC75vg7p7by
3dkybPKw57oAgLyE86BtQ9l3HJay6Io2aWTOrTzD983yCfrcQHWw8HdxmP/cYNr6
zSWPypJIRoR0+0gxxm/X+RVKw44KdJEP3RBTNSALUZ1Is44owuZzMM0kwpnIj8qh
pnDRHRKdXmoBoahNYZiOuLfrlCeWo6jpQ2RiMq4jdN9gRecOjVH4B61fd5Nznd5K
f9XHw5+xyvpdlxtDqPhwAUHUYZ11PA87s+CB8y1rX2T8i5u58V9SsNvEad2odl48
fAZDN1ZweWbTz3aw2kOmNOD6Og9ijmAfLUZzkb/qF7dXsb12HyH1+iylabtIl7sd
8Fw2bOgxpgxwcRPhTuxnsFwfBnOSQ2aW5e2FS6/1cita3vH55Q75KRRLK2cK4lM3
G96Qx02upWe9vRxleMUsaXDAcsVe+kyZcdTaLpdyXCn81vJmC7Ej3AnPj96mI5+9
uFf8mHJ9LXx6+BPg8Umgu/fXqKdaLSbI2W8flNMfeNCAkQr6dij11yfAVFI+OH3H
b/D9wnBuYgdsvyA5kxSUMZp/xrPiGbwhfoYd70hu0siy3MCvXDjhPfmfuuoKZ2d3
7V37C4dzU06cGWfBfXsbjdOJjoJEAYc7UczQ/GNaw6kXA7dp95qJt/8VvX88kFcI
0mv9D2GULMyCgx2KgoVcV/ctwSJjUzardNcR1PKFzMi7byIicRllzzsOsy/AWES3
S2rmUVjWQFpowDLKnplkxubY9FSs8X71rj3CiUp7TR3wKlHNmW1HY4Bmt4PCsrKB
1mZQj8Da2z+vTfTpfh9/ouydCND1U9qazvV18ZPmI7eo7Sj8F4Qxi29PZoFFEGnP
88NkVGBpi90/E2VkrN5vGVvnDh72CpNx0lm9ohg8opgvCJ6zh5INT8Mc/gXU9PZL
VDuncpl8BQ+gve4pitMg3uCvkgFkR54bbLvM+6kmhmDssJR7kHZFvMuOfpIohOJr
YQhaUh+t7IafLXWZEhdG6o22jgBtgAKs+lV1v9Dvbl5ITbXREH4nxXT4rbuJE+FC
wfXNK/vQRmHEVee4te9kbNDxWHCnJpW32JjQenvE9eSD2uSBIDD0TnBntTtPb55M
Hg08tjKUTxTr3OzG4sWZA5auJpfyj1/YLm7MG2NddR7c7N6l4xy2k1yjOp8D9IBf
dGInafMiLTvur6zmCjcB7LRtZ/V6oRGgRJNT2RR64BQyKXQ4qVHvTsW/3MCZyjWF
jR3FseQfFF/k4WA8vWRd5dd2cU2x/M/HtHbkP6sg4bs7uEEMxXQX5+75chAkv/BE
f0Q+TocpefugEqAwhm+MQ3O19IovA/YqPjn+qdrjjr5hzV1zpYML4tN9wIzrg1yD
y0kOo5ivZESFOsCYEQ8jaWbs5+KWnEYIsKyJuvWsyhCyD8YAzUFjyyoTuDHJxsat
L9/NJ/kEcCCBqI++KFeXRgz1yJekH8pYYpSpzGb+uVd6KMit5rGNvlUI/3hdQVSg
Nqm4MI/7cuRWZs7m/bBrCldzOLoO4HGO+LmVVLV04uu8eLhGyhGGxzKlBAWYIUTF
Ms7wwIO11AUrTQYGBgbR6cyr4w9bU3F3XtuuKyT72LvZxB6l000p1bOQjeCmeKn6
V2jzNy7pM4yuSQ4JT3j0VzduQ9hvC1y9/xdymyqN2SSgKSHPfHIfSiwfJ+7v36G4
9548z1Y4NXtCUjPEuPnUw6ii7g52dZV1k69wClVyBuV1w8HqsKyaqjLOqBtj++Z/
eRCCn0iaUNsAavSgugZfJUPZZLvC5FLE/PgU3cb6YJApasd3iJFi5LTlx6cne4Ow
NLwEoQ7iAVliFh2c0FLxu7a860YlF/c+WR5vvcJwuZjjqeTPDShj1lWc+MmxmIAU
SkzqAVhFieC2GD3S2P3QvlzuKxzmTN8QOhHetBaPRQ396eCtoVAgb8qr9ffvnxwc
BrHj6nvrTYlJTsxKZPhAzXAYRmDn8zKQOTIN/hj3CdDodB55Hxy5zhknBSeJ8TOH
aGF+b9im/PwSq43ej/WUmGTSBVMTPIWV0sHK+NuhNqt1xxIzfFERRYBU98sdCw3k
KxCgGg4Mefmk2blFBuZi9POv1NtEVAkI1sWhmFTpi78UlcLmsBvGnPCjoO0ieoMa
hVtevqkKksVPEva5lrXQRA+xkms2Kj5zuV3CoWsyWDrY3X/7BnBXi9hvBpUaZf+i
ZkY1ds4VRSHJ6Y6FHbpNQF8xRSbUSNLtD/g924BGMyjYSHySk0I1Pd4xb66/mZBQ
zzDsz83Zl9OULbH+gVdQm21IjiJp/qdLf9FdDWfcLPgaCBhGchJF3k/L/V8l5GVR
8PoYTWpxbLqjWRZddi2IiiH0qlIosi8psd/D89pGRLvcFLmBO8MbPdQmNZ/brP0v
bNI6o5c9rBNfEwzZDE2NcL/MmKSZ9G1AgLSVN+vBgMjQteJVMfBOcVkiVje35O+/
PTcEeoJ5zNAxdG+4SZhwMAWm+UXkpgqHiJJHfq1NRRMOntRPsP5L18NqRiYJ7s5u
wQKgQPNxSCm7n4eFtt7v1uAooC6SWf1oYZk5e3mIhOaziCDkL/3+uhbCfwpQ/CPp
pxhrdEixF6JITEBux8gOeHYkk8saITBgJqbIoJmxSDjKl6kOojk38gAipzHzNWrM
uHFzs+FdOISvzeEBVVLcys+zQjUAJLI6NNmfr6xCzIeIYtjCn5VllwJSUPV0sJhl
Dz2bAekV1H6HVhYqYuqUcErZChlQdLXyf8nO3VqLyHQUC/hm9ERb0Z+t1vAVsytr
Yhah5b0iY1McvIIgTuTh7lpNdD54runS1EtwST8b5/X6+C+RXaLqfXDqHEnq66iF
YFow7MOfCQi2Z4/udhen3YXG6ixDKIJHHHRr4uF7N9lKsFywmk6r1mD/XDDUrmOH
X1UEkwjeXQkmAGahsMm13mph/AScfajK5L0t9G5X3IatKEwt6gBMiCk89KXENFlF
BHdOpgxcmsNhSSKgygSxtYu2MzGDNfOXxviwhbYhnbZuOdAXtI7va1tPv1uxt6Ks
BfbWRfzYjj8mOFwNsmgLqn+TC9WBEDjfTCDQ/sgfPapa3DtM4+RUZtM6n9NawDuu
uin83sAD79B3gpBfoqrTXK4tqY/wbkJh4mVQJPbdf9r6YkdE6iXW5rkSMXP/vxcr
IGWsvK1jDUM2vymEokkg4/viAmoi7XBbMbVxZDb2hptDo+NgY/zCAi26LttGMyuy
DVdLui671jBf8ij9FO7EuofQE6b5xSyuspWQjcj4WuRK6lKDSY/58aV031PQC6EK
Pe9HFUrWCNdIlhAkMQSK36nXItSkHuw6Weg1CQqOzurbszN6wDdSMK9cgfZH5EQ5
18oAK/FvL2Nm5oomEHbs7WwcEmWyhy2Bx4SLFXqFTKrLf/D4kPoRb+qEO+VMwepP
8qN9YPl79/NPAuDxVDSreNshyCwInxgWF8MbZl6T9foxbkVwm557Tc1GTaSpCH+B
BjIHSOE/mfoLK4F85Aq6Fkl3mA71a/NCjup2gMngA8ElAxChFTSrCtej+pDwiLGn
zCp86xz/QDO5AN2NQs4hIFnh4dXzoa6vvWgU8OZOerLSMLayWHnUh5kgP3BSUdcu
Vl0PTW/7XodhdkA+viX/i/Q9HexIHXh6fvZcAz5+llrrf7qU8aTzIAmM5jAlEFLb
5BCUiQ2YjA8epMpBrCSbUcThdTxfhxvvyQKdC4dLQiAZhgGbMdSDzSv3ppod6o5E
xpNb46ZnozuEJBMDNQmlMYRZfvtS2rcHU1V6ldjy4Gh9hLAzDJ1jZuHrqPSmPl7W
Hc8aw0VI9Drt4lGcLfrzu6Y8OevYt1uSN9K08kTN0mpiozyBEyGjjn351PA2zF+W
gOIfRtDod9KizzSrPZNqp+Bj/GEB1gNKu/sWQVPRUWdzEOpnn38NRAgx5ZAQKUIO
FrldlRPsZYcUQPwqhxqT+bJpsgWSzIcj47ahSMs/Zu+lmonejYV1Bk7kwoA+3soP
WIkT/S64IrjKtK9mnCPuuJOeBMCO98q7nLEO1LKzSW5Ku9mpMHwjesRwDmgQikPj
Wmi0ya6g/HA/njpMwAH6DDEXnS492crr+/zC2Rykxv+tltIIRibL9AuJdVcMcxVi
G6mZV7rOG5xrG2mKuN3cQmJkeZH6FjCJBLXBeXYExlbIe8H2P45YBh3hDrjHk9+5
5gHp+ukn08DNe/ZOC/jUPe3j/bA2W3iJ1dZhPlT/70pzC72haPtilqhZ4HelwKyV
T+Ag6TuqSe1k3QJx6AmkIMEyRLBiPnvub04WNevSsCF9TGLYc5TfUvv+c5ULWH2q
KFBIA1oBR09aKvkUjXxG5QekQNBuCoUrCLDoVuu8E9T8LtVy8RsDe7yjTz8RlIKk
KHB4NGrtL4OwMHeVSma0fK1EaSXDqbYRNiNak7QNn5U/E3VcpmjyHYr+K7qG/KqG
lS7RHua3U/tCRflbTOFrvmUA/f1IuUQt9iDzMRRmMIzjQpKjpyxGPT1stHvuL3xI
w2QyhrQUyiD/p+nYgbK1a25Jmk4Ull1eY3fj4gscyM5E0So6CTGVOkGqBBdukYTH
twEdJrlmU9MLIp2okxaJB2V/OIpQS6DUZIcU4fOdpgTjmTCNBgunb9us69Si2IB5
7Zu5VsdHnKsmwB4TAT/ZVPAfZLNPXIjrkPlvpv5lY6MzPsNTPdDRegh+QibxSZAS
2cxWLDCzqW2K4pnIjSt5iOUdLM99rY2aCWPsFr0bDOzhoWIcdNFouHyhMYeBpnNs
tvvTIKsuJ5al9ULTRB4u2nmm8QxsEo1IOsz2+Z6qGipbI2eY5lZoDr8NQxCdSryk
mCPH0xbthgbEv9dEmuR++2TGt2kL1vfQTGMTsX4mBHJ8DjyWn37RBmUosZ125bOL
VqWjFn2/SfP7K1M0cJz5vG7Y3VuqNzHz3Qa3dr4whlE4LrztVRM57V6cslgRmS5H
h90I6ERbm+oPbQtbuXNj3Vcz7eBPsErg0XOKHhRd68/+ZGkD9hDujEe5hY+bwomm
xcjpICLutZVKLOUFelDsCWEm52CirQ+GiStxB3nIVILRyrii6fil/OhWwt8mzvbj
zxgYsNiIYxxXokPRyNsfK9+YIqzVNYY55mpgSQbkMWjNHuB607Om4BQvXIAWPoDW
pVGn+ftY1F4LCe3dblsTD35MWp63xYiUcM4m60kKljD60LY9ZfmxI2BN6qYbVeOj
PUQLxg2+QSbkTp3Meq+haxzZ33PMytggQbWAgcMwzg0FIEGvf4O2TgvSR4ojvwQV
uYSV0umP3xx35qIAbICWJBz5iHublr3ekBMrfHQP4Byu8691Tlzod/izUDinCyAr
t1FaYy16owcYdvZy5Pvtc1JUu3KeMTYqbMBwQrG1Ke5VRCUd5JO+4X0FeZXVZiz9
Ibmo/qratvPbU0EmLfM52piuUw0yw9Lf2xWLsn38e3Xk7YM4/JbsNIxYV0ffeMQ5
D1dKlFecJZ3PSw7j+FW4TjJ2VZClKb103QDdE/YvihkG88PR/UF3KVN6F/PjOUxc
+Fyd0JFxgHIYcawioMvDPTjFRz2kpSgoyk9AC4JhQ5e45FGFgrYNbJQjiPS6uMb4
9TUTld6FF7S19+e5P4+XTnaqTBSC1E/n2k/9w0rGYTpr84L5RpqZVlMBze4C7pLc
bgWDkS+SW+Ro4ND+MojO7SQrhL8HiJAAd+P64GMR5AZh/DPZq6B2zSBJmToAlXkZ
sYHDxQKTNH70HfagLGlEHKofPisvQAk5OPAxolV5B/+JNyeoSdr7FlTfzD2AhhFY
xpnb5Bce/xUTYC+jTmf9NUymM8TOYWVb0wTPzAEokJQE4QLMdD45sfHmpdsJQ1Na
PNFcF5+gID+XxN3vZIgeyZfH4jnsSxWV5+Tkq6x502lUqL9iHub7npYMgfKL88SH
cAoZZPVPpn9V1xpxU6zIC7bbd84LsBWy0OKcrTqBnI2oGxSvtqxsd1/KNIYqPtDG
+elT8ohWseFd+m0cRCsDOR55PqndNqgpdiZHbFFkQsKr9YfMKOWwVAiq8A4S4tnQ
Nyc5+X/LFVvPrxf6GoDnPUUmz64UVCd2BB8KiIlrGes+X3wQHgs4pLjzsHgkRTQJ
SwVx3u2N6O0QXcCR9Ix9pPbl14jIiKp8PRvgOypKQoXxLSyYM434n1iL9pF/9W7s
Yb7rH2VMS9pKbzi+BL6SKsDxNW0jhtCmZpyayNJTlJ8zAupLlKNjroCAnPu7dRLh
w7Sx3UJclQA2GR+DW1e/+XJjqU1BrdsqPL1cunJ8SQOENdoqn2cS9EX6kq1hhi0T
MWdKxhjrcTwshLG1XxYL7YmQZbdYfOjK0t8mxXkG/zlqcU4AI/mqwz/acIwFE1cA
Tldq0Rapf2Sk8JP/4w7FHmAf+PO1tsLrNnqMAHz0Suk+2dt4RHu5orvus0v7yyCB
SGPO1ouIrZCwNUi+89mkHh+EhxyAj6GSmeoGGS/R8U/vGR2Jm4l6csFIVnZsU2Z8
prYoYiZNo3BCrnVhSwH7notWF0pVg+6Tn+gB1pOY0YgbpkEGPfJjTXeqkXUisoQm
rFf4kOz7dkf7AGKsq9Shs6Y6n0oUHvyVODtU6MMplfcf3a3a0PYBmfwd75VyE/Io
GWQ/mAzVY5Vkqd/t7y3V+8fIMo0ZPhPc329N6iyoRBNod2zygRUHXwzI5btNwkWy
Jc2Au6+Dfo+HwedUtNsEnB5kdLtCSyY4vS5v2p2mIjsk9POmykYan7g8VKAExlJs
RtpYtMJeCMwbx48GzLXWd8xUDcsJ74lb0CLqEwLiaqrcO5ppBjDR81DWALk6oEvU
wU2nL1tUTvT8rEIYXSwdSEESd+9fNfiyQkzJrq4NTduymt3Q8A95qHkiEmOjBroT
jJukWegTaRqkD43Ni5yyfD9MPtTHRB1hkcTnu3sRAhZ4n4OtHBezsjCockkqQs3B
oRhreK4o4KpePAvEGdlSjK11zA5nqzgGRRuHfPtralqW0IeD3wwOxsHdL/0Cc1eL
KxzJMdFZ0tpXkRthi50e2Cr9qkZJNmwSqhSGFdubR6KHf9MsRw0zAz53ZtoEgDCh
AcQsQ3AJl0nm1GYtFU/VRtI53JoizX8ALftwndaLQ3hcwrTWlUmg5ZQ3Lx2VJYSV
FRDo11a/H0a/X5tz+I5c2FfDrOPympT56NIPzkFjhh/F7mfQokJJo4KpGuNbS97i
7A0fOBybNbWiOHIoovMmyBr4m4CCE+q952kkl17gbCBK8Um7QkRakcCxJPo1JpEB
fWXuSKcRZyhsxsRY6C+O3A==
`pragma protect end_protected
