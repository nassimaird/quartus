// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AbKBSpefN1IW7dPWoWfcG1hGR1OhFzRXbP4HJmbKOH80HDW57v5b3QCgx7AgH4nTTHOAgC4kft4z
Jo7tBvluAW9CgnM7KAY+xqpj8VWCD8uh+v5mVcVXTn07157itbNol+VPyadvPY6QaHbnMo4MTdqb
8Ibyx1VuqHB6uLMvAB/sOLkWwlU5gE9c7mPx6V03tKioK6qmEx4jDevkY37fRcSmy1hkya6AgNZd
M3DpgZSSaXX7yf/kgCQroUpJ5eP7dyJCXoLnkb7duHy1EyzpyOQ07SWHdQ6ho+2Pz5QqVuNV+Xb/
+nzX/0o25U6k8C/bGOY1D1HrHYBi00biUxVLIg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5888)
bSPFs3J6xA1v4jww1ffczI5K4pc5hbI0d1abr9AVdkVKJiEm/jZ7GzqHIhsTqfJXA5Ri0BdYjPrr
tibKsYnIxY1jRtMGlv5Awt6dpGDbmb8017soKKvVMlhPcP4nL8ehoi1XVQQlSxjhcS0m9D1cJAvD
rt9vIU4h32U8lZca+2oEOabwNTSoF8aF6VaX5sAsNDvEAl7VISJKGklpy6MeXITWWYyyWmxRM1uj
92Dn1Jb4wQLSBZSSvJmSB0LhyWoAJKfMbRm1WpkbEzgKq3wG83l/i3orK3mdHJ9lKlpNuftagNfH
wRxSJQzZa4MH0ISY6VjKrVM80mBJqLUeBZz/tHndGUbLUs0M6ITTisSDtOEXdKpxXhUnUouFY3k+
SS0NTvUcLFXLNVW11avBVxlmcjtgJNYJFNcLatcWpPA8LydC7lDnPuuiBUPS56ut1Rg/aEgXulRo
gSN8fzmcGDxTAc9AvX2Oy8B9YAFQWFLdHRgTNoYWd9jENrcHY3N3uAkAK5IK9Bcqje42mXuMrHpu
OM6dYLHYIWsfo+XzvckkqdhFrLsispa4yjTmLXq4djAYH8ravG2B+7GONKDFVtG400zaW4pQJiz+
tNdZGKT66bn9zGF4WKePn2RNuEdbb5g302aorr11KFlnfcEVgXTRvL1h1TfqSq26aDPRKz4QAXhX
7NNdTvpjsGHWq/9gMp6es2qNpOPAV7bmVjYyN6POy5fUnYr5t3F5ll6Xu4DsyjIO25W2MWsznvuT
YzdvXeYHQnunua4FFWonMuyL4ZqLFYfYRhQueFBQ0xsXyT6v6G4sq0aHdcrPXR+JqTtij7o8rn3R
6gzrWoJcfHJUKcM1MT6JhT+5XrEyND3iJxCsKkwIt1vbxJHOcvmU5wUmxIxQ5lWtHJPTm89i9pGa
75ME6ImJnJuxwnhmhYTm8rAgwQAK6RNsT32pkHFJMjTfrym4tejsuvYNS8orMuv8VoRNkAok7a9h
wFt5DdqegsIKLZMYqtJwhaJCfyEHhl0PAGGsqxMK526vuYteai4/CcY0saZA4wbdzSR+kcRPJOQX
S6J3O+przo+7+PGf4pcqSoKpK0GS5HUA7mkgPKO5PeWALlVkZQyvEKWUhnBjL2mgkMeLdveRd7F/
8WWNyQgRu1NkRxVGDLMKym5JsqNrB1cYimRDLrW2IqTXnLcr09rF9bSD6fxdlS6dlPpS4BYeQHeh
8x6wQEhjZBIFDGZKjjqqC6GXA1HMG15nfU2TWVN06vLtZUrILh47vFOS9F4bum+nBFJTWqyVMl7q
2Jg3xiRW3jVdVvmjoo/6YLSLpxd/pRCAVOtNq2UXXM5ZvxorEi9KlF4VIgXUHKnHmww89xpjlejb
O7PK0tNr6qi3DwNnBReCuM01WhbnkkVtg8CWNN2S9bLGqooSxZabI5TOeM1jx1RDktwHZqWQaejp
6khMml9/n4/4KeJJhkZb/Qi1ZUELVqFaFOx5bFFjVCZH/M9wnEUsw5bP2NFOyBfTKrVpJuIGb0sK
BQ0JEE9cwMsXQbpl4ecOgkeHOSZOFm2z2QLIPf508Q5Y0De2JqCIpsdA9Sh3/i3DqPanpCerubrC
gkGmt8BpVKuQzOxsLFUkVdKTczV9JW5NycxSqklt92FALquJPoE6VychHD1bpkvr2EWc+4DjWydi
Z6Dxxu5wSqpjKRxsGOK4jqUa2ZQ6WxoOWazJo5uok02F/qn8RqwtvTatzuR8q+34TqwmoHoGC85r
hIuONxkbfQXPqrKXy6U/tdWZJONcizaotqFUr989BTKUyd7ApXk6i7MIhba/tlyWQCVym6sI07cV
eIDbmbs6ne0akVe6p60Y4hDLq/y1UO7AYDiVVx/NnEGTDWSGEy2sXSlK1d9gzyaXsV3Fx1RNNfJr
pG5/5F5qYbGngfO/2CLbcyyeOskvSGjCpqOw6+XzT7Sbjy0XIHm8ht/Hi4SOOGzZFSI/ZEsOM5Du
thOBliYnRoiUanfbLBOkjE8wzcQgwpRPBtW2GnZCVme8QMhII5KWDjs65endmsaKs/jJW10Q3ugB
2252XVNpyAep/tUD5SRV/mBZFY8mYe60P4X1jB0ziam+j83x4d5AvVYeXZm7fhF8fjZBD6e6XYC6
+YXxOUXHgSknLeBTMYHBIgJhF7gn7bif0pmGM+H1Do0ylPDulsNQYDXb69YDK9sJZFfk1NlWBL9b
wYjr+5RZgALvm9HGKGTaACdY0JuFAAlysD5NOF71Pze1fFn2Y53pQb9FmXKAPdjTHftOJv5G+aYU
hPFcgxMvqpyp5zMi1U5CGHZNZTGAPvWh0a51YfburUXsfl8jqqOSf50M2Yy/MNuyr8zWexLR4iLF
Z5joHoBDfzBXlBmSq9ODc9g4RVwb/TchcOp2A2Kn3OEiEqOTcPMdMDd4WuSylzDEV3bgi0whY4Ru
cTdZ9N+HOzxsQw/9n2OwgX2ph+3trd3RZQLIPYIu+Hj3uVZi055FuSc4zL1GGZIyZxrAzaUP5t+I
gocjkVSZGgrzV5hYQYZCwkL5kgxRlRKlOSwtaXVaT6tRspREtHQL+zqz0QCVTsieUo+W3/9KQmAf
c1lVACR0gndAM9DCWzlfcK20sS/ijr0EPNHbh6mb2dceX6K4vjYBNy4GjgpNPzdtbSTW7nPYtVmt
hpnXTVptPenhePlAesAwB0zVrX2EPKQ9+eoNyckE+0V7DncW6OkfTjyfb2XGNpgwFIMqZsDohLBT
e7UeVBrHQhFNdQqZ+0Z4wOnShqw+C1aNjTceR7dSxj/s9QJbd3smrKr2ebu/kaEFWgEE5/IHwq2D
QECmJfCj83yW1y4lxZ7PAgWKGdcPXgxVAvN85xG1hDCkSmJNQNVttmnHRUzAU3c0qC2LfeI0JEm0
xTpgZcFdLtHG1gZvfSIqKorpSa5twe01Ypi5ATTd1fMnTL+ByJ1t5Hpo2ftFYuVbX2j2ObRYEwon
tcCM/eZvl9VkL3gzRUejHh+s3+JiyS5zL+iDKhxSUyfBanV/tT2GzTlokT9vj6oT+9DUB9uuAhsg
yh+lZjwWPQn2Dqvaa1qA2F3QGUJjjoCJVLixLoc+dT5QgVvbtnUvPXuotkFdE8Z24nGCFl3B6F2K
LbOvopxYGUxuo0bHB681W1+h+NppG1venJ8Vn1grK7qnNbHjhK8Abe86JrOsS6F79+yfZRfF7J1n
DPH+w3jJlTmRPZj/MO0zFVPm++6xNJZqFJK81UNu0g6ejKO150dIRug4c6dUSu+j6jITUtwlhlcB
eBUs4Az0bJ28NUqxzyozX8vma1yVUzO0/gFfXPRHp3S1Ji7B47qaQbikOFEglyYpWEJeoeq4dVIg
CXWKBojB5uObEEY4j1SId5XoBMFhPsfJYgkWf+IFrQU7vFuxddw3dF7vHIeTjVkJix51121YvTv8
J6XSYczm2jnG3ylZIo1EdstGuVtSlinSZq4OKOLOIqEidXLw9CmHocidwrPc6H0l+15CYcRID1VX
FYHQYIxaWzinnD+Ff+g5DMXDR3iTKH0WDSDQphXLIF5ljHK3YbKTCHUPtACIIiiLVpx59NctCAFh
Ll/cQWbYAgjgt5JgPaMryJ9+TFvixjvxfSw1LeRpPorbPy5b7AOObaw++r6SxgTzUbC35zUOD27m
+5QbsXbxYW5STTPHN4qpJQCGHaH3606pk4sHlZBBidylbQSe6Tn5OWOAJ6muqDZBhF9RhhL6lyaT
SSFkpc25R1dTnjV73Eg9OVbBORxKz+sAemZqqWCSL45t09TdL3+Kj748ESpHnufGJlAdjoh9oBV1
SImksB4pNDanG7YH4vE9ODBd4nKzIKd2wS2F3vs8AwvDOebMx9bn3iHw7/XnyUqh67OhtYZtdPY6
DEGnST3eSMAvZ8salR8IIiNbVuf5/JdfLeVX+yMjXvpc9QamNOuKAS9/h8Y8KeROaJs1s1vz0ZPl
UuCRRq7lMs+ekLxu1v6PhqvxIhDC4Z6+5Nok0Mf/j974GBQVKuX2BlEaCx7sEe+CM9L00CblZ0Yq
xOAWIv4gElb5IMiMD79tesiS7ymyMwcTpbERyJ3dBhGoL9/wgs+HDt57XODp7XW9e2TvUFuEyZot
/cO6NcMP2pTCB6WIwrSzyAjGZOw9ss3SY5wIUCCQXu75ctYlqWMPdeTIJsO1lgjz7EeE55tyfAIn
NE1qRVtlGaGLHt57XqJz81eU1ct8DkmZJBcR7WrJU5HuZEKum0oI9o0VZ9OcguSFp4fVvXHys89j
4qUmpYP/xyxuoNUab9H8fdu409uJmDqy5BrY3ynH4IPKC+xc6uA8C3p2tjtQskY59c1hIVzYNQ1o
v4txXHaR7auwvl7+ZII4H0HA2DKJP0SMmA6m5WU6l5XaJoI8hAcE3b0aGAnHy2eeuzkZMEs7Pdl1
24mgfOB7m3IzamFqo8yyeRsgkX3ebzfLjZeAPIzNPcXl0zlil95ZFwMlEofKITfYfR+NtyZSj6Js
txyOrXLYC/vMQPlGJJzNf2mzhNZt5VtY3zRt/p4XSVaxBFq+OenU9is+UMxC+uag5zsuQkkFgSQP
RGmbcvexUmDz9VUPqg+ZyBr/6XVQwDp9e/FqQw3Tnz3zgiErvfGlseZIS27fdhVCLohxBn7cBe6p
z0D+fks4jwlV9rNW2Z7Y/LgyY/R80Abh5pkKUmrNIDo9TNB09VCXUcQfxGkgwXq6L9/5kNgKPObe
Jm8vU8nsJhDw7JCnqq1bCST3sK57UPspy/SEVfS/pfZoj7RnZWlVlwUQQD/0YK4pVm5xzq3z2pGk
pb9MD204EbAgdev/c02qwQV1LH6DWydlT4MZac5TU58FSq5N6tibSl4Nf9WYt+y1fmtJhB08tvAT
LeIaxJMX72sRrkz45bKOmI/Ff3q+mgplQb9eEu5pBMz8Vo5HcpKoj4UnOpUVDUuojBEPmrqmwpSt
eU7LRDCTK7rlks9uV+GsDuLnAS8EFYsgsEucMzkmbETWzTUs1AcYVqk/UFLgof3pNPazu6KiPfCv
fkloAlOpR4VP/swYfXZQP9UjK7nIaZ66SbGMvkgi2ry1YL81Kb1ah/GUkwc0j9uDITPcX8RrtIeB
LjkXY0PR54B8GR8GyWSkPyObOvlBMWyWiao82F9Q9v7lmoCvSWvN7ZfNQSFlitq4T+nVjTzZDsQJ
JVqzwQKYGkyYILytBqMUWHBEkTiAZoeVhiqu97fiPfkMro9dpY8teRsBoNd+jWpykH1WE2ilSXqE
O/+ObepcuXKFpxug6yIP9tn7EUC6XPxpx0PJB6c8gmUyMAGjWwLz+lRSVWrFOhGLt8plCnIEkxd7
Hmj372wdzAJnTq466ywDzmYiUsqSkGicCVu46JafDQ/JceWNBvqtfihzFIy+QBNetd5bj1kcQaxU
SI2Vwkqez8+TTvnXlkH9SNj0VpxIXcTZdU9hd6xAGFvzXKmulvYxqV+7Z2aEQvvUQ5Jby4aHC4uN
2fGbqcxHC1jRv3qrgtEIOjS9T38qM7Bc8q+aUuxNsCD76yIY/V8exybrmRaLwpseGEolHpRm4Ubg
w/AkVwwvD//DpoPknTK6L2IlMMqFjpQgBKss9dhnQQ16aAgZNDNOl4q9yT2ReIm5UhNgjzlo/xqe
zKmPf3tIo49ccDav/af6dmwehTNnN3rDVm8nOfs3LdnwKL0WK20tAzkOO6nF45lDI6ZhYAtMCD/g
9xyroW0vxAZ5SXGrv/zA5i8DO9ZiaIAA/xzSQYnL9LFUKoZnr87up9BGQKkYKFGHoNrbJfvboDzK
swDe63Nk1Pqv65u57DkpjcRQisUffuVy9FMWS78AaZSeroGnSeamAo7E9dbwE45KYyCd74rEP/z4
AhmgAN4fidENDfppHM3UFTD5IDA2pldLCFB6j4AZbPuAMFJjtqCEB8ucrSLX9Wb4tct1jHGqfytT
sUjMkPeyMAC0QHEjDfGcIXn3NUC7TGYFXUsemk6FcfcZIQt6vRUUp8M/7JghudE3trTAMTE4OAuU
aKalTswOVSrBPgfIQA7I0dBBja+nz3wQJbuqNETdvKSoYfTGDWslqOw3CD12tW0IFOpyH2n0RrS+
gLEVIHW5zHcoPnubvWGUWfFWpoIruBtdVsG7yCVfOd+TPi5uixONpSdTiujtGNnzuNjS3SuqjKiD
0NMmFHek92x2fAtQZjKWMCe6yn58PEoR0+jeqZOPMxkTGMgGWZNbOJu6Crkz2whkiFbn3bh8i1g3
udGUyOtrmGZui+bDMw9OCTpaIdlr2E/vUywgqjVtdpn3kxZ2VQoAXCq0d425vIJI22vt3bqdGOVz
76Irh+CBfc5r/rLF0Sw/X+ZZTmJaazxRh1KRcUdKuDvVEu/DvPesrr08XK4dWxCm3bWbKPvAlEad
kncSfy3eADrs80WzEtBd+Audsdntxr0wBnVw0JSbTUFQ8i4B6auCXyRJv7Y4/k2C2vCOpnmM2m1K
uqP2rmuQxrM3IxoKFyWrWZqDDUIbXBCtf0pz2xoj/lLpTJ4d8BMy1FXBGZKdk6iUIHU9VMPBeF7M
NjI3c/DXklVz06S7Gc6ksf77TmUAS8pXmeK1XICt6QFHOdMuZc9NE2LIYdTf0uavj5vJlT39sAc9
NDiRus+Znkn3GsmdpZwzNt+G7kWyi5XTwClvCougGf5dXXbIhaZnyWFxoyqitN1Zfq3ZGkGmg4hV
u5B7f0rL9gQFrBgX44rl6JqzLIKAsfQqpOU3kMwOWM+yLyfq/F18gaDV4BL1X437NkllkbAiOsY3
qWiNTGZvrzoNqknSvw9JwDzV2jJvSKRgN79AYoaXTNk55KS/yd08wJaDaXeoWW9FBbSxBSS0scYO
AREDgZbDVYfvHxsmRLtCS3NUJtHdapar6qVwvoOqlehaH/ND8/CP/ef0GW2Q47QnYt7PrmzK4eMU
pKhFgWIph6V29aflOEdnIO4o46hTLaTxsD0eIB2DaEUcjOJUoH9Drx/15YUXHxnh9hcjiW2Ky78T
z9Pfg47y372e64VvhRu7vKHoq34/4DQ5+cW+ZGPdH5X2sEfVRUjO/tqjDCLTMiGtvHS1m8DbOgzw
rnUv3ErS3BJImbrKui+jEajrhj1g5cOKjHhBQEdUNGiSCpjMvVuYsa2MxxQ6ZGJWhVIS6qKcbXXK
5aCLws//A4wQmyEAIE/gzeV/sh/0udoKm2a4fP2yFGpyhEatKNLVCQ/ateuk51DAuFFUftLWZlGc
9qPUy/pNcLVr2eu1GPVTj5TYvUcuXerreKqmwTKhwNSYq/4MK7HvmodqDikDeLhoDvzS1k8V69hW
DVpCcPdF+X2Z+Z18ur3BPz+r7eAmw3keL5/TW0vXbNQg+l0ys1fBTxlB4rtySS7jwfeljURDceRO
UcoqGiaABfFeUSPu658fhoezpaeuA46JWaLhrDFV5W5Yf+oN8ZqkPSfgyJVYmulNLL5micrZc2Bl
eb5wqNNbMKh+x+nOVB5WqfycpHJ0wGP0YIqD7ZZzbfsoUlJKPsxPkpINV+IIr/zs6Nt/XosMiSF2
0zjUYdgpisFq/ISEcvmA4p/O8yTgRirajRmMOcbfTa4pO7JyPQlmTO4y42rbdWi4IlyD7UBtogNJ
YIJ/iwyH8WFrOe8lk4AAbDtm9WlnFCOUJ2GKa5LmHhRB518pEt24XBmeNwWuaO72QyHCr1RL7fLE
jFttzZKjHs2LE9PO2tOkVevOFVL/dOn2E7b3Cw8ZyrfvIOwUtM+LUagQkrsIIzDz42UPnom6sDqU
5ShpPo3IYqrnv/q4xEUkPR8mMHyK1wKO9ALvdtZkKP5vrU3zuPhdWsuXPACbcUkgwnsj3zszYLK7
VEx48B/sGrK/EhNW+U//xDQ=
`pragma protect end_protected
