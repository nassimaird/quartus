��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�y�ϧ�6�F��.��"�Ln)wk�p��5���3�">�@��|�L��?�_�N��:^J,\��[A�TI�?���'G�J�5�e("R�N
ų<r��b�_�b�x��(��f<��!����o��=�_�6$?0zV�p\-w�1�`ܦ�	2y"���]D�4�c1&y`�=�C�����[/�9[���u�� ��,���b��\��J�#\�K9�%��t�!M�� �*ͨ��K7�}G�֞��Z:H�=8�W��_u8ҝF4���GK7s�y��CT����%��z�*�C�oW*�i6�c6f,������ �3h�|�����i&rX����]\�ͤ���m���>�{FJx}��Ԕ�/Ң{�s���q���;r�ҭ+���m�#��r0�Z�T0W�'�9p�P�Pxd[.���2Fð?��D���ݛ-uҾ��_܏��и���Lt}�W��D�y������J7{M�X�^F���U��o��f|����:L ���ejIWz%��˹��I~ɛS
�8bӧG�����#��&]�������]�/��Җ��&��B��Ŗ�Vn�/�F��I���ݫP(M���mҥ���[���Q�L�����v��Ṽ�|�yu��P�r)pZ"Lbw<A���*��w�َ�`�S�!����^�E���ׂ���ï��h\�����vw��$�J	^������qw��|�߁�,�A��f�ts�q�����p^>:.�V�w���&~{
��$��������m&G��><a���I�:A�97�� ���E�Ϫ5������a-*$�|Ƙ﹒Fe��n<��ˉ�����,pW���P��	GC��EX�+�+�'+�x%����>z2�~*.Q�I���ze�C���x�kU���~ӿ�^��8SW��/Z���?H��:g�o���n���QM���	��������o[0u�5�.�^::���χ�����V�T���OK�T�-3�0V{�w�4��s�o�RU'^�����D�Z����#Ň+.�ˆۇ�N���6��$A=�A���D\�O������e�;SH1 3�vZ/�s���_"��t�(B<��|���5d9yu��K������.��X�Z��*��fA�e�ͮZ�a��e`~��+�4�;I��-�H�X�~�7�;XIg�4�M_Or�٫��p�*���?L�P0Dԙ�U�bS�X���Hl�a!μd���'Q�Ƚ���m���F�������qj��O�}�����Z�a����b�##�c�$򐮕=�K��1sS|���Ε��y1&�K���gp���Za�݉�ٟV>�9�x:��������XC{I�w$P�����J��r0�1P8dd"82)~ufc��04�l�Q��9ul���Y���*�~����щ��T\`��Gju��^����k�P��%���3�S%
��TT��y�k�*^�&���b��KQ�BV�nPg���[:����ɫ�	hi�XR�wl�8Dq)}�[�b�4e����\ަ$�,K�6��k��cC2�_��� Z�3��f�xՒ���: �v[�+��mp� ^��l���v4@�y�'��QE��Kl�ӧF*O�w�C��5EO�dLpM���O���٩�^;�-�r�S�G-� ����Fx���hU�h��%�u��R�Fmp˞[u��PHg赊��;(c~�|�� P �<<���T!��ճ��B�<�G��[�,0]����E�PG����]9v������ً+�����ģ��&+�_ԛ�CCC��zmL����������x�2B��k���N�=�Cl�Ɂ	��2ɀI�>ۥV�!M�z���� 7��/�:�zNSb�g�;�:k`ב=�o�q�x���D3���%|Å��>�|FN����,8�������)��2t��g\�E�i�Z59��S�F0ķ$��O\[D�m���/��}�2��D�He�xc�*X9vt���fy){��#-Gfx�4��m�<���6Y>���y�I�����=	*$�
��.`ѕ�,y?E�\�T�;�iLH��>@Z�W�v"y
�!����}��CkJ'mh.�s�Nt�A���O��3����!�LdIB��:&�o�;+���|�����G�z�k��Q���/r]\Ca���Z�^���Bv��+Uު�,l���˚:$���iU%��-E�Љ�Y@?m����>�H/2�K]������eO����݈�x��D[��XM� vK}�״pQ���o �bQ
O��:�)2y�@�ɛ��@(���8t�}j<��Y%4�J�Zc�
���Fd_���	��'�`�X�cM۟hOz@}	�]D���~���͛�0 �a]p#�����Q/����e��UX\��G&j�ch�ac;3�	g�`Q��%L�N��=q��	`�P�!bmFpL	�N�ni����,��UV����}�M�r�<K���#�Z���`Ú��r��O�?��X��r��"F<q�\������h(���u�h�kj����|�91*�ɸ�U^�#
��ĻG}|6��>Y��S��L{ޟ�&yTnU���~K��!�KN�r;��:�9+�u]?�/�Ɂ�����W�('�S�����m"�]��P�ｩ����W/Y}5G,�K��)�ϳ��`E��OV[���H_�� AUsU�W�f{��c�G�Hp3b*xrL��s�.1��+�Ͻ|d��%
��l�T}Gc�
�J^S�\��C[�ǲ�~rc������N�4H��%R54�^�:p����%���b��r����_㜅!����]
�@��W�eK��kY���6_�"w��(��HD-�w��uQ(}1؋�r����7�&�V�g�E��o���E���Z0� �WU���́�f&5��U򧁨�W�;�?����t�'	ժY�0�Γp�}/�khԛ�T�c'��z�>�n�	Jۗh_]�~vڑ�Ė![S���W��AW�˾��g�k���I~�r�;o_$z5��v�,ǆ��g�[q��݌���z�@���jp�D��X%
��}5���H�64�#�>���kӀğ�I���K�}K�uz�x��GK���Ѓ�K
#�|xpG[n��p-xEa?�Qm��#��a}q��7�8�����G�F��PM��r�R�-���i�>���l�
�2_IB,��+	His��\������6�íQ]�FDK�\�Ũ=�a�{�]7t=��{� ��P�!a6��8�ƿ�L��v�B�K�`4��e�)�ӿ�@WDi��)��`F|B���{�5�
b�ɇMV��o3��Gj��pK>�1��8��u�<1�U�b��A[Rʹ��%�j!ٱ�zO�`Z>�[�Yxdn��/=�Z�BO�K$���:�r����FlXŀ�F���k8.�ڤaυ��#��`ஶ
,�˿B��u��A�6���Dv}�"����~��!6ژ��Vj"��D�"f>��#��i�+�zG�WP$u�d��I��5��V5I'���ߎ� ��.���`WG=����w�x�Q�u����f�H���j��h7�f�e�b׏"���P#�&W���\!�o�:cM�=Dg�&x�<.�(Q�Л!��o����X&��|�W�e.�����f8�G�i�1�ʏJ���BY���D����0�-.`�*ܧ�q�Z[��v|\Jr%J���C"�����wur����]B%W�ph��ҁ�Ps��`}��r�H*�Vy��
� ���\����T-2���B����)K�h�!E�����P��1e7�K��r=���vg�5�<�T�/3�H�����"F��X
x��>B�J�(����[�3�BUП9� ��*�.8q:J��I(��9°�t�� ���0�c�D�<��!�����l��T$H��W�26]\�9iu�𖀼[+�]���)З��InϘϥ���'��ΌY`�����ɡ���P��X@o2��~z��oc�?u�3ww �S�ߴ�U������@n�ȳ�	:���m�@H-y�̇�>x��%��g�lV�z�zKI�T���� ������^��n+jŁ�>�v�i��=�����k sJ��X����CjF����oA�>wP��/����4��+��q߃hFc>��e���i�T��JN���6 �M�7��4kp)�(nHl�z�l{���ߏ�m立���>�z��������q�h�U�j�6I������ʊ,���VJ�Ɩ��|�x:]ȣ5��+d���:����f>Z�R��ݝ�R�&=�v����Ƌ2��H�~E�ph���=������§j����K��Zygh�+�j}���u��d2՜w��O,�fMY,�8H���ϝ#̡��f�!*���J��������Xf�u�����O�Z�<�;t\��ݰ��C�C���ѿ`$�PMTd�B5�}H�\��g�a�ϸJ$Ag��A�(#���b�Y��hո�ip�GYT�`��J,1��M�tt�������j>ğ�Mx��C`��8��x�U��qE�#�F!�H��."X�"��B�����D��!GK-yHl=7�@�I�f������c����wF��앴��>7sy@�u��ruBIc�s��yp$��!�+�q,)���9�M!m/	����D�U!�߭a:�*Ԩ@�6���ݧi�C���W��~�i�����3�$�W�j�N��v�D����Vs��)��CR�|0�B{h���$�M��e�W'ҚkU0:TI5��F<��<�� �%0<R	{�%IZ�A��Ci%�o�!=����6[
�\�݋�Q�3���m�h����]P����a�-tǿ�f���6�"���Ѽ)�C"n����{uU�B�>VS�"���"R���¹��!����C���;t�a;_��k`�DS3�����67H�EV]�r�<fy?-wJa�.Զ��~L�ȱ��w�v�5�Z�Ϥ�� ��x��q`0��Nt�Kcl��'����*~��+W5'ͧa$��qe�s��}='B�Y�d'$�X� Ž���(W|z'\����`Fum��b�+�M��|q���!X�n@W�@�r�8>��3��5ˋs�? >�?���x=�Ζ�-�UN��g�o��BXO��X���م�q�k;V�ZI�*IQ�.+���*_#�n�����q��QTQ��>����T�I�΃Uƾ7�/7�ϑʸ�ަ_�vYu*Q!�BvV��E>�2����,��=fٜ���+p��3ӕz�h`�GV[;��&�fr|$��zպ3�diZGQ����sJ����y�'�b��\%���Θ�s��{�=Sdt��hE��.��kۺOP7���Kbب��" D��`R�lYP(��$��I4E�<W�q%dI_��^�<;b���
zU�.��ܨsZ�[�>\�������܆��ET�T�IX/�����z|���;��IMP*d/�}�QD����Jl+n&�aךy)F=%��Y쮻*�O����@a�T��+��}If��I|X�G;���*e+�vծ1P{��y��:7z�X���^�=ȕᏢ�+����P�?
���*�����%�{�w�J�]�B�̵<���^E�wX	V-��ge֦��{I��:��M���o�ͺAA���ۧ$���Ж�g �q�6A��ä���9�o �ORƀZ4�02��u?Z�N�:�ẘ7�ͥ���������0�/�Pu[@�w&�B݂�o�j����s���hqX�]�đP�Z�P��h�j=]
g}�8��H�1�܃7�SQ<��Gu�����a�����_)|H��!�~M��dټ�����qkJ��`�-�!���/=ڿ�#���/61�[y�EQ�4E���h��u�* #�&�@��S���WW��c��H����4Z��$���6�Y�~"]7'�H��؍��z���%��E�O]&��y@�V�c5xq!A]!,����q-�D�Ƴ�M�7յ��E'Yrdԓk���˷���sEϙ����6�S�:Ե�툲�䰻L�j3�d���0s�:��g@<�i� ��Y��tdo蒓u�q|�-��_x���A�]
CNË�o��5�a6]8*��5e� ;��*Y�C@��ΧO���!_f�c���-ub�����ڼ��MZ�4�H?o)�%�T���i����u"��A����+Νsz��xX�5��P��-\Q-�3�<���xމ�.�7]�(�x2��W�����j�#?<6�f��!�V�W<55w�`z%S<R�Yw����u��p��AY�����	ٴI�Z!b��+{����5�"5gMG)G|Pk�o�(�4����"����#�F�u>?�r�p����>26�X�M��C���;ߙ^�ݙ�$���_��v�>'7-YdbH]�1ڊj�=ޚ��B��:��O_	٘pFE0�`>���6������a8���[�	��p�J��O�aF3H����;�0\[@%�}���f�~��IQ��#�1���V���_���+�`��8<��V�%���c�ߢֿ��6P�˷��j
}���+�L
l�%ǖ��3%�ʧNĮ�d\v9e�[��;�4�X�Z�\�/ǝ�P���>I~�/m
Z�a��#���˔m#R���Bc*4��G�x�ɠ�O (\rߘtc���!��R3�n(>�����	k
-�z,��)��ũ��r�~�Ei����ǽ����؀��wd��0���M���3�,�qg�(#�D�T�ꩈ�X�{	f����?���8�	��f:l)l�U��lڧrd������N>�2��M�o����k�ͫ�Y��Z������We+�$�����2�k17�x4���@���#�}�s����.�yQ�j�z]m�sp��gc�@I`BQ@�n�w*�Y�L�&�9"�.�!��C*��K��	R�J��m�QL]O�]�wq�����N����#�|�Yۀ֪U+u�4�e}�J
m}��'0x[P_�`c��d\"�(![�[�������ST�˸�f;�����u7���K�Ff��ۭ����69ƴɐq	vy�I�G)R+��K���ޞ�hJ���>z�fUD�KZ�j%���&	9��L`_���*�A��4����&l&��)St`*��q�<�2w�gR�Ҳ���y*&�Df���� \(�䲻Ѩ�p�*�kr�I����x�D� ��1�ң\8z&����!q��O�(/-��������k��X��9N��)h�Y$�����\�2�@ď\�޹�{�b������o���SL��|�K!�֮�db
�M�;s���'�)��V��3�-zFA𰌁fq�8&#t�\H�o�`��1ܿA_Oy��y����zsJ�S�$YM�+���?m'���6J%��u8I'�ʔW��N�Z���H���t=�fgQk��g�nǘ�?iS֒d�&��DYb��%z�S;�W
�ӝ!FX�'c���U�4�H1�rv8+
[v�㞠u��=<�@�'���0syL��N\�#�"6�IV8���E4��k��2c(D8�C��ȅz-c*�k���-�;F���2�O�~��7 ZL�7A�%�p�� �՗��"�A�$2�BU=%5Z_��!�EH��ݤm;�܅NYS�3�c �v@dE�ixX�~݃��}O%�9�.���|����lXuR��������$[��s�z���4J�F3��h4I')<Y�E>�'�����bE��������DRAi>��BqŽL	�����;��I���)D�{���� '��S��uK�p�
{|	�Oz��RƤ��/R���k�ֽ>=k�25��ܺ�}\sƍVx�RF���'cgށ0����L�YkpR�u\K�Nz�TѮ���7��?�Y�%��	20�xB��?��Ho3���%N�*_WzM����ιe�$�u����ا��=��pe�>1�!��y0X��ZX�-�+Y��r�Vk]AS������램'H����g��Q��+z���
�J��R_���+�g9�����Z�Z��<����r����M%�vJ�P�tw6ضqCv���a �\lM@swuH;h�Ecq/�
oBR-�6	{|إ&\E"�;M���j�K�t�梞�~�F�J9Q�eW�q�;\LFN�a�Ò($����x��3�	Y�)������v&vP4NE^�N�0���Z���\��rV5$��H1%)䘇��'X�����C�����W���(��.�A��n��\`i�Q\h�۱_�X�?V#Dq�/S�\�����=q�7|����>03��cg_�-$j�~��b	�Ef��7}zUVk��@S�X�h��(IO�:�Ѥ#�E#g�od�>~Y��x���a���Je��x��?/�@x�+��߂wJ�׽�:�4��6l�D^T���G����Q���b��kQ&r^�J|�\�|r/N�v�+���H�T�ͽn�50���G6�L�s0�~���,���e!�]�ٍ-�F����h��#�u`�U�W��� �0�I�L:�q�G��v��COa�Ѱc�r֛�0�V����J{�8�/� �Zd�u�¯��F9٠��Wg�0 ��ܕ�A�-��z��x�΅��Q���Hޕ������T���o0�
Y3s"Ì�j��*? }=1Ρ�tw�j��\z'{�Sy�ć2Z��>n�ʉWֱR��ɪ�S+���)��x�ں�27��`�:�hp4"r"U��>�,�-� �*q�j!Miyhe�����Ԣ�BȈ%�{���-Ǚ��}�a��'�dmU-Y
O�va�}�Z;e�]�I�9�Xz_���e�m�y����:���	�jѸ��!uc����\ʹQ�_�ˍ��v��H �$/�ϊ�B�ފ��+�璹�(��O��zARɞ�_.;R�`��,��I�K���ԫ�oj��'�N���{~c��ŠL�����=`���1��,q��.���A��I�{(f ���Nbu6����}J=N��	d�|]
�����By�M}�Ǝ��m�QJ=�&z;T���;����B܎jb5���WA���fa$Q�w�q�EC�1M�AbG�%{l5����F�N���u���4��"a&WLA��>#�^�7F���a3w�|8dG�¹I���[�֊��+�!�����1���2n�C��t��p���v�d��c�MH/Ix�e������=��Ufi��~N���������إ4���G�Inx#D��=�7���C�g�J����rIrMlH��P��U�6^�R�.��#Z�#4����:nm>���Ⱥ���a��y�]����3Sf��A������q�m]4@#��%�<,죆�RH|��K��Έ�;0��.��1Q�v���j�|�z`V��vL�=��e���l�����F5Si0��N��Ǹ��@��~��#�({"�A?��n`�K�P��fTr�.�暶n7�,k�b�C�ǆ	k�z<�P��m긲pTJ[F;)3I�F��觵l�&�{�u��mu;��g&~ ��	Q}x�����dǷ�j��f��φ )9����
��tP�kA�[�J�r]��%�I�qٹɜ��m����yg����U\2\����e�-��ٽ'BxU
<�Z��[�L�B4D�Q��1�*��]�!�"�KVE{u�ˠ��B���\aV��U"u�If�� N�)d�m��Tc�_��\��᧛��fԠZ�F����+{x�C"s>d�5�+�E���� ����M�7U6>�0��`����+tJ+� ��dw�H?!n��r���0�%�)T�z��[���Y����G�u�`)��ۨv�-�.[4QbC��>�all�{�����k���sce��!l�$P����l����i����lf7�%{����!�]n���D�\�Z�㱁�^̋؛2bl?�߳öYO$ȯ���bTAu�z˫T��)!���Ee�͏h?���=jX��Z;��ə;p�/9߉0�2�8�	��a 6���4��� (y�)�]\�_�I�a<��H�E�5B<���ug!�~/���Yֳt�������5#_h`Z'-
��Sj,l넲Ղ�Z�Y�Da(״hH;��$�#M^�����ΘB�����`q� ����޽���$�J
Nڂ\A��I�cIfk��	]٬�,��)����l�D���5(:���D����[ot�����?�F��܀j��3�dK`9���Z ��/��;��H		(P3�	4�&UP7�+J� ���_?wt�WZ�Lj\4��yY���.ěC��Y-�??5y�{�m3Uܩ~u\2Fi.<SD�j��<������X13�&�OIW��G~�+s�Ք�^�.̫CI_أ�3 &Q�H��$�EϺSjfF�Ѫ�K�?�aB�q��2���}i��)Z=-"��r0�_���$'ߜa=�S�8PW|��Q�n�)�Ue��e�ќ"�U�6�i�^a�o�"�?�� )��=P!���������:��r�H6�m.���Ѫ�2����L�hXu��Xt��O�_�����U,LݦB�w��${�'�_AKCK7>�@�V���_��=�A�7�!�I�y�)u�]�}�p�[�������T��k���r8�f.db�P���Ř��H�.����Veu�����٣r(�Wn�п,.9RX
���,��x+�93�v���h)�������� s�?����T1sV�$���W�6�*jߟ�D�6']�����ٔ�ɼZ��6F���:�yÉ*���A���{�K@�*��N�B�h^.�Ti���͓a��
>��t3�;AQ��N�-՗��~e(Y�e)��ѓyV�����.6
����atCq@՗����Ht4+jp)�/�����I����r1�.�|l�2M�b������d-9Rg<,�ws.�t�&��INp�:��=7���[b�t��D&f� ��}O��>�k�<�
9�.T���c揄0֨�F�PQ�����5Rʄ��)�VG�I��F[� �4+�C/B>����ZZ?�Cr���+ #Ϛ;�\�B7`(���.t�I�O�)ѝ�Ҕ��@�nj\��;D:���m�����𹍃�z�V�*�j�_��$p�u�A����wE!M�{��[$�H�5��?P͡}N����t&�{"���3>��5�H����;�%Dr��4C݊�j�65�h��ܮ[�Q��~	�$"y
ƿ�熢d�.GtV'�I=�@���)a��b�.����%��J�V�4�:�R�#����[��T���jY��m�.�o�{B�Q��VF>ꯃ��+h��,��D�l8��E����!`*o^B7��B^!�;�]>a�m����0�p���Umմ���UlJ�[�K��{2�g��J�b��53���r!�_�2JB����p�?=���Mf�&M7� �fF��ϴ�t��.�Y@�����!W��S\��*t�)�E�������WJ'N��lqE�ZV�s�d����2�˽�ȸ���в�  ?`��)�,iZ�]����!w��Z�����r-�1O)�����ԭ.��p�c]B�ד��������0;�����z�؛8�^��?��K�j�"��6�{�g�ĵ0�m^���W�{�)�X�$���Q�}�N��"E�bQ(��\�S�{�[�hǷ�E��V���}e�I��1`8��.Mt��R<��c�b�w�$�?�5�Nq蜏9
,����NX��ץ���oX�3B��ʛ��<6r����`n�8�;\rH�)}��ӯG��LD�}.f,=@����rQ0���A��k�N"g��7����H�G)V�&�걉6Fڌ6����'���$�%҆��="
��O�/��:	��ڸi�?���UalA%��l�a!�)����?y��,1h"@�u��$��?�3`o=�5�}�� �j�S�vnF��`&(��&
r�LVD�R�N��z�/���?pS�G@����z+=2�9�!>��Y�2Wv"B��B嵈���?	@��S��f��<�m�; �J���\�6%!A�3N{/����� ���s�t�%86C���Ψ쭠1�K�m2t�i2U���)YzClt�D/hw^(R�Pk��w��:���<5�J��c����W��v�̲Mh&Ɔg�/�CES�r�Q�^T�V+�bQ�P���Z5�c���@��7l�(JW��/��{��;`_?�rQLnz@�E��3�0��g��}F��sR���y���I�/_(��J�A	2V�Aؿ�sO@d�I�R�V�����	�/\�8�p#��ڣ�+�z���)Ú@j骍�-�O�>&�Ѱ_����MŴ��v��V!%�!;zZ����&��d�YpDNQ���$�3�^��?��ՐX�%�uW�\D2�Vmƺ�h�4R>�_0N1A�� ��f�P�� �A�%VqW��gZ�C��l�5�J%��=��$���%p�r02r��(��G��d�W�/Ӵ�\�,P_��Z����H'��&���IB�r7BX��dͦj���W����F�E��U+�k�5��Jh�Kl2�R���Nv(�B\�ɋs�7V0ng�����%�-�P����G��sG�w���,��KmL��*���!���p#��o��c�wq�|z�AB��3�gr�n����c�o���P��17�)������8�J�b�xd����kk��D/�xʄZ
���;=<�^��=�|�L�ds�6�X��u��v`�ȼ��� /�`N�|F�gLH^�N~�sG��~�����T�#s�Hh��"���S��Pw�&[�n?@����[�X�9·��7������O�d˩;�[% m�m���M�-*Yr�5�t6��>p�[=��oV!��gU\:�HY�����s9���ß�_���%�#��"ӌ�x#B�ڰ	�SJ*G����h�/�ypG>��0��!�N[$��T51�O����ٓ�Ї<�+>���W��4��P!��� ���U�z�r�ʦ@���fA_�Mg����p�?P�� S:�=4_x��&FY�_(�::��n\��$+��N�L��:8:_B�s	.��cqv�/��i/y�����n;(
��Lw�>�C9��(�o�{Ԉ�0yE坻4}��OkR�(7RDS ��L�/X�f�18�	�+z�v��Ɖa7�%*�/ٹRb����k{���E�g�zq�54	����n��ԭD�Nw�%���E={}r?J@�q���O�>��|�������'�5T�R�3�e��9Bh���a���e�җ�:�����k:�j�\ލ�-xv�s�@�j�2�D��-���!A����O�c�\lQU2�IRg���Ϭ�bz�FI�	��Q'g���%O\��ڒxVw����Ĕf�Q�,�*�����͸:��'>p�e�
Z����e��߯�m\��h��c��)k�E����g����h}���ۡ��ƽy��Be�D�7���qo΄���g��,��o�GD'g �dC����q�T�o���'D�������Tl������\��%��T?t����/���蝀�,�� ���ҽ�����PV>hH���S��qU�k�i�1N���+����.�J��u^��!Э���MXU}fg%������Y o'� ��1����Qk��߷���QfW�}f�Sw`}U~R5�j$�=ǭ�֛�M�5��J�Q�fÍbx����p#Sa�,֮��Rƣv�k���/C��<:���S��:��]v��lb4��S�֖����!�r'�AZaW]���ޥ52H�"��{���"\�W�=�y�!٤>G�ֵZǧUS���e�w�[F�y!��$_/ ��9Θ���F=�#橪G�2I"�`�H���C�w6���y@��f1�	�!_���>(��A�,Tl5�i	M� R��#�0��U{1�q�o��9��3ޖ���L&� ȟ��Bd�a���ݶ	B�S�Rf�j�D�P��1uhSWbݑa��v��
74�k�yY�ߙ�ڳ����li�a�j/eF�E�k�{˕?�1�.rW�[̛��:8(����0�H�֕�qq�Р|�露G�����ٿ^e4���>h��Sϖ�(Y�
[�82�A��MJ�!�~��N�ϫ��.��6�x��[\Ζ����K��J!ƻw�SeJ�M)��V��~
��0
 @ĉ�Y���:�w[�$蘛�@��*L$��W����8�����b�Or�����o	�3F�bo��;@��A�u�p�[���tV�S���<�
�ņ	�]&
]���BXȎp��7���n�uG�U۶�s}�q�X��-��е��0�O��i(@rp!ˬq�Np�t�
Qg:Ū+�8Pkof���/��o�E�4H���̫fI�2@�z���]���@�<�q$�p����=,�|{�*����������UI��ª��*f�e����d4��{���D,���~>zg��]�	~��(r��<
j,�&���}c��9�I����e�}�Z��T��km�̶J�;#��ߝ�!��,o�EL�tNg�	,�՗��m�J�>H�;�x��jy�.s�{P��5h]��Q��z�A;@SڰY���K���jb����:����b�D	7SR�M�A�p�ɼ���g��¿�Z
��V�O&͑�}�Q�����)��"�#m�|_sxo�����:ex0�^+�z3���O1�&U�-��>w�v�9�&.��kb���jYÇ��G�[�1C"���78l���R�W�0�e�6״��|�߳2Q@QI��s 2	. 0�������5q��G�33C�Ҁ�0V�hD�������=�@<O�s�6n�l/��*�Xߥ�(-4bȫg��B:�Q�6����~�OWR�y,ߦ=�=���)�ܪ1N;TK���_ڬ�[s�qj�&���E��r�>�
���mA�V\M�X�����R%w���rK#��س���g��>L�Y��/'QtJy���c�"��o�H��B>��y�k������ɯ_���"�'�N�	t�.?� �
CGGg���f�ϓ1�õ�l��ظ$�*��x���~O" ��ө]��sbfUo����sQ��Q���Ԟ��R�/�Zo�V�e�Y5QU$���,5 ��K�45��,&�^q�5Y�-?�Q��OŬx{5AŴ�����MA�?:"oA��xSz��Qh9Yě�+^�󔓙����,<]����W��9$�I(�﯂P� �Į��"C�[t�&G`�Cy*��^�BEc�r�~#��o'��T�d��$'�af���2���w����hاǆ��D�i���|�������ĂLͼΔ��3�5-��Q�!<�Tz��!i���O�*�Sr��fc��=
H������V�e���GLB���B� "�AЍ<I�.T���d�kHIqD���y�ys�A��u# ��	�m
3�d��<�H�O���>��W��^�;�?��¶Ҏ@�}[�PG��b�ص���n���0!/|d$i��}?�n�_�@�m���$�-��3\"��$,O2ɎF�v@"�X�VY~NCpB-��k�J�����?���V��x�}�[šV_b�>Lפ@�1�����G	1W��4� ,W�J_��F�T������8��@Mϯ'l!=��Pp˕[[IM,���m�)L,���5�x@Tw��2�a�L�9�tDy��3��{��*>���"i��$��%��KR�5�\7'�g @�qĴ4'�JӻϜ�o�!O�����0��"u�Swi��Zr���B��pi��o��}0]�n<Ur8���tS�h�F?{�j�if�o�pe��DX��dJ7`�����
__�u�d�KR�fΩ��.��;:��m6FY42h�E�cg���۩�|����r3T�����ga���K���>e���ǎ���H�	������س�Ě	��]rlB�.�����s^��N=���zg�[�Sn�,����U��<�2_�Ё+'nOw��X��g ed��oy�4x��6�s�����.�0���;*�,��pv,�T�FO���bg:%�OʣIDT��R�`<s0ďl�#gl͊,D�EңB�$Rk�/X=���:5���-�O�R�T�p��ǰ�)P�u�k�c%H +�����}�uMz��Bp��'�Q�J��gr{����f|R�O��n��m+��6��I�����R�b�qQm�H�B����W�g�s�3����������O `��P�[-g�J2�i��UE~ї����;�K�x�6��R���6-��f��݃����7ؠ��-�6$Z ���cѣ;]2�������2n��(5������~�g),�3fqp�u�(�/J��?GU6��+����o��\pZK��;��u���*~�;a�|��(Q�
"�ar]?gҜ�I?O��g*4�i�x�)W��{�iN�a7���]5�p�i�G�����T~;^�GCg��ۅ
S@ï٬]�Ā�������k�W7���T?'sY	�����Y���\�=չ��������K0gXl�E1$X��;�\�Gݧg�0��xQ���^	�֖������hЅ��i�i6	��f6I�`-�W��`����n���ל&W�#=�rKׁ������d���6C� O��=x�la���ٮ*NM����7��_�b��P17�d53P��&�����-)zTJ�WE���;���v�Ӑ�)�S:���R�W�ܕ�"أp�z���u#{�b��<�]����"��k��X���rd���Z��)eu�-�ڮ뒚yM����?��<���q17}l��- �B�TX�E/w���rj������z�ZEm)̿c0����=����7�uA*�Wa�2��˂�����og��G�̆ Qs*,��vh��X�^?����[Ȳ_�Q�N�qZN�
!�τMv�` ��t5L�/���=[,߈���.�{���M��$�T������8���~jּ��e�C�$�u���'[}�!��%U�t��I�}7�Ly��a�s�{�&<Z��� �C����0�f$�`T�ֈ��򍉣Z�e��?��%}S��.a��H�K���H���{a�}M�)6v!n���9	�r�,�����My|������b���>�I���� b�VS�sYR�6ce''��'��~S���XV�O(��
�v�i����Ś�r��ڏ��։���F�t�hh�l[�=�d{S`9��0|B�����7$�1����G`��e�'�
䮇Fsƕ�!��(�b�M�<oO����'�'&�̂{K/���⇞���������5���	J��5��Ʀۀ�X�eGψYW�^L%��`�ƃ ���=|����Y��q���Y��N`3�q��3a�rξ:��~b��"�kfZ� Tc�|P6yƩ�q@V�W5T�����67��,M8XB���UVC_z&UG��re@����tW�L�fюo�ӊ�J�j=Q����2�3�4��B�����U���w��Uf4~�I��F�<O��V�R���o�/�]A?�W 	�9����y]��k�A֐h�4~��rj��5�c�b�P���T�y�w��9�j���k�t��7�۸�Q��e,�ܟ��(7fag�4|�	,=ڤj,�,ڡ�|�)�����õZ�/f���1 1
�R~0�Tx6��&>���r�3�@�X��@Ȓ ���Q�(�5 �43D��X�6.��l�i��v�`�T����J�
��+�_��q���T��ۇ~�Ǿ[mt6Ɩo��O�φ�P��{��?���~�����"ɡ��.w6	��n�~��ꖛ��#��VN/¡�'^$/9��W��;E�v�OETc�����뉧��8D�d����P�[(�M+u�)ك��)�K��c.��C;���"�RRi�x!M��j� 4��,�L��XYJ����e�.�6D��������@��l�;gp�h�R�1ն����rtI	!�)+(Kd�=��L�?�8��L�Y6w��-x3��5�N����e|(뤏�3���	3ǰD����?����6IH�Su9&=L��j��usV�U� *�T�Ȑ���$�? +���[[���a��|�P�&s�v�u
?Dmp*q�rr$f�/ևf�`;SM��KDG�6d?[e1�.�1���z��1P��_�{:Vy2�޿�(�j�nu20;�c�:HS�I��%���^A5��.QD5q�d��5@�,hxo�B-��X��?�N�*a�P�.�m�5`5�:��)���$����PQ����,� /\��K�0`0��sG���-��7]����e���>�H��(}��h�w�)��NidEc����f��,���[$���[���g4�eϤ�� s��m���va'cYr����`)]vS�Z�t4cٽ��?p��ȧ��2>x&Bh�c�U��>`/�/�<�F��k�X������J���pS՛	���>���^�؁0X4�"~��*�t�8W��e1�H��VZR�A��!۪c~�n����
��6�*:E�7�M	��1}��2�YV+��-� �f���i����
�)�����א�
�����s��ܹ�Zid��M�YO���ߙ�q���e����?�Ghز͎9��X-?@u!�(��X2T�B��*�3�H�zDp$B���^�#��J��7Hj�e�& ��z�Y�,�b�c��]~�;n�?l�P��,M]l��~E��f��m��6��2��qI�挛<��ɿ}����it9�#Y%,���~h���I%�z�Ҏc[J��f��`r�V��v6�MLPZ�߬�kƭ��0*��BHz8v�y���5	!��J���a@H�S/�"Hu+�QR���n�Ǆ�n�zw�q#Nu;�e���=�3'o8���m��JH�V'iF ��y����?��ό�0�T�� ���s��TUaٯ��(���_�������GH��!�=��s�0����͹'"�
�t���M��I��;7��F#<r���(��l�iff$��GhO�e��~YrD�촶@<�>����j�T��`�ލZ}��e&�W�����������dɤwM�b�49F��3G�8����߂(���q��T��aLxg�]���V�Dj���ˑ�L��Ո^U�6>�Z��bl�)����x3`��m��9oy9�bkC���40��B���q/�$�O]-�>β~ ��H��]�v����ZV"�j3�3�T�r��v��f P+,�H��VE��)��/u�_A/�ߍ�^:��/]}H�L��4R����/'(U
�ϯ �1rh���BI|� �Y8-�Y�#�&��*-�t�����`rR��	ت�]��uC"#�/����ݨfA����j6F)l�4K܁����*E��@�E B���r���b�<����9��R^�	���DǱ�������b	m���y��a�jt	����o�:�P����R�gN�Yrl��~Z�D��j�<����C=�$8h��#�|���^��j�g������<��_�ۉ��0�A���M,K��	7~�������,�%d�L��lh<<�0}f���*�����{y����u�'Ec��q):9dȕ�����@��7�»NOZ���#�{�D`5ӯ����b}�抌P%G���ď�T��ف�Γ'g�`����
)E������W8��.��ni�fc�U�ȤĞ@����M���zM�'~���͇��g�#IGxE�~X���T[3�Xfj��8�V�6Ld�IF(6��Yf}��T<��4��4�>��.Gg4PXx�+@'tC�d���N�39���
]�9�d�Z&�SQ��+:v)ٷn��0��{����<Չ_���^�߾�O��깦�OF1��ĳ�����䙎��k`��0�"t����F��P D�B����f�a|��nc,+F'���j�vl: H�c��!�]i��~��سq�\��&�V2A�S�%��`:#3ޖ�e#BḌ���v�_������i�8֍q��*Xk>�1k��DLU�!jen�A����&9�ym�vƽ&�cl���.S�$���௜���9a���bc�� h��GP�BE��N\~9p���p5g�֊�݋.q:�����$�\����D�� �XոǬ\�E�-�C���Ԟ���[����o�6G����yo�]\5��U:�)�W�A��3��I�b���K%#Y�O���6��ĪQľ0�x_dN�ͤ�T��
 �] ��Ϊ���{|�l�bɮ��>֪f"��-jK~֟G�Q��3O}��UB�n����6Oa�hj��3�p�@6��b�t��^'Y��=lO��,����jG�}�n���}g�� ԉ<��y�I�:42.Z(��A��7@���:lK�|�%�IV�$ Y���wB@��F궣]�"�'ܘ�M��Bq;�#`�������Y�U����m?�e��'�ؑg�ڄ :qv�{��8��&���ҪBPƣϧ+t0��o[���$�����\�"�M��ϐ�3��6��C�4�B\�kǘ9�R��Sp����y��i����»e7�^�~�y����j���I���w�z�����n��Zd��
�.�`�=QS_��a����z袁�=�<mXP1`�~�K�{Q�Q����A����R��)UB��V�Ж?P-�f|�X
 M��F3ଇ<�'2N�O���#�� �b"�fn�{�JA�rL�)ޞ��8H�xɬ���PEO�<�X�Y4aԚ�;�Y��xJ�ϑ#�J�s�Z�*Q#X.�
�"�s,�?�_b2�7֒t^'N�Z{`m�g)H1�+�jz}n���|����6��K:5���#������45dW�!P�驷5�#1��V���B2����,n%��#����7K�-8}u�8�E�g�us kF�$���S�N*��I�q���)�� ɜ�{��o}�1惾M{�AV���"�����r��҉�ߣ�\T��&Z����R�qhN1�3�2���}q��Ъ��7�)�ye!��#D�B�j|ڞ�-)l356�U{��;&����fhD�8.:��#�����?Y��B$���J�٭^дzܳ�w��oj�Z����ݪ�0?Z���G�\Jj�	��J4/�;G;1���
���/Ej�c�.25r���M9�=Ԗ������:ώ�j���&�FBՂ���Lu�I 鏂QE��%��������L�@T ɸ ��pm�kg�_���0�Z���ߺ������e"�O|�K/Z�P�#@3� �-��7,<��Bm�&@��N��S�si�;=7S],QH�I�X̥�I���Y�|ߩ��TtO����i6+�����Zx�����B���_2�u��R-:�s[���7��M�|��/$ڦ�#Ёk%�`�oJ��	�ZJk���H�#�b��/ZQ��#�Ȝٗ{����S�r�����b�Gu}OCm5���G,��%�j	���
��Řʻ�ƺ�%���٩dI~�ܘ3y�������h?��>�N���u�^a�=�ݪ�e�ب�ҶZ��p ]�]���@5�� [T��	����G-G;x��R���?BӲ��#��AT���dy������ ����G���E���
����f�K�hIZʖ�O�a� )����1XEY4g�m�ҵ̯J���׷y���^S��uO��jr*:�~5㰪w���a�&�<D�Ƚb�j)&QŇҖ�{y+���e[���ZI�X�H��>c(��h�=��PT�5y��T�� �z�{�Z3��K�6N����޽��4P�A�p�I󄲳�@!h��p�����$s��T	Y��� �=��C��B-k�`k���p�ї_��������TO�������:'	\�`\�U|Wx$���$�soN����nA��GF�6 촛��R˜���y��ۡYޣ���I���`k%V�&<.*�#�ō�g�Ғ$��4%s��6�joQ��c^-sC�hñ3�s	V|� �j�{�Z��,�+.Fl��>	������� ��^�Y^����Me�ȃ������'�*{�J�b����hPU�����}G	����:h|C���RrW��?���H1��f��f������7e%�[*P���c��P����9�u	�ُ02�!��t¨�<RݫAP�)g�H�6nr!v۩'����OB�$fM���pXʙ`q{`~)ِ�wQ�pʵ�Dv�u4
�B\o]�v��;���\����~	��7���u U5x�`�x��U�H�[J�&��J!V�M�=�_�r������,�^�`����Ϻ~�*!��\d����WY:���"Q%� ����,�����񫡩}�R�A�g*�#�|v`;��.S��Ϲ�f��I�P��FN��;9-���M�vz�u�\C��T�
k��b�aO\A���>M��vE�%�:?�RD_��|�D��2��䡆ã�BE�<�ǐm��Z����e�_��I}<�VK�^K�,j�-�����|*[��B�g������K�7kw�|Z)oi�X��W��sqR��^/JD�qm3�=�.%޳6��S�l��ْ�=1�����Z��	��"�*�&�*�nYXP�}b�Ƕ��.��JDe��*�y��5?	���xP��aL���3���܇��DC���6k(|���%��D���TA:�w�@g�nzdxpYF�jW�v,�%�@n߱Ɩ���Oj�|t�?0j�����5j#��F}_$ܖ�Y�E2�JN��:����	���aG�:���Sg�� 5�Z�]sh��C:K������M����$��Z�~���D��}a)@�-
ŝ�\����ִ$ղ�
@�'5yF�$��I������@��+`�!�|���:F��݃�tyH�,�Φj�V�I�4_�.%�!'XI����[��k��@�0Ff	S�N�-���hBZ����%J֜�|�j>V#�I���'e��[�����s�T�L�:�s��Ր>",؆�},�Ќi����D�gqJ���;�["^��x���M���{�� >�����e��{��yh��_�3ER\Ɓ?珧{�wǣr��T��gK�h��V��Y?\�G $�%�6Ty�3?;+�>����ԓ�*�����e
�^�p��Wpa��pO�=��Į�#Ly�����jq���$Y��3�]V3�	e�^��c0��4���@���e�E�7"	W6��G���)�f�~x�=ϞA����~�p���.g�cn���ة�G�K��Pv�g��sg��W��i�B���}"�I�y�d6"�x#R^�@. ^�`JP␹y��X�ԲQ�ꚑ�D)�Э����熫�(��:�ާ�/�ԥ���VT�Ƀi}y|�՝�7��"N,�+�2K�t�n�`Nw�!�Vj ��!�#��4�hB�4y`�m��k4��T�(UC��F<��`����r�U�?V��0Ï���!qKvR�'��U�E$=U��J%��5$^�*���j����Q��Qb+����d��"�2ɨ��m=�Z	(�I]��T�M/�xߎ���x31$�P��!�7F�D�>̢h�]��%}�|����n��+	�h{k������5�O��ɎT��Wsx0�ش.�W��DF�=�i/>�[�M�����a��qf��d��&տ�f�vQ�j�'�m�W�)FQ������o��\G�T��ɔ$�R��n�c�bzV�!Ԋ��C���_3�w/u����qㄈI\�[+�>�D?	��u������)�	7��=b&7����.���3��A���l�/�^{� p�.'Xո㜀]~�e���-�W�S�Ge2���!RG�<I;c�9������	TGw�	hQ~�9� c甶����hXQG�k&��h��څ���xQ����U�%�c�k��^F�������W�e���S���K��({cSQ+��08	t/��R�zF��~��B:aD�m�ˢ�p=��S�h�kR�a��-�){#�ݺ��m����B�,1�PT��&�W�f�!soYb3"	E�c���K�3�_w���"��CO�5��j��|
�̙�~��Y��z}�oxT�mY�Uk�hU�3�Q�{?���"�3V�� <��L�ɅHW\�^Vk̖8ph�?����6c����%�hЖ�u�6O{��$&*?{��ĺ#x��	mAx���҈X|�LC�ǉ�=zH��m�?G��ͻe�K7�_�V.�*djbI�ʓ-�����A�c#x	�:E��`T��O�p��O�u�j�@лW��Irg���n����!e�N_/Sm���\�B���#u�jtE�.@:{��!Z ��PK!1�w�(:ۀZ�r"G����V������2Հ2=��:�;���%�|�5,����v�h� �����n��:ҙ��4�v�i�e�֞R$���&<F�şV�}��i�E��V��\�_9�B�-�dX��C���8�0�rȓi�v�9����Y=�o��\K��0'����z$��aĆ��� 13w1!����$9_ӌy�F�7ء���[`���*���y�ܶ�RU̸�`��5��c�Qf�cΨw(��:}�B���?y���ny��2����gg���G�Ф��_�6��q^ ������k��uZ�V3N�"W�	G��E`�����P���� M�4���^'����6��ʵ��A:ۯZ��C0���>νn_~�(��)�d'��]����`Rx���6�6U��z��-q���)<�6=T���+	B�P|5�L��/evJC�;5�=�'t}�*i<V�.��DZ����[���$˵�2_d�'�Z�-?w��U)���a���L�J����F_٧m������G�
��D@{������Hծ����L�F��4*�@Z+�;�C�o�AV�~k�7� ���u�a]WH�9꾫Z��t2�w��#_�uT�0#�E1�a�2�%Z���|��L�|����C��������e�4�W0�FB�*�#�㭝�;�|-5���ȆH���@�ⱀ�}��;v�?љӵ�H� &�W+��(���:�Ñ��P'ߢ���5���썤m��_�ݮ���P+��u����eiVL�#�u�y�x�Z�ޯ ����H�-�D{�5.fA�$�Nh�d0��">@3TO0/D�\g�A�
G�8�Pt�������}���Δ��?)�������V�)[��F�1�H���̏m"АNΟ �ZV��<�{�RW%T{z��D'݁�}�%�F�.��3����Q�H�:�I>mU��M���/'����R�|:�mֺS�?��E�tDU�u�u�-�>����F�� I��DX;��R�
�fTAvN\�
 ��Sd�Y5���o�U�v�X,9�WA�Z�O�� 
`��ʱV%�!j��'}�����G�B�*�Hj�~
��/�N�I�ZB`��ODqj�F֯k�Ds�V�j(,L\ٓB��׆�(�Ɓ^�>���y��SBs���wNq5����bs�Swe^���q7F��E>�����*����
���vʒ����!3�V"�W�G9�\�	����p{Da|瑱5��[�ĥx5�H�M�? )�Q���A(S��Mo�Z"����z��b�.���۰�Z{�5�_�n���l�MPgB���p��6}q��Ax�͎�u�u���ZW�.7Պ�����зfy8�%D��g��۩y0 N|�@���	�(��i�>�8i�=y��Fh3���_#ژd�(�	����RS�����n��	���?������jO���u��{4.�y�s�i�7�nC��'�H�M�VNM���E�� L�)lc�f�!���u���47=��a���dht�^��9����t@�ixu�N+�&�|�
�(7�}]*�\n�>hI޾@'��/Kh"؉;�]kNW_e�gC�z�EČ�*��>^~�� ���"#��DzDz�y���\vҸ��¨"���
�F���WPW����"*�A3�0���᎑��/_���]A��^��s�[ۘ����%��ې��o%��e0����S���A��=�5k�{�#��%��V�`/s�� �.���]�A܈T�{��HQ��3�?F���4��	V/��0�s%�m����+���.��N' ��v��R�Z�p5(���c����^�n�{�@����۠R��&��;?�[c��9��z����g��!_Q.r��2U�N�&w#�Ԉ����� ����G�u��O��-�٤C9\���B�IUh?� :*���:bfr�W����>O�0�?t�"�2�_
O��b�����@g�\Zʟ7f�\q�M+����������
jc��	�x;�u�u�|��ŕ^�u:��A��҇0�nWӏL���3_����/��`Ƌ8�&��'�¥���v0Wu^͙a������*t�SDa�Gj��?�' ��TK,��q 0Pw�Y���{�JH'��N�p�(�9�@���9�WX>�~��S���Q�q_�����5È+���#�w몯�s�oo��U�bI'8��@0�������ݼ+>�mq��CT =�S�1B1j[�w�O��6�6?VdE��8�<9���'O��/�,+�Ӯ�;��4�~�`�$��t~W���\n�p2ܥb(��К�.N>��J	
��ි�Hl�c��.��`v�Q��T���;�%Rmm����%�:�5�"t���1�E���㜞.v�?lYѸb7E!?~���4��T��3�{F���o���쵨Vu?�w����]��'$)?�m���|������8|Lz5�}72�*Ga��&��(���+��^�:�Xxï"kV���`�y�o製�G��u�������.K�@��5PO�����(��Z�z?[�&����o���uՖr|���.I9��Y.
��^ﵚ���!KF4˘~~m�.��k�;͎� �sg��~D���Q!8���Q٫��Nj݌<;7H������X)��'��`�u���T���cg��=qɍMH��܉I�Ip�(����	HՁ� ��Sy)��v��_E�#ݙI���lj������Y�O�XUf�1Ȳ�%���w�C�jl?��!IB�j���my	��hAp�kP�T'�ܜ-R昂�r��?�'o��O`T�4�O�
AO��[�+�^Jk�0�TuA
�}��5/�K'�&��d�*�P	)貚�P�R�g�A <�~,��-��nX�"[_�.�,�E��9���G��m|�5��ʃ(�����H�$��oQh~�;-�N�X.C�Y����_� 7�H��5b�0���p���YB�8��)��Et�H,m�Y?�ٸ�0���'��-�^�:NSfx��� /��e�pK|�_��XG���V���yXf�2K��#g�.C���j�}ܺ�Qy�q�"� �c[�Wv萦lpMԓ��a`�7ǅ��[nQW|���@��p'H3ק-Y��)���$�����?�X�;]:���SI�Juz6��O7^������VCsĹ�h��R�#��f.����1h���� ��#alq�u����ʡ�m�"�D?�r���9�<!��qws�pw%���S� -z��zP0;2Rډ���O�ݜ">;Nʖ��W�E3+����Tv49��*|�r��y�E��6�Tj]�V��1�Ӵ:���if;���	�|�27�bM�]��#!��u&�z�U/ل�[�+i�c]�,qP)�����r�J٭A&��u�c{B��ǥ;�/3ͅ@��.���i ȼ�"�N�Zt��b�{N?6�<2bN��d�D������ʵ�6w|�&���qee��㧙5��q���֑���Q5���TVw�',&9���UHn�=��[M�.ߠ�Y ���)-v+#dN[bp�Z4_��@T�	�u?ʋ�cg���Sz�z�^�>� �7i�T��.^����z̦�"� �4�A��{Rդ
ʷ�u궽���v�2&��$�y�|,d՛��=�:wj%������Y�#�Z��éf޸��0��T$�ա�d	,��>��f�cd�I�>̵��G?�����C首�P���=F'mL��^��x|w�h�����ڄ���F���K#���(J>�$�1<��qb��`)H�,��1����y�bK�ꑡ��T�Y?�&���r-#�� ���ñ�Y�|���$iXa#�ʱf8��+A;���9�e�����Ϡ��r��t���ѕ�����;��ϖ	����Լnth���K�����VQ��YD9J�\f��C��]��BMr��em�Nf�@O�U.�,=�aȂi

Ѓ{
�5(�m(LdQ-��p8�cU��l,�}R1<��B0����}��q��pw5��������R��tҌost m>�M��JJ�6}c��ۧT�&��/����4* |���$����lF���Nd�"C�]����h��!F�)O�D���*��U���gU�
z�Mg�D%\�=���L�-��&�9X����O̺$#��]�Ɗcۨ�RٜZ��M���Ml~�����2!"2lc>�2��<j!5`]��H�QZ�i�J�I��n�9eq���S[_��?�Յ%ij��UN+}%2�h��j+�w_�=c�����lk���x��~z�����[����$�͟��p� QB��O�,C��0ޗ�r"'9ݔ��m�?�nˠ7��%��MY��ų�S�x�48GN!j"k��� �����n툿$u���m>��.���u����Bf���gݟv@ݠ�{D��!7{8�L�R���@@!��:=4�� h���0˥<����8|M�Ѱ]��N��B�M���f<�;͋#��"�Y�<�?~q)��gG2�ˮ��n*�rt���fs|⿜JWI
xY����O~��?�tɡ©\��H��@�e|�a'���y��c)BH`�i	Ǧ�;�Bb`�x�b�ӌ9��"s�z��?��9'����5�������K7�M�"#�n]�Ɯyx9�k=;�{��Ϯ"����oo��n\F�DZ�]����U
 ��WC�{p��٤�w{�O�g��b;�!F�����X�A�y��It��n�|�X�|NUH��7
j.�x�u�x��#�]4(�м�/Q�uHt�`��Ar�Kf����"���u��m`��K�?�z�l�e���Ф�t.� p�GT���}�g�5cD��0�ܜ�kbp���wR�6��V��mK�qQuz�p��+F�1`he�=^E�F���x%=�D
v����J���`7LV��6Efw�l��Gnv�_�֬i;P��z�Kfx�Q�4��{�|)G24C�Ζ��[�I^$8��M�*Щ'3�4�1b�\l��ب�6"tj�C�]�y�H�0��qi��U�ʾW
��L��q'�9�k��P�Y��_H(�9��[K�'y�Nn�	��ʳ*�/�����77�ڻ�"���(n�}>���[7��i�&bñ�ڻ�4��Z�
�NST�_R.�lD�3�;I�3�"z�8�'�ێ����wY�ǆho䬗pC��3j���NP�r�O{҈�q�4�,v��������*��B�����֓ǻ�T\�/���Ar_�x�OV�,��Y���@�n��X)��2��@"��jD�Q����=���@���o�,T����ꕘ������?�kqo�k1��v���d�y����t��E��`�y�-H�NG<(oR�{�j����&�k��N��!=�Sv�I,��j���'W�nWՔ�S�c~[��CCn���F�[�|B�聬xS��C8	�T?i-��&�ꚃ���\:ǥ%y��	�f�����Z�Ţ�w�mn>^���K0�=���R$v7i�(ġ�������vN�,�l���/��	CqהLe�u���hƅ�G���衂��
��4��M�^�!h6 �N�t�'�B��xZ2��8�]�5\��gv��P�o+��i��0 ���)�ي5h<���2�X�,����HԸ�����C�����4]��hk�a 2��{k�=n!���9��y��������w��������z�+[�������Q�m�����mj%��-��zt�ŵDO_T�[��t��ڊ�n!�_g*�\U�p��~�ƣ�'��އ�5�42u�MJ��.ǩ��ک�y��[�=���5�3�I1��o��X�;:+ ��Gs����B<C?��Xw�/�K	x�}����Hh(�|k��E�H�!S!���,��v|�<fH'�C�L���Z�8������7��x��TZ�	�~�C�$X��~cIs���`�h��V���Wy�\~I&;�W! �;�U�j�V�<��P��u��d��*��f.c(f��)q4*0a[���� �=��SW�q���l�t���� �5�/�krg�vi���c�@7iAт��q�;P���7Sm��v)�4p��ϡ����2��-�P�Q��985p8/��y6,�.>�q9��[H���[b=z��d�C[4����ht�O��嚰$����H��@�_mfV3υ: ��칗W���|�����u��o��c6���+�Yt����P�!�g��=
�wR+BQ�q��J��Ӣ�G��B����\)Ǐ*����Y��j��qn��	&����w�fy��NA�%���|��k��o�}k�+�y8j홰������ ����g�b�q��(���Rh[wùAN@�F��f5�nR���щݑ.P�!Z���E�֪�69� E��[�}���D��e�qz�Z>�K�'��b����T��Ķ0�@�/��	Ӝ��֞��$��k�~�6�^���{�D#|u@�h���`慟�l��,]�ʶ��^z"�'gG���$������f�Kz��*񡡨ml�&�Z�9P���JW�X6��J�7C���*�-��u����zi�P<ad�c\ oSNj|�W�v�@/���~�yP�D�n��l�Ŗ�~��oL,ȝ����6��A��M �D���Ij�K���r
�Ta�X!�x��ݻϼ��A���+ˤ���]�������D��}B	�,m6I1)]Te�Tq��ް\�1%Z���j���N!����"|��r*���ᓎ�` 1W�h��V���}�U�'��}�tg]+�0�kM;&u-⬸�a?�_��3�ɕI�����z��K�P���} ͵$�3#d�k��@�`�P�u�����@������l+�1�.'ef��E�]};N#�L�ȯj�{��7'��0��t���Ocf��;�uuX�oa��EQ\���ۦ���s�����9բ�:/i�t`�V��o�

J�_�	�k����"�`�ů˃g����������$=����W`�LG���$���97uE��ˌ��:̽e�.Mos�}6i��R�|��5)�(j&�}�ሦx����]���W�������n��s��S��N�i��U�s�B4�SJU	`��֛8^�l��T���{_v��(NF�y���LZ�*6�������a%���:�������O�}�t1�T�o��H����k��ˑ��Dd9�@/��'f���k��{C���	���e7��'����L4@u<8[e�S%I������S��ZFVef��M�$d �� �lY�.�s;�.��Yö�3�
����_~���%�i ��p�7�R���O���M����Y�	J,n%��,��
�^�����w[����i��T�Z�pW��|u$C1����s7K�VJ(�Vn8��M/�{�'y��w�k�A��W�+�Q�4/v^hkL����%���\��]�Km�awo�_�����4?���)�p*9�� ��g�����S�ʓ�~W��F۰|� X���dh囌�{��.�q���t[��xUnv��R�}?d����-G��āsM}�A:�"�Bq�bX��*'y9Ya�r��Ζ"k���v��S�M�3�J�
��Xy�Fj�B���s�~���5mI�ćj�@GK}����CֱEI{Iy���$-M-��Ew��9z99�����Ϻ�A�G�Q<Y�I�)����*cQ������3�\�"��i�����{��S"D��m��=��<�}���pF��a�AWϯ����c��"N��ӧ�U ���3���`�q_hz3c�������0;�l��Q/�ҿ�8�#VW �g&ߢ��,R����M�}���!�~��
'� �ǃ���o��q��8�ϫ] ����Cs�f�GZ���Yal��[�%钞�2$ ��=������Tx����ϮIQ#��Ko���~!D�6W+HM˳���m���p^n���R�=1���_�C����40���u��(����xe���d��F��隝W��@�{D��7�_��B�����d� �i`Le���Փ��la�g[�S�fa�O�K�C=���a����9��fK�?N�@��nы��1#*�_�Ӛq|�t��y�ʐ���`��2B-�9b�{��[l��h�H�c9a̢��yi8�D��R;��hIA����j1W��j]�бTE��D\���3�v�:��#L�Ľ1����<���>��C���� �@�����U�̽�*�9�b�j��리�*�U��#�r~�3�y���
|�<s�R��&�ȓ�w`e���tflW�9*�{"x8z �ʞ@0WQ��$��z��1��)~-ö�MGyZ7fR~Y=?QHo������֍m�^RH�3$�>ui��Ѳ��J�ʱ�3�Q0�u��e�/�&z���Ɂ�`�6� ���V��f�=���a-����*ޅ���	�߽�d��zA����	EyI��<�n��P��M�]�~]�Q������p�;��௢\�Ն�@g���S�ǝ�����v�~^6�Ѩ	L$r� Ĥ�]`'�<Kc�Z@�}�b�³ \�L߭*[8d���
a��,�7�ٷU�7_�&����\(��԰��Ψ���6I�(+X���?js��O��^��Z��i60���B!�En�U?\����i�" �0�A��˕߹}a�5������g�N�6?x�$�9�ȿ1g4�.�b�N��y�}��iG|Ԟ쁷.��Q����px6��Z�K	����a�}�r�#�Y�2/�;��Ձ�G��XΑ=���:gk�¼
	�Ϩ��A�s%��O��R"x0���0�\ۻ�8�$�1��z�s�E^���n����`�oq�<Gl�NRet�����Z��o�§}e��숿��ӻ�9�%tjF�ޔ��A�� 80H0�n'	��y>H��۔����;��Fc���|���=A���x��}?�白;G�p�3�v�:���9vX�k���)�Y���0���vA�T���l���=&;���Xc���1@�|08�դ��#���-�zM+��$�'B�������^��6�Y��&��~a9�:T�!�ȹ�\ �lDoRA g:=��@fYYWЯZ/��4ͱY�C�S�rV�l'�o�1{���z҉VJwL����é�+D�-��K��Yf��"-��j(�
DK���n�:0, �&�=QCͼ�f���f��^mgM����@��QK��r�t�z�B�p�hV�ыܵ�D`l��D^8�^|B][{� ����|fKZ!��۾�':)��]N�)kf�]�MЎT�0����X�aw��%�\�FQ@
�㪋�a�*�T/O���J;wj���<c�pȦ���4�<?-9�O]��	��&L��ʏB��l�B�7�;3k�����g]o���%A�G���lbV"7<sR�cd��D�������C<g���q?[��'լ����@�I	�ڔ�΍�5����P�^7Y��"�	�ِ�#��5��_V�6S����2�<��Qr�D#D���~ձ�� |��y��%�k�!MD@�v#�o�]%ߧ����.��b �U���ak��8�(|�����z�Jj�����ͤ�*�5A�a�1�V^�ޙ�F �T�-�8���/��pY��Qe�S�l/Y(�U�+d���A$G1B�Z���9k�4{��t��%�w�S�����)_�X��qom�Ҫ�3_��b�ц�5��ln,�a`6̽zYcyl��������aۈa���a�
}������35�q&���T�u�
�·�W�UĪB�`Z�����vm�b1$U6�X�+��_/���!m�mRl+ ~[|T��g6�_/��$�6��tA���L���N��x�\�B�7����G;�Ǵ �B-�����k�?����{&�)[�W��s�(�.:l�|��B벱�޲�y$Eh1��R�C���Ḟ�<���F�*E�O 5�>�����Q��(g��}:6B"Z|4~��|T��BSM$6�oͷn��#Q�4�O}�3�,*���@
�N#ذz�j�S`�V>���y���0��7c^�k�yF��ޕ���a�ҹ���͒�W���tF:�����:f���O���hxqʿ�&�����
Vpq�U����Ns"��jT�r���,��SE���&�_:mꪖ1 �ܦ�Z0���|{^}j��N�d�ِtw	"��EފQm���Ϫ^�,#>�j�Qm�:�1��	5گ\�ը6d��p�u�r��U*/�K�P��)�w~FA��v�~��<�\u����1neUZZ	��&��Kj�P�{j�ƥ��v*V$�B+�Q뵉�=3�6d7���8ĸ���r���Ygͬ�IF3S�A��s����JX頕"ϲ/׈�9V�M�6��HNo�a��[,�sܞ��@V�.�M& ��ˉ��9��aҶ8����im7�Sj��У�z�;���y�m���4TF�t[Bw�i��G�m,�{�ql���9d�q��Pu[Yl��p�_ Ő:���TJ���l��s��u�C�������(��J��+�mu�ғS���&`��
y7�����P$�<�G�u���p@�;���\R��b�*n`�vؘ�&�)�� �»�3&��O�#a%2�bX��(wQS�X��Ep�`EwiC��9V8�-hTP�@4]�37�oC�;��۲��gG�pd��hP��h4�� |N�բ����MjZk�(�@%*�T�����͠���}[K�R�a`+߳^�(x5���G�`�=g�b�6��,b��"N��)Gi�;�;4Q^�T����)�HٰF\^�2��yJ5�i:�L� V���aTe�K!Ų�ԇ�?H����q��]B(c���y��l�qw=g���}�� �O1�c����H/�>Al�����l��)�����32��w�k5��� ����	�6XE��m���-�0�7��G���Y^1�\�P�I��Bt�<-���:��6 g���F�����,#����NH�6�4i�����o 7�͏���T�*zu~2(ԅӛ�H����Q�q5O��Yt�s����q=�zW�1SY�o3�$~�d��q�$9�p�_��T{(�+��M����#��:���__~c��
�$�E�rb�rM4qˣ� ��_��<��w�[pFA}Zݛ���0���xǀ�Oh��_R,�;=�t���sU%ܨ �~��O� ��['����\Bi��ŧ�������S�38���a�σ��i���H��G'y�0���ݸ'[���c�W�&��4�{�D9��x^4����1Ɛ7�5lzKp+��Qӹv�ͩ~���h�ޚbu0׋����E@kB!~����	y(��s����:y_)x�1��pV��\~۝q��ճ �۬��s!-�$#	�,��_@v)ؾ���[~+u����@����\c�l�I����Ȭk0^�`��VJʨ�io�V���-a���ť�r�� ��XkV�R�{<�adc�9��V]��!b�G8_�籠��@q�7Q��p���(���Yº��\0�;��e
Q��c1�?�VPY0��̱y=���{6e#��"��	i�ޤM��MjƩ3���;&�\��h�� :�M�ڕOq��/1Z���5��H�e�z,"��)�`�v��0�KT�Ѯ-�2KQ�J�Ķ\��s�����G��tV��TFl��b������6:n�E�e�]y����w�5��(6·q@کV���:��⇱s��B��}p���9���H���=���Ҙ{�N"�fT3�����D�*lu��V=��S��_�b�oHl;]�"�լڻ���]�c���� ��h���z(I'�V'[h�?���o�Lp�^u�VG;+Ӥ��_#��'��`?VcB��f���&�?��)ӵϞ����i��4��3��_�NPq��h\��p6�Z��H�鯜���6���10UA=4����=�U�����6|�SND�oE'��e�P������@>���Yu�h-�ץ���a��������֏dS�^����bmM����]��-�釋b{s`����
'u�42l�:�Jh|�]��� G�%����L+Bj����jA�ŭ�'����0L��[:���Џ���/�x<1�]3#���=gM�2��53O��� �	��׬��j�6�@��N�i��3�P��5�Ԣ����c����YQ��_� �� w������)�?�@J��3���|whTO7^  �*28��?�ĤE[	Üa�uǂ�
"W��j�oB�qni��!0Fr��y�nг�W��)?����f)/�<=v���->2���ߖ�T�я7
�Px�sR)J4�Ǔ͌A�ϐt�|.	Ԝ�?x������i=����v7.@דN鋐yQ�]���F���Q\mt|C�+f�!3��c@{�y�ZR 㧛�߇����a�b�x4���h'��V��2?���D���7Z�FdP_�A z��Hs���j �3A� r~gj%=���"p7ɲ���A�]�
DZ"�~Nōyq�T��	�~�|�<,D�c�L�5���r�A���z%p�4@�+��3��R���G�	膦}6�瘀�z�� )[��iJ�+_�.���D�����N�\��sF�S�G7�K_�4����%���ڽ��A0���x��!|Q���ɨ�>x�w-�n�ْ/�W�i���U��^��)�@�A�����![|	��덻n�L+��s�����R�&Й^��a���# H��#�Tg�珙V���[_���h��=�NQݱ�߫��y�zy�I���p��k!q[��q\?�ψ�e�|�s1��ld��:@n���a	p��"M�ű}�5]b� ����kg�C&�}Ufn�ð�g���(���z�gk�;*[<���z�
�DM1�Jy!���&	oh]�B14a0d>:���2�<0�g��~vj,ć��_��3��Ab�lp���EϬ�`�w�\~��D�g��Z����+���}��:c"��������r��C�>�B������IuW~�]�gs�>��n�cy�pp�I���f�{8}"2��*q�P� �#Mg�ʗ1���=�~� d[;x�d\+��,(-�cb�O���;��9BԂF��� �~'̙9��=T��8�	hm�Zq�t�Q���d�ǃ3!9R�q�/���"f�錏�J����.		=��t="Q�<���;��i�5�"�"��C����)J���[�é5��m(T��߹��خ[�+E��܁KV���9����-��.�}(���e��ٲ[y9�2���4��6%��x:�*a��񬣋�El��@t��B���}��Z5�PCF�ot�u�p�k�>�(0�Ӵ���p�"ʗ��}H�`{mc=�����/P��nXJb՛��~��n�
.쇋�X�eNTJ������+�+���5������q������؞\���2KI߸�d���
㚒"����Տj��w"���̕w�ﹺ�48���F������,���Q���P�K��r[�{��D����+B:��i�Ě�:[����ٌFa	H˓^Q0>8��b
Ec����:������R�����@2݀C��A��D.�	�����H�����b2�U/Z����͓(��燳�����ܤ,�/TV�*H�)��t&Y����TÁ"E&����G�|�FR��Ebd�����T���ϗ�C��A�3E�i�;�Ҥa�c'�E��7K�`���d��+�1;�J]�� t��\���:�I�*(���V���^ ol�9�k?u�M���tn1h3��S{����G�ِ��%ڢ���D��`��XA˶+�ے����(���r��1�l̞�-g�SֲxfU�IW�F�����<=4T�S�3�(&�d\��uXҸ\��m����4Z���ry�mؑ����k��ɡ�R�<�HPz���BY٧)�PէDdJ��Uɳl���;�K�!��&�h`#��F��<c`w]��V����8�o���*<-6�:�����h;��(�@�	��*K�nF�Hc�Ya�Dq:�俧�w�x9i�O�1�a�	��2Fo�J����m9����6行sJ����m��re��C��I{+(4}DO��R��4g3L��w�����|n�6����H����B����2��U�b׉��ݗQ��`З��p��9:)�=6�:ߺ���c��Fu��00�9e��X3;��ǟ�%@v�ɶy� 4�g��c�W��.ή[t����ڍ�戴� ��$E�������?�(�����f5�FJx.������F���츊SjA�d�x�%�>��D��n�O[��n�lO�mۻםPK�z��<�����k?�M0��g�Mf�r�X�$�I�s1��,u\q:}�^p8:��U���jV���@šS�E5B��5���s0ֳX�H`1/���1����
�� �5P᝱�A'�)�|��P�m̃��fq����5��ȱ��e�M��݇ь���w��띥R/C�G�Ķ���[�A[���L�X{���:7�_�w�k�������U��=)����^9�A�ſsF7`:�%���-��ƪ����@$0��G�A�
=�Pu��D0Xu<��UL�+F�,�o邳�
�_˪���,c�=�|T�� �d�&�i����@��V���N�nkZ����k���d>�if�`���MtW�"ϫ[=i�0E
� �<�;5�4pI�?�����"��ۖ�̲������(y���J%�\f��*U��i}m���+�ʻ�R�f�ަ�����/�{���m�&�g��O�WZPT�_��'��^TZ��`�Ƨƌ�&��^��H�^,�w�N���L:�"�
��+zǓ�����0�����>�IUS>�LY��#U�듛�Y�_��Z��S�a���?f"�M"��kc��\�KΤ�b�B�cCM5 wt���w���s[�Ү�Z�Y�T��H`k˶�L����K ��QA����^����X��+���x⛤p8�aG���R����Y0���يZ�W��+"Էá3:�[��t���w�{�5���|U��ż����?٤��̐UZ����ty�Q����Ov3��ۣ���hF�!��*$��,��V�S<	���B֍R
�ljI�Z�b�a�b��׵!9�����E ��1��CP�� ڥ�XL�֖�
��s�v�1�����3�����*�	�{��x��9�ϔ��G	��uR�Evw�V���f������ʩ�������o�d�BYw@We �pw��F�p��}��C����"^B\BR	����4��[k��<O5H�JȦ��O�"VQ�h��q+ǷgD�6쭐���j;��>M�ղ(�kc��{<�����cBk�}�3���	-b��2#m(�ik��lTѶl<BJ#��֜��k��b����g��5�ouX����[.��[T��η �#�tP�>� ���Ȧ�`Ӝ)��Q�A=���,|Hv����������o|�����(�M7�w#1�ېf��ʠ�j�Y�}���ۊ��)B�ݣ���F�;p�Eq��0��]���s�!{�a�3D��\���7��(*{��,J�B�ѴS���R�E��&"����a�֐�b ��U��&,�_D�?|�2W�5�S�[�`>@<��Ww����+�:�^����7g��x�1�e래����UR���>�z[O-$��q4Һ���J���BCEr	u�|��QìH����2�^�t��N�gSS�;���A�c8HC
9�:B����dٞǏ�DYU{Ɩç��\E��:}�G�y>��Wk),��{�9����,�M~�9db\�]4PW�,�R�5$d�(�%��`G�-��S��EP��]�w��S���H�P��X��}�t�H ����;xO�z�0�W��F!O���ű�np��xA���r6����fl��Җ��+V�|٬�e�\�)�0=�Mږ�����E���]0kgs�ga��zf���rxU�i��Cr�^<\ۑW�|kN7v�V�����us�H��Y��>�p��5��ϰ�e��A� ���@��d�s��%C;Ɯ�]�']�/�rUI�ܱ�
����j����1-�]tw�w2�i�*/��rZj�Q}��3�[�B�������8O���>`݆��[�!vY��*�Ez*�fp3��	Q�bc�ݵir��ʟ�Gc��(�����"N�ER
F�Kh�xqs�8�	�����d�N�A��P�AgAa=x���g:"�&ۤI�4H<g�.��$lB_�>K@`农�ܣ+|�[q��B��NzZ�XMM��'~� ��k���-��h����+�&�cR	E����n�5����m��1G�@:��,/O4>��V�亂Z��{��V�3�f���ON�a��ˊQ[$_?�x���d13r.�u�뵳��Ń���߬'k�Y}�1�)ǒf#<�f�4(K�{�;̐�%�=�y�<Q�N�crv���r5� y�����0��\</w;�-x$�L�§[��Gt(�l�o�jﴐB�����$�:�r�R�\��`3-$��]�">d:r' �d.4��&�.o&�lP�},�Z!ꨁ�T��I�2�?O� �4~_��~�ز)v�8�*=��XLܤ�oʐ�) �:���\��;�Q�'�I��s��*)�3�Ȱ��p�ك�h����ˆ���r���-:	�2�O9]� �0�q��c�@���K^�*�M�䜔I��O7U����~�}�cW���{x=����Q�n})s$�ж��}s%al`���	��S�E���!��n,��jeY:��^�Dz��:�C�	�w�;!�Ag%�{�H0��y~�xo�9a����7�J��7�1�lc��q��+��h��\��n� �_�R�SKɖ��O2w�c���gt�E��A�j_�s�ăTj)Qr�g���Rn�D��| 4���ߴ�KGE{́��p��El1��ʆ�7�Lj�ƤC���E3{3�(�!�K�v�ߢ���AR�D��n����sl	����������칕��=�ɚ���� k���~�@�l�"X�ɳ����rd�#ϛ����S�U��4�\'�ǝ�(Y�5U�)�t��?{/���0pr��}hl��@?�I�@��Ŕl�� 4��pg�M��ص	�X�fP�`5�Z׼Z_�F++`�����R��݅�,r��!@`�4��M�|n''�8��$g�G*��?�C:�E�}Y���ʝ���^��|򗱫�X6��F�����cS k�vS9wU��^��Cz��Q��*e��Eʃ���$���9�݉��P��xr;T��gLu֭���;��g4�ݎ �>i�Z���U��6Z��y{2���鞝`1�=��[(��2�x!N�D��&��u-@� O4�:��!���ǨDNxC��D5�
y���)���Ȝ���V�D�:�
�]�;����3��#����v�����������h� ��q��|U ���
�B?�?��Q��/���}��c�$�K���
KlEq	�y�}���c����	QDCF���b��AңCL�n�~�Ï��G,9~8�L*`�5ǧ��?�"~s�a��5c;�I�f�g�mAg�F)W��0�z?�ᨧq#�7�MFt�aX5K��A��Z{�*/ɜ��1&2�sf��o����$k�&��A�{ꍇ������?�i�^/��ދ}�_y8��d�s"��^w���ԫ�J����C����Yn����>�I��8������@8�y(1�k�s���Bo5	?�:ܠ���{4��#W.�u�'3/��&�'�j���W�ӂ�Lr�_&�����[�e\��w�`,�L8R�Tm*4���%���NW��L�ܓ4a_)�ĺ X�ȥ�2����NYn��I.Q�j��!��� ��F���0��:gѭ��H��2H�`���p�Q�+�z��<�~@��c�?�Ǚ�P�X㐿������m����"�;����塷u��y�*`�#���5�@�f^e͂�ྔC<T����@{G�ob|v՝�=
	�YHn��>��Ìk� ��^�I>�T*�+`3��FtC�R��ߤ�ѩEc.SU�������W�g�>�i���)i�1���8���3���96ٶ
3A*	��\�Xx��N�l�]��%��\��ݍ�W80������0�@|�-Ś��'�4�Kg�ם�����JQ�蛆�.��j����^�k��C��3�y�Q�W��AU���]�зM���#�.&�$�p�� }f��K�Fg�A9 �/�l�t����e�R�S!�����!��۾Ճ�k9�)���������iH�z���������`��>���T�t~7u�z�3��Vt��~�����9�����rX��#��GS璹��2�wlɪ�!*Q��vb�ڌ�r��-SP�F�e��^Kʝ��R�5�%$�_e�R	9�C5<�!t����X�$����_�a4��s�y�w��
�x=^�#c8�hj�ؽ�f�=�씲(��{�m{x�u1b��\h��X;��Za����{��u)��>��A����}>�}Ű�g -�+��)�QF@ФN��k�~�}�{���`��kr:R���kv�<��_	�|�6&��X/f{�P���+*srǭ�<Ԙ4���I���%�iq(�\�2lk0����ra��߿̓x��y� "AP�+��� ���C�:�U�ma���\b�A���{���� }��.sD�Xe���/V�R�=%7 ���P�]����W�}b:_��8�jv�F���-�����Q�����#�jp!f�0�6�g0��WxK��nb��@r���<���	�!�﬛�Ejiui�p��z'��I n�B֒��Q,I�lBe�n}RIdO�&x3݄�-�݋�?�]4G[PF�*����gf���ۦ�V;v:2юi��d���b���{�(����+]T�Y�l{Ч^<2PN�� �憕Lw_�f��)�aփ6�P�>g^���ˈ�6Z+d�z�������>Gh�Э#g>D����3b�o�w�&�z�����5��������	e.�3���V��7Z;G��ݮe��ͯ\�}��x��I��N�C6c]���J� ���P�Ȏ�52���X�ȱ��R�Zγo	�tO���U&tA�e>�eA�ⴑ�y3 Ƚ��p��{����z�
.��� =�w��
b�	?���Y�c!���h�C��vo%�������*̭�i[��T1g��j��ٕ^�.��N�#9���DyGV	�G���l&� ��F�(oԫZ��
��̃��|.�	!��֍���ϢrŊ�A!�30�Y����	�������yQ���N���������p6~Ҋ7k=��i���1Ά*:���<XˡT���#�DI֜���W*�L`�� 'R�閨�O֡�Y�'E�����+>>n�
���U��j�^0��Q�����[�Qeo��vu<!���C*��4@�G	W��`��/��N��S�c��YC6�ΒQ:�Fg����W������f�
���*���g$2Mlf�Q��Q�u[�u���`��K�D:*>6s�%K�ԕ���so�D�~b�#y��_O�(�jD�qnG-H���������Y�*&V�?��������Uo���{8l�z��XZLx#[<��C�.&)4|r�*/�ߗ�vǻ��{�Ʌ}[��@چ3��ѷ��P���o�J:�%՝���s���t7�r�1�&�w���x������rk>A�C_tС�l���3����5=�<>R͉	a�L� �]�yoc����wQCVz`I:���'�q��2�|�협Bm2��Z�b�Bv��q$�F�t���=qc��E}Լ\�W	�����4薳Rז�b>��d��		���3f�a�d����Z����G���9�`y��zv<=r�W�~v[��.�BP8�W�@~��(e���@}������n�[A��T��;�FYG���U��1&�o���S
��ό3�#.x�`��M�pX�i�f���jA讄���O����ˇԮ��rS�J�.{qo��.)�͌HnL)�5����jU�$Q�m�����.�2��#�BiDG|��Jxl�I\��t'�
:D���-[��Q-��12hD�����dq۸@�KW���_bN�6��d�w	.~���ݸ�!�H�A�	���AbPH��Q[���iruCʙN��jh�H�ϻ���\d��BIeWh�cos��H>ԛ�;g� v
�+3,9�9��,��Õ�gn9X-Z*����M����=�� ^�j�2��xG����<[!04�6i.��(�W��-�ˋ�{|����O>���Bmh<��i������z����J���:�c�ၽ�RԮ�7I�,�%�`�`\����y�'w������z=e��&p^c�ѐlqn�f�i�W���j@#R`�}�xmþ�1:�6��8���E��B��`-�8X�ŐJ�������_x+c\vqlՠ����ֿ��K���S�5���hJ�R��!x8��A�W�a�ҙ�Dx�=��KO����4_L�j8)2�t�e�(�jb�|��o"����/�jdӔ��5uH����Y7�R���/t	�r$Z��z�|�y)���f6��R��u�^*���u��O�}_!�d]#xkwV���r���j��DA=�����̽q��<0�6-�s��b/9��sF�m&�Hu���ͫ�J>Q�F��)���h"BeY����c����m�D���"/B��nE=	0䜌�.�������d5Ļ��|8�n����K�;�%U����;m����ͼ����=�,@���g�;�d����M�xrVf�{%�4n��u���� �����0��_��ZIc�;��}�3�E3�
���Fc��i%�d��f\|��C����B��?�34J+�<LC-~��[B�͗�8������:*��ڋ��:~�7�o��/�	�?��v�sN-��v�4��P#+x��2��o�@Gj����1s�������I�>%՚����E�>�:���ă����{������YHA�*�0�%��N��o��u��$���#�{04p3��	�۔\�+������Ћœ�
�a8Ӣ�ݷ�:��CWNV�3ٱU)V��3�3���@�1�9�;����_B6(��8��@����~v���Ǆ��Λ߼;5>�)H1鳺��g�1��y�<DR�~��+1Ő�m@�],DAȓ��6˝�(��Q+W l{m���<k-ۘĩ#��"�ٰ�l�!�!Y��2�^�r�I=!�Hh2�v	����(p�'Yl]�n۪� O_*��W)�a�T��]~��=+��/F̕��@�,!&8P̶�'��J�W���;H���Ҕ���G/��-���Ϙ��-�!�6��[dm)r!P�g��IL,X�ߌp��]�����_��#���ޓ���U��H���׉�����$�����hU��|�{�\�6-U<U��U�%i�����+'?�FϘ����~?�pW��u�� �y��ҾR�Y�Ӟi6���x�����*=��
u�\b�  �J+7�cZ[}�{����*�e6|
��;�e��U�~�����á��
�1���3jb�G[��3����W�-G����!@ro���0g��>�Յ�BЃF'�e�ޗ�/f����n,�� (�~Ogi�S��R3��Dwߐ�C_�b���������fO��3�ۃ>JU�c�H��b5![9j@m)�D�̨[��w,7�"WiU��G��J4/�3O�x��&�*���=�Ɗ����9���_�շFa���ؓ��T�'!�$�+k��˶g��f=��@�T�On)���IVz9������Jr�΄�R������CN��b-�p8�$��[�P{oҡ%L��	?j�C�S�1�p��*��k��iDqb�uP�/�H0X�䩁�]��&����R���v��+K�x*\2G*�T�BrPr;cT����ȑ΄�քC�I��s����_2���O
FY��/D�$�_$I�;$��Kҵ���$b���S	[��H��aK��m/�&�]x�DsǄ�P���j�w7�6S@e�4-�s����y̅��"�z{xyeW��s^�'e2�j�q�@x���V�	�l5�MlI"x\�P��,"�E�+�b�����E�%[)ל�u�l��l�u۰��6��S���{3����)l��8U3�?{�j1�����C>�>��-��@9;~3�ᰖM�Yd4� 0.�P6�7JH?��1��
5V�U��j�k�����E���.oњI���ZVy�-���b�l�A^����%k��o��ue�`�yC���E02�O�*mW����Ԗ�%��u$�e:b K��gI���>p,��g=���wR�SUr�Y��{�EK�Q��v��M�!�-Zq���4��6�zu�rU4��Q�)�������5�PV��n�f��^i[L���N�ї� 
0�#��0͙�=���2��!mNI#ɧS׵A������+͋D!��x�:�"*:j�R�IV�bMM����i�4�C%��!��0v��_׈���knw �B�2����M5���˞�R�`�kDC���0<&δ���cd�&�)�U�nu��w:�u;��p�G��c�%�����B�+9'L�;YSl�{�E�/��Ph+qA3�	�}����M��#E�7{�>Þ�ǲ.��.q��m���ȩ�������Tb?�sӀ��	d����UC;;j��AάM�t&k�En�u� ���8��@��)����>�m�5����z���I�mɂ�L�3�M��Y�&�aķ��A�'����a�Sm�LU������Ԣ�M����[��ic�g�*�)_)���g�>H4j�Қ����׎���E+���:Iw�0�� �#6j�~��_)hTk��`K�j)I)=e�ӊ�&t7�Nk�0��G�/�Q疕EWW�Kڟ2�N��rO��xg��-��W:�g��T�?087���"y�!'��I�ܯS��8<�o���3���O4���0��/�$P��X	�i�o ���^��<�ޕEZ����*D<|?Ra��]ʠkR� ��OYʤ�
j���X*���%��e���E1�A�S.V^��I���IZ�k[�?�>^�F&��~:�"#\�Xgf:L�7�hw7�O��ԛў��t�B(�Ь	�A���\��st�䳡�O��kY��`��<�����|��&��;n��mde�i�� uP$�S�����=�M`��A�!�CS"�'4�������P��0�UJ�p�a�^.���.r|�<�1ۻ'���ę�j�}O�_�u���o>TK��2�(����I�pǐ�:�P�KU���ߨ3�JO�U�C�Cc�h���E����`�l�xo/��|zr��тBH)�c��륜�Tu7�`|4�p�vA�O�}e 3x��6�`2�Q�F�]�]�5{!���P��n�=�y��%�[���>�d$@�t�F�m��U�u��!����`�&f窱ƇB���b����%c>��ʺ��We}c'M����T�M$�����~�
U%1�٠�&���L�>�A���b��n[d��=*��T��aQ�g�ʁ�.��l[�H:���	%�G��f��kġҲ��*�`ާúC;�����2E<U��0�VS6Z��8j3�#.5S�L�+[��YE��]�������p�`��7��\�=Lb���"������o�o�m[0宪�a�Ӽ���4O<��8������k�Uw��Kǆym�XQs�B��^���'_M��%w��<h�F��M�r����}�u��kB�v��S�?�z��vȈ<�� �ސӘNo$��/� �y��L�))��;�Ҡ|�7KĘLu�c�d/��)/��]�8I�@_���A��F.�6jn��J�Q�U0a��� 1�8|e��#Bl�Qc�Z`8f�c�I��N���e06��(�*�H)DZ�vZ����i���H�+����a��~,�V_�4(��l\�i��}��
���ѳ�-~@��
�� LV69a������OF���ByMñ �p�͉�Jӈ_���tŊRt'��I���AJ�ٯ�i��n7BCӬk5��Н`� r ��6b�����j�D�t�l�%ȬɆGiC;��U^�t|!^�?��d(�R»�ͨ���隁�/�e7j��r,�2W�՟d\�e��D+3pٍ�ɶ���fK�9UC�� H [ڰ<�#�)�����l=D�����+�Xۉ���@���i3R���r�dl0R/|�b��I�	*��5A/Xȉ05�=?#����9�|��S����ה/�n��N�Y�Ư)aÂK��D̋�8���uIـ`bis�I y��Ј���F��Eri'A��_L�)�|����O$� �+LRQ��[�����W�@c�L�o�[�!���D�dR�/
>���!e11:�c���[Z�Ҿz��W�lFA��:͞��)ȣ�$�(d�1�T�8/8�<��M�����U/_0C�	���kT<G��b�*.���j��bl��f�k�9�@�C����Z�#�UO�H|��2�ؤf��3�� �2��Ὰ���b�l�~��k��I��5ݔv GK��="��QU������Tzj5zpj��g�� ���6�Ԕ�URb���a���N��r�!Fi������tQn�:��ڟ��f��2����G3(?�{��R�� �r�I����!��"��f��DrP�5�:I<D��rͨ��KD7>J&�?�ʣC�H.�he��u��*�+�	M���t���gF��k�*����ئWb�/��Y�6����jR��Q*\�J��Y Hg����L� P�}FC���sG�ȞNfD��;��b� �-�9`-�5�7=5���A�r��@C�F4��1ŭ#�#��Y��w_<�����= ˤ*���#�B[�ҽi���q9.�A�QbWKϣ��E�C�~� �yи����ET<;�w��'�����vOe�#�@ێ��p�U���-j'�����?5��� m`d�J�v��5mm�͐kR�5=�� H`���-	s�`Ћ�'=Ǆ�P����}���{'=ݚ���r7��5]*��Q��K�p=�Ʊ��� Ѱ2��!R	1���X@y�]4+ώ�|LZ��g�rI?��[@��ԙ��A����jM��'Y�ѻ��^�]�E|�������n�����)��b*>"]�[%p��@-�.��a�~�V�&�{���۪��^�5�N�WLY�&��s�A�P�G�*n�"��%�ҝ\URAA4�+�j�>�#�p�.u�d'�R�M��%�!Ӵ3˼!Un}��"��; O�����{MC�x��42���}�aM�VT�.wL=`;�JF�龃�B@�#����Ig ��^��b�Q尚����Z�jQ`�|�:��0ǽ�M��	j�;ZB���	V��I,�=���6��5���it��v�:�y���72􅹾�]��:��̀��ʠ`��h���y$#�\�,�۴�@r����'n:K#��*������{e��G��@��b�� y���,R�U�0O���0v��?9Ll��*�{t��fA�4�[��9�L����N /�+˰̶�4�k`V�!� D<r�Z0ܻ��|��IY6��r�A�N�d$�xVĚ!4LO���?�#^ه��J��u�2�P�	@|L�K
��L�ۜJ�L|��T8.+�=�_n��g��������>B�Wձ���K�vJ��~���������N�����.O�-�X�i6�"��<H�~�y�c�������r��4O�#��>9!$���b�����$g�Al2u?�(r�q���Gv�/��<ҽO~�{�d��R~�gLӔ�\[�N+{]���HM�?�s�)������sS�>�4���K.Ku��hƝ���y���?�&7��g:D$�4(���}�<��,�=���
�'�/)�cGD_	���!_�I �`Z�Q�	.��@�u�x~��B��箵���83eG���i���曰�/�ErQ�Zp���2�#�@!xH�����:��(W����#��򬪀{
��u�#�+�s�@e�a^>�=��%��#%Bē�Ƣm�ڄ@Z5���q����Ų��:�͛��s��^HI����Q%'�z	�����%��E���Q./c²|�&[[��Mm�Le>��1F��Ki�.x�]�䔀{�X>p��K�����T{�=7�� `���a���[E��%�B~g떤������r��.W�-��,`"X`K��A��FXCi�!�՛�8�˘.j�3n��u�*�q��H��}�T�]�\�Ҿ_ֶ�P��C�j�XX�X}m#T��|�};�}uw�S��3�%��RR����P=^w��1ÃIBN6�c8@k���r
p����?�>���dC�t��H�[�V�0��n�C��m��7j��� <p.�	.�b�����uHZ}�A��Vs]�
���a��͏]z:q�_�1�����?���O;N�?W&�8��Dn� �@�w ��C~{]^���6�wp))}V㤷��Q��=+03(�G���؉hNAE������d|��'���q��*�5�����ĕ%�i��)��%~���/�+��w�:�UV*��ӈ�-���Nn���&��h��k��1!���EA��uå�p��B����{~�N��c�EH�é������m�� ��!wљؐ�RC��y��D.��~܍4T4��Eb���;#xvg�����w{E:qz��_t/B-1+/�*~�!�U�b�X1�~���e3���Ǜ)��ևG�ئz���e`"��8�~�����"�?[kR�<-oeO��`����6�D���d�J�0A�:������Q;�p�9���<��uM�.o�'�'�p���R}	!��2H4�\���9n�8�_v��d�;DGgS	�5��IИa���õ�sf��z�`u�����["B�"�mJ��`"ˇ�7u+�8� `\��[���R?��77$�R�6w�ܦ����Ԃ���9?�	�Z��.��|v��M�3D��i\���:[��	�qZ�Eb���˨�_�$[���ɦ����N\�?�(Coa�B��~\X�G3��:{_�%�cɤ�@�;���$��d[�;lk�Rg�l�=r�	�;3��x��N؂d
I^;��s�U]��%�����e cc��Xd�������>���e�N�HD!�3����J�I\��e��'�p�܀�6��Y� ���=�� h���������/=tI�*�yx�K�4d5w��[$0E/q7M�-w�$�
C��?���w��CT�"+���a�FP7.�]{6 �z8ax&�q3� �X{�b����+/�#\[NrG���M����
M0�BIM3Gϼ8����l/C��]����3J+ Ɇ�r�D)�R9xt�?)����b 5oS*�WϤ�i�"�<�_��t� �bpr���R͚dճp�x2i߻6��W�կ�(O2T׫N*�@�%���Q�a#)����ySݝ��X�N[�h�n3�|w
��
C:�1z��Q�P��`�R���oJ/�4~H�F��T�8h�0�Rf�����Fډ
�0�;�#-4Q��p�)*`����^:rD��[�Q]�<�.�8��P��>�U&ޖH�Ɖ�a;}�9���P�1�Zr��]{.�r(��C��U$/\f|�`Z�£&?�Į��&1��J������}�ڔy\��b\(U�ܬ�pc�����&dAΧR�8�n�R#G�u	XG�� s�5��i���M�=)��C������zw1�d�#�G'�p�mv���;�b*Jj.��ؿ�Y�_��!1��?��A�}u�Hhv�ؑ�6��y���&����[▆�ɪ�dc C\�Ĕ$D��
��@IF$��=�R��eH󄴣0�޽�@Jpj��΁i�wT�P���w�t�]M�fdƗ�c���Y�I��xh��ͣ����jB�e� �;��b��;�������%F�'LT�Zǒ�
bK��*&te�Ƣ�@�H�#�R	�L�q��Re1𛆊��JXK�zs��7D'��,�E��NL����@��0�9у�1O�Y"9��]n�F�������M���Q���J? �� ~sW���:��ğst��+D��h�K;����_$)�6c��ʿ:˭YΧ2hg-W�Ga�|�Y�U"@0���DorB �>�K\¹wó�D>�j�$��1�5�6�g)��z �kJ�ǚ�-o�}L����fg����F�=?�Vyϩ��2�9o04���i�1#!MG.�a&=e`��WW;�N�+DR�%�N�R��|E�����PC�f�M�Ja@�8��21��7>v}�Z�B�c�'���{�^����B�q�J��8�A�@7����2҂5�V����˳R�nW[#�UO1ё��vT����T˔7����Fa��$w�����I��єo7�-D�>���@��r7�jy߇�7��t���	u���ohc̵�Kg�����.�e���f�RH8���n�@$�]S�q8�S��CƸ���H��<��Y�|��6�H�G!��-�����\z_�	|��(L�'il�	����tۮ}�~��t���T9����6��^�ަ�h�Dx�}�"�t�o66�Zk��[	�������� `{z����x�t\����p���-�
�_�\��L�y�}�ժ��FPze��-l��h0�X�2�R�:�>c��xÓT����w�3��3ط��Se��e5��XlRm� �sJ�"��u��d����1�2���"e#��
So���%}��M3Ϳѐ�f�»����?�_z{~���o�,��
���0-�I+M��a�sl�u]Mh��UV23�G�4듗>��b���������G&7%�P�Z&ڧw����p�6��r$ƪ&�"D	� �^_I�@@>���׻�ɎW�,8��(�4������eW	��v�l�"�e��:O�8�N���;�o��ە��v���2�g���5�8��Nj��UC�1*�J$F_8W�|��J���� Dq�<�%�T���G;��$ĩeV��t���.�_GZO7g�Ȼ�|9@�m�8G��`vJ&-&͘��M�*@t�i�inf�jҫ��9�0��"5��B�ǼH��E�"sT��\z0�e7�eJ��+�Ϧ=��?½qK�KÔ�@�J+�1��<�0�O3�C���C��u�p,����x]���B��U�k7-���{\���+׾�V��?�˾���Me�G���?�Q
rؙ��Ul@5��6��9L�i��:��I�3�U�.IeҊ�ex�$����Bm�A��F9�{>���kkCz̎� %P*�v�鼩�F�b#W�c��Ƕ�Q�B]�r�!��)�^�/v�8��������=���P`�=7�gU��$���<��4׎���@����
z��e��~��\͋�d����� ��T��������W���z�9�]ۘv %�|���9!�(,��}�T����-�ι	�z���"Y�
Ё#i>}e_��})�_��ٷ%����'�Y��h\nm�"_���/g����ϡN�`�@�S=>I��[e��j�)u&?B�k�᧱��K�H��⥮�k/ݤ�߸��]/�\w�y'�p�O_�x2}�p��c�V�d�?�~��#�p-?.8A��J4��|���H�|��
�u�����XV���������svV\k�>IN����BR���#If�nh2出"��CJ D��v?�r�.�Ц��Rg(�ڇz��֛���[Q�+條MJ� ��_L�G�j�7N��+��3
�i��T�m^7�[��j<M�SKU�Vv\L��pj0J��ڍ�,�7�z,Y-��r�I1Fg<83d$���`��ݨR�}��Z�Ih�2/H7eI*�ͅ-��G%u�;'�9�P�e=�J�^��5&�_�e�����<��x�j�[���ⶀE���T�5��jߒBa��@�TƏ��Zr@�>ƚ�q�%�Χ"ZۇGX����k����۱�w)x'"s�S;���}>�3��5E�'0%�G3A_�H�H��|�\�9�Wѳ>�S�bd���T����.~ɘԠ�")d�v�x>�=��$߆)�� A~��t���^�!����wr��Q�0��R��4��!���4�=�X\>�K�};`�y���p:ƐH�ܖ��c���Ɲ��'��Q�����)6� n��_��1�6|%v�l-�W���[�Ǽ�VJ��{�F
�v��x뙜�Op�\�#N:8>��)C�,�n�!ݹ`K��u�Rڱ�a9 �e?��D,�B,�lő�� �䕟P��{�%�fU��w����unf �5�KL���*e���44�"����*����|�&B�N�W�'�,��&(N���f<\|A�fe ���5���z�U����R�޹��p�cT�������[�>���f��e1�C ���6���}Ͻ���
Uj#o��fo����SS�v�kA1SW�Ό:7���_E`'���[���r߫��w��w1��ޙZC�x���W��2�������Ĵ���8g5�sg���D�9 $���N#�f�w��s*�3���B�!�y����j�}C7Ĭl��r���F�hD��
Q_yM���^��`$ND�U`�`�B����^$�n�nt��<�z��k�"���_���rl'�����7���H?;(��_9Wt&oQ�0}P�)�Ŧ���>����O1>I�x>8I�����l���O�Ly	Ǟ���D΢aȦT�$�]��S"[��wQʢu�J޿e������������l+t�l�ni��S3q����3�N�@�D�-��i�g�4��Ɂ>a��2�He_Ƶݝ���X��>�>a���?Ac�����j���Q1���RևǗ�?>zXg�+LG�	�������6q)p��_Lb�{�ѵ'�R�Hd�vm��>�%���v<�s��k��"0qWU5R9TNrt��|f���0̀��UN����N�>��z�(T>n��,���wI}�^�dr���o�W�<��O�P5e�}8}�<�5��4ɡ[���*4E7u����*�z�m�񾰡�d��4b,�A(�"���.\�L\��$�e��uF0�t�d���=a��K姵���b/-řV��t�����2ت�z��|���߇��[�Ɣ#�� %`����8ȕ�����~z�qٵ���:id;����S7$�Q�'�F_J܁'�B /-�zB��l��g�=�}�걶л4��f"�=H��ɡx!����R �6��Ag��Gz���KJ^?@�yl�-�o�d�!��5Jy��R�}v�Ϛ؎#�O���~�-�� ���񸸢�� �4 �x!��LAR��A���h���[�Mާ��!����}��ٰ�l\_&��uuО��ێT��!�=�oj~b}K?��F5��^;����,�f��Ζ�J�<���zmE�[6���\a|��*@�.rS���m~���67��)�)�G�9	�!�DX='��b�^i���d|'�{㛱ց`Yu���I��k
�y(��o���6�$��݀��_qG���4��/�񪲢���_��R,Bc�P�N���(�`��J�!�%l;�1c�!�|`!��W�N�!��O�A�.�iI�*���2�k��lv���~d�Ɓ�fQ,Ou�l����',D����C����PlD,y��@��6���m���x|��à��
W_w4�O@��28C1�*�لb��)�:iV�d?d�m�j�Aw�6�"4��K����y���x�����:�Yf�n`�\��F&B�y�ۓjۼ"�"���1��A�G[���><m�����h3%��gzr��O_����QKH�3i�mN���z�%����#{�)�W i�5E�2X�_�����*EG3r*C�R~1btC�x��_<��T����W���0�lT�:�4X���?����JS��&8Ӑ��<����r7NTM��\~���%?�/ɺBPD��:�m8 C��0F �h�0$�*Hc�I��ߤ�R�T���,*;EM��ɔ��K5�<'�&��[�?�U6�D��ޑ��g��'�n�-���~!3uk�����4�1�K��'�Ҳ�����W?^o-g���hFc��N��OC���IXO�/ �m՟��E{6ʓonm�>S�u�y��g�1�:�*0�T�����o㬋�x,����ɔ�8�1��[����1��cԶ[�����gWX�Î�3��K_�$�<�����k�w���2� l�B�⣍���k+�|�4_�|+�ۤ=�3��p�fK�%ʀ���[������p�w#�b���<�˪��D���i�y���Cb�:�V_%���L�gR���G�٪��Ϣ,K��Q[qG)��x�g�a`dq۫��)W|��)�����L@�h�0L�tgM�:��=�]�~�6���I��m:��²���v�����7���Z���S�{�Ra�6b��4��z�&˖R�O�����*'��71���[�$4���h�I�ʇp��H2�nq�v"�/r���^�Uv�Z{��i��k	�8(�8��m�b�F+0�o�Qe"c89�SϜ;0v��^�'�=Z��3��9�B�g�0R*?�FӖs-��EC���6W)#h������#�N��Άc�Θ��Ӱ`1IM5�I���^�س�F���͈��hM��@�n�3!�=����w��F�HtTL����/���m�ozY	���F�D.���c�@�v�p]=�8:�(,:���]�*�����}���%��6t�f~El�'������An���=���EȎ{թ��\C�T�<+~?��/T>ig���܂��l	�a�ɵެ��С�?���"�E�%ep F�2$����ڵVB�����U�o���m�ۅP�՘�9q�,��L�b7�6��I��N�؇Q&�	�p\�dDu�T{
s�V1�!�R��`U��֑�T�q5�v�&Y	�=�Ͻ{um4�Ud��/T��&a�g�ە��l��b�����6�����i���f�?G~2�5rӧ�R�[A��e�3_���KY
 6�7_�aCF�us��=S�W������a��!�ա��Z��ur�Ip��V�|�y�*�Ԓ���AZ2����J�o��2��zn��1�U���f8��Ya�90 0'�ڑ0d�K>#L�O��|є`�*�G���c&H+j6��c�	�o_{�5p���\qCП�j����Qo6��7��~
ުQ�U��H��-	����"���pN������'	~�o���M���0�9Ɵ"Sq�+�զg�uxU]8�@b�� ޝ7��Vv�hj	j3��:�n+�Bk�--^j���=M-��\r\�C:Pf����61G��M��3��Ϩ{��}���`S�<�'s����ߧ>�P
#-��n{��UO�g9d�>u.2��d �t6���z�����7����W�Ml23V�hE��S��/4�M��5��zX0<�(Ȍb������N4i[�����ay�M%C�cf��]<����T����Fj�_��]HM(L'ð�c��휲�<J���.6���A�ט-�i��F������a��Է���ט����jўP���Ֆ#���cNl�c�.��.Kۙ���@jr��:w��䟴<��X"��\3W�k}.����c;�b%���-���%�TVW�*T<~�8ը�4l�zi$*Z�2�����*[�]OH�Y?{$�7i��C��t~�U,�To�=�dѐ�JL&�4����*:"8�'-��Sc�77��/Ӽd�6 ��t�:�zƥ/���a�=KOz�&��P.���y��_F*�K+����0 Pt��A'^�s2C�",NJǀVq����a�?pJ�ynN�������A�����j���p��ۥ�g64�r�����Rl:Dk�����}%�U�t�F�Lу�D�X�Z+~	��'�k%G_�YP̿k#��~U�$�0o� �
}�+�k.1 ���S�[�@[:~��^�Ng���E��#0k�p����|���ݹ�W��޹A"#�ߗM�&��Ѻvq�DvM�`괇�t��
���8y �EQ���b��0�7D2�����B"[>��A��@������N%F�%��� 4x�B\e��3N�]i�I��q�7�Y1C������C+�V����Pά -X�]��R�׮�@FP�ם��֥y��H̡e��>9`!�0@�14"�#�=���4m1����b� ('H�&^>o�7��T��!�Ol�hΌ(���	����Н��?fh�p�n��� 9�Ǫh�'^�ʊ����EG7�M��2������ˉˍ����^�`񣅍��I��o��\uRm�8>���f����л<��X��ҁ����.��>Ϸ�/-�e�������>	�a`^�F˔��PBٍ+�Ӗ�ߦ3v����&��$q��\��^��w�ӹ�G��WT��$�&md�G@:�W�(���� ��e��\E��
j��j�g=:���'�:WR��;���y���Uw}�^��od�V�s�~H�Gr8���ʶ����'��g�g��9�����={����$�T��	�w�-,_ǘG G3#j����o:�J�᚟I+O'~؝���qG,`�7N��g]�r`n� +R�JtRD�isc�c�_;�b+5�[��=a>z���Vǝ1變����V�θ�ò���)sZ��J:�7�"�?��a�Oe�i�D�"��B��~C� ^p�۹�d��A�К��:�#<��&o�늊�̛=�?�
���9��[Y0�!o`����g�
�QO҂?�sizOv�) wgЧ]@��5��ߡ$��!�P�S��mg���/g���h��Ϟ�Qbh�}�ƈ6N��P K(a-�i�0�2 ��)��3f��]�1����9%��� 'V���K $�r�Ix(����)��+)�g�<�-['9<�� �����U�������<R���D���b�\W�=�
k���q��{���s��6�S�h�ػ�{wv��B�(wʆ0��=fRA/�M�
v����{��&�ຼ{(�����S�F	�7��V���py��=��@H��#��e+�S_�r��\Vn2�gC�s�k����hUt��]{CB��y����{���5���]������/-�eK�U�t�@��8$MeĨ�*e�&����F�)�XF�����������0\]�5F�pY�+��iV�^�dJf�+��4�����7��o�,`�[I�ۧ�Z��F�|�d6���-It�f=�E@�%��u���p2!�`�p��<S�b�W��,t�}C��1� �,,���Ts,/4P�>�p�CѢ[)(M�&A��gd֧[	4u��]��c$�wfi�{��G����1v-'�@<Ǹ}�˫���籱�I�D'V�W*���P�������l���F�.-���{R2�]�)���V�ہL<����D{'�� `��x�e��@<���� ���i�J _B��#���GpF�|�e�v��b�����S]�D�����7q��{��R �p�8��#�lܝh��� +f�-���"Ô�Z��Ģ�"�;�6�uO��9��(�uC���o�%�CM3���{���N���	�ҫ���:�q U9�L/�I!�`:���;�=�5��a�ġ���ip�Rc�]��beK�y&���E>al('ެ�ko���b�洴d���2��]�5�o�{�ܖlv#��o�Z�l�^+ZfL���P�ۛ|oGU���8�w��4�(:��wI"7��
�L�u`[�5���Z�U���V*X�q2�J�7����|_"3dN�1�I���9��2bl����^E�x�T�bO��o�1�b!��u�Q�vv%* ���U���Z�bU�f>�v6,w2hF9��Cp���<��5!��䪔���,"F&����i�K_�,#�*�_�'R9�g�"N�q���� 7��=;)ܝ˙H�u�1�'�E��8rN�F~�')?@�򓮤�^82z�j �w���q�v�1R���>qS���>��� ��Yi�5v7X��Z6 �u�ߨ��Q�Ba��:z��ٌ��E �H�"��٣x.�!���h6�?T�%��3#�L2��ڄ^9>��T��-
8�Ġ��q"o�b����p��+�^>^U��>�Ʊ����A��`-� !���~����Hze!kRYe0C��,gT�BU0�eb�,�r�6����
�z�K����Iҡ֝���*kٕ"��/YϷMbܰ�(�z�{�Abb�&K4��wnD��K�9~�Fߕ��]4ϙ�ۏ��x��aH�ZeN��&�".�+b�ӘS����	�0����3N%J�x��I��?B���PUm�u��Td�����CΛo����G�߹3*1��s��N�§Dt�ѻ����s��v��)z\�����rU�s��~�-)�dj����|Ⱥ_�N� P�p��������os����gs^1V:��5�t��7c��kYS���"����K��Y�Q�_c4�¤�Lo���/��m	�r:0"��7��؊�'+�+�%��0P\��6�������P_���شɇ��]f���^k�����f��˼'�W�s[�<��e�G�>+qo�{�Z�l�.Ǯ�k~O�6���M�����]1���Y�l�y���b
��c��`®o3�ڐ)n�n	����%��a�QF��wީ�����J��s�ƮFUf/����J��bX���+�4@��H.[�-�R��2�ֈ�r$��2j^;ۯ��g�z*kq�	C�^{~�Q�j&k�ʆ_�V�	9�J�rm�����l?�!�'u�P�4�ɉ�NP��
�AFuch�%�zq�:�n� ���Ԯۇ}��p.�z%���I܂�Z�ӫ?�;Uv���b�S��*�8<���R7`\��\�.�U���֕��Ԣ t�t��������*�bۃ��i�p*5�װ��iك���v��0%[i� m�S�{��*�A��;�G�c�h	�?�-IV�s�t���rQZ�3O���Xڔ�P�<)&�T��T�E�|���:��`
��Q�9H��n�)6�OQ���՞_�`��ب~��0��\�[�Y+d���QpW���ұdN.�£�<	' P�6�B®cm�ZC��E
L��I�D2 �o���Kk'Yl	��/�ݓ��P6�eǍ}=�p��]����=�\#���۽�c]�k�+Y�8`ى�Z�sZ�n��Tn�O ��"�T`��,L�v�^֌�=K�%�����)y�4�e:��ξ�7���C#�w%�ë�:�������),�o���eW���BC��R�܏�7�5�slXl���,��cK�t˲b�pB��3��m=���%�������A�P
�Q���2ʺ�s>��~������=:��f�Y���X�Sx�+׫��2�ݚ���!v��;YU!ɼ�����P%���b�~*M�3Ѩ��c��lw�H������Ω����$ƺБ5��g�F�"��=�J�=�>�DH�,ek ��D�H�Ϭ�����^���h���Q:�\v;���}�A "���8|���|ʱt�!h�Hq�EH�}��m��v�O�aѳf�ɋ�b��X_^�4�E��(ۧ�� �m^�+Z�//@�i�}��N��exF�L��4�k��F1���go��G"&���n�9!躌q�8��ΐdҏnO+�ͲG9����,� ��ԡ=���*/����☍�Pº/m`ro4T�%�_�W���\��P=���Ԇg2h��L	�nN]Vp�VlR1Za�V�dBϑ=����ތ�[&�W��m�@�¹i�?wJY�g=�ڥ}�[f�:�&��[4�{��/Ъ�H~�k�N�R��w?i��}��R|�Y�j��k�.���@�cc��.ӛ�lλ�t���9�۾���]��<��o�5-CwmgB��aD2Q��A�s�{���I�r����-�i��\�u�j-Z��H�˘�k�?�!X�ĸҟ՝rs�@pe%$Va2�'���	��wE���lؚ�"y)���nx��?�:/z�=���_����M7��;^����6q�7.�s�
�Qj" O�.$��Xx
,�	/J���
���Z�j�1�sL�~<�ȍ�̹����DOOQ�($o$�v5� �|rWu��^�{�PR����<�W�nQ���!����\%��cj��w��;�߅�=[��HqNR3�o2{:���La�uB .���(���y����q�ڠ���u��@_m���YC��VP�"ۻmV�-h�4bpO���]έ�:Dro���Y�
j��'� 2���-��3���"f�N�^q4H���㳘�.�V�:cY��]��Z�i8��*S�~��?�Q�k�t�� !��7�;j�VL�{,K�����Rܑ�7�����b��:h̑mY��5z��_�Q'�y����b	� �;�k���b��%�5�O���E��%�5j�?�L���#É&�ٽ�l�D����1�o�j	!R73��(�u��M�Y��L������ԮW�44� yq�/z$s4�Hb�l&����p��ok���ܝ?�0l�,�X��֯�ƃ�PW�a������u����@t���3Հ���\��$H4�K���̀W�?�W�0������5�/���6��:�O	FS��խ�zN=��H�f����C�85֔;�����H鶢��_��6��nV۵>�fQ�p���:�!�d���k#�U� �C�����8uZ�(W��kSW��ӅL=����}8�
򙹋����c�j��� �Y1�2���cϹf63�(��%8�����+u�!���g���b�2�&� `T�޹��^�9�eX�bn9���|���?��8���\���"�}�$�ĉϱ_(]��ϸ�����}��#���| �h�ʎU��70�dc�*;˵��Z����D[kL�m�?����Np�*��8���$���MHl��� ��"�=�	7�m��&� ��I�S��n��l����u�8V^�
4�A�|q��1�ch��o��Z����e½������c������e, +ҽ��.5cV\\���� ��6"�NL�b�zz��()Я=�W)D�������xry`��YvE^zʏ�����pr(��z�(����"�������O�~D��̫�xve��\F�P�ȑ;h��|]�<4ky2�vs��4��@!��r��/*.S��!�?�Ͽ!+�Ei�O\@�A��!�{n�@
�D2fDD��d�Ik\�V岚:��Fe���+%dq����b|���j�Ul���+�7:�N_�����d��ܠp;ҍ;F�&���a��b�T���8�l*d��I]\�P��e�9�T�����\��T�^:��!�����9�3���į�{���z�L;�=w�t��0���Z��ƅ��{�柀w䜡4���g`B�T�۽�9̄�q��OЈs�)Lf13����e�*��{ϵ]��=^�[t+�I�eu02����P�T���[�F�L�yƹ��m����&� !����Q��2���<�=�c)���,Oh����������-���(*���)o�V)s������<@�e��JQ�_�U�y�T�)�I�ސ�j��m�O�?1
����5<˼C��S��`/#�Ĭ[R� �҄Zm�D�z�A��� #���[x6a�R\(}V{��w�~�I�U��Tց�V>�R�t��$�$�@A�WƯz�۴j��Õĵ'2�0��Qd�"�T��p���D�'�_ղ����)�K@�g�K~�5��ǵ*�2v6X�^Z�&,v:�.kz�H�c6�;��&u�����b���F|�U���s\�̃�փ��%@�fU��8Hge��bxLݸ���-�z�������EpG5��E�xc1H<��Ϙ��G�g^02i��k�3���P3B6��X�J%��s�8G�������{P��d4�4�GxT���&!76)ܿ6�W���KP��C�[��y���]f�u Ąn�` ���Q�q�|�2��u��<�E����?A��F��"��$?����$��?�Y��J%��|�L6��&B�������t��@o#ӵ)�.�e
��7���͈	wf��
u{l�z 	���^�q����:Q���O���l!9{Zs�bCˀ��K��҄��w/Q��k�	�%�N�қ���'T�E�� �:1s��L��h�GS��@˩W�6�(���%�N��J�6�}h���=v	��[�!`��V�f�Den�GPܵ=8J�|c#}�:p�Ȼ�2 ��NQ��" ��!�	�� |�+yg�ɵcvW�.]�#�a�B�qy�6�L����K%�n�vFns���˪H��.����r8[Y
��,��������.V��Gd�]N�h�F�}����B��<ʺ���\�����'��y�H��t�w�{i�80�#���������Z�z]�|�{�Ac되��k��=�T�1
�a���Yl��K�Nu@�h��T\��� �r���AJ�x41�;����[�r��\���|�&KJ�Jh�:2�1�6��S&!�઻X����n}<�*Q�Ѩ����P��p-�z�6���_�,�jYU��r�m�Qœ�8Kel��� �S���X�i4��t������N�z�B�t���<��ra���c�v�V\�O��Ci:�E?YM���1�ѳp�0=�	�R���g0|���Z|V�z���db�����S����?9ߔ�m�T�3�:|kՠ��kc����Q���J���&k�-1C��Q� ��"�UmD6�T��N����A���AY���"���.X��(�y����F+�B��� UQ��[�<f��n�$`��H��}S',~��qd_Q�I���=��(&�zY�4B�X���6��^>Dr)L�R���_��?���'��&ѿK�������[��J�i��5�a_Ɯ�A�~�hK��v�یMJ��g1 �S�֍��6#�ј�qk�^KzA΃�gaQ�|�K�� ��1M`�%/l+e�d���D):�ޮ���n�έ��i�Y�2�q%^/���w�Q��I͌�nEmb�W����]�
ө=�<]��@e�}Ы�Ay�_M�e�]ݍA�W���y�=<H9������_u�d�!�"�bqof��|���UM�H�ޛX�K��l(�k�K�+�qt(iB@A����Wt�~,�l�Q���n�{�@���g4��<� ��G�k�O����8՗�ܰ����P�gw\�rk��K>"�7��H�1��82hI+qt�SG��x[�N�Mۊю熸q�</����C�"sIo��_��7�lI�Z��}x��#�y���7b�.bos��6Hԕ��t'��%�jl1P�u�آ?U���Ӌ���1p%@�x_���c	q�o����s���!4*&�@j�.#\QdSZ�C �J��6�-�y������dpZ@%�NXV�S�5R�����rb�=}a�չ�T}�i=����>��`p���kD�5�O�6�|gr�x�k�׉j��K�(:l�
׊ޗ>.�2.�N�� }ʋ9^�5:O=��~� ��Ŀ��|���>�s�k���6�� 22M�q�-H4X���f��R����S�tٍf#j9;*�Po��S-=)G��,k�.�C�o�.1@g�<�?�O.nx�ض]F֦y���t��t�xsf�AԦ��Oq!c�$�r͍��H�e��7��H�+�AF["v�uXH�]��5�6n���)��U�!�����8-�>-�i�:�Lz�<�?'�9�b]�T�����*'5����[���U���&�+G:9ͱ�c:R�υR�+�6a�Jw�ȇ�������pr�O=c��<]k�r5Ч��q|%�mE����P$��N_[.�l=t�J��v��,t�?���G$βt��������
a��yr�5���A
`���y���9&`0�}&��G�}�Lm�-���x:�kPW6	��f1d�oX��`&�+���l�s�$!s�?cB1����O��_O]f���~���O�A��5ɯ_Ab%��;5x�Ona�]H��lXU�ļV�0���p��l��k>� V���R��y�݌k����M��y�ȳ�ʾ�/���>=�W�R�K\�!w�X͂��SC�PXq��m]
���#J�Z�=�t~Qm�S����OH�?*R�*�A�qC�Co�Uh=j3��f=�b�i������銻J{�A�D%��#1��+������J�-��-ozaW�.�U	��@������[j]�d�i��g�%|߰�L�:Si���DYB:�5R����������[.&̵��;{l��X��u+B��u^��n�����eqi��q\G�_�V�8V�u�^��锖��$�N�@���=�0�a����֢ ����m����.CA����1�绘~���푲�8�{�`U�����'�r.:u�^y �|����|'��Kh�/Z�5�ٷ7F�1#mQ������X�gCna��lv����n`FV&ml�8�+���	Z�K���QO	��$�J��y��o�~�9��!#<�t�3n��5}��B��s�p�=�ۚ,Yk���IC�U���Gxn�W��a���{�ן�.�;<�E���-6%�	P�4�N�۠L�ا�A�:�8F�ݡ���W�=��{�W�#�dP���e��aR�~��H���宖uE��m����+�r�	������q��� |���	�4I�*f��h�]#�#�z���|��T��aَаH/���J�҆ݧ_w��>����oo"7����Q�q������{:^��I�{u�n��7ɦ9�-�h�R@r���d�z�k;��]��neًQ�7x����~Ğ�%5kv�̭F��q��&�I�U�#�.'�/�b�8�VP�VϦ�*|P�`v�Mz�Eq�eT`_&�S=����1չ�FFh'$$ʧnwq�}{�}��gF�xzoM{�z��	+�?����s�f.�W#F���BB|x~CH�^�"F������6oVD�]at�]�� L5?(cH��-q�ے%3��*:�۩+uvp*�bۍ���.*�@+O+��`*���?'�3��Z,fWh7x�,8���t;�u|�W����/	�qM4f��T<��ХG;�y��t��x�I�6��ϙs.t =��Bi3��a���e�!�(x�$�����1�N��ߗ�ُ����V~c	t6&v{/��%xhILUcn,��>���t�[s��=���a>ajh�_@ƟΒ,|ȁ��&ߖ�gн�	6��Dp��C}�/~��'@����!��l������(�S*ߊ���ƫ�����rf'��1k�ыGL����Bf)
�q]@AS'�FI��М�
���W��;���o�F�hX���4��d��s�ʦ�P���zԀ?bF�<!��ĞiZd�1g5� ��*!�'OH��~@R9��;���WB�;�=:;��J�8����=�Û;��ϛ���#}�7���G��:�-�nM)��='.&K����f�Z�T�=3�c� ��L�]-?�5YN9As�*7�
2�2E����hz�$K~.w�zTQ�q�GGw�<9�(1(ǃT`$iˢ�O�����r)L�3\Ѱ��F�Ta�BF��&��G�H��]��	�Y�,}�uqi۰*"�P<�J��:��j�zM���������P���{֎**��`���*(�����V����sS���
�o$P?xm__r�X<x�n��6lH��}�?���5�<4�����@wn��pO�i<`�a"P�IxX���xZ'5�R���џ	.��o����db�\�6X��j��a!���J��N�Oc ��C��:�>�)%��M ��*���������ׂZ��hĆy^$�o^
��E����y�s�ZC�6y��~�+C�$qj�KON�˅9�]� Uه2Pu���M�iL7�ڞ��1��:�z#
���ƞ"j\5?y>z����f�g�,X8q��/g{���MaphA�o=!H"j�F5��*��s���נn���oʎ�~����w��f=�l�<q��0H�n���97�g�N�2*q��j:�{%x��D��?�G@!���Y�)���|2Ά��Rm�EP��'���=�	l�kM�yfTWS@��11x~�k��8���k�f!�d��
��3�+�gͮ���^)zW�e��f�A��>y,<q3�_������p�Oq��ni��ݤ'!-k��tt�U����0��TR
�3������nǗ�*p_�e��R.*V�Đ��&"|K����gnc?NK��&z[����7#�Թ?na�]��[Ѕ�:��r�>S�}3�)���\+���7�MY.�8|\��#)��4�`*`�1dU�P���̫�O��(M�<2Z������
,7u|U���@��c&��
��Q�'�བྷ�d\7�Yv�� �k�����k[@]ҲN^�Rpf�藳&~�>Ze�1.��vfW~!�<�r��h���%��ZO������W���E��2�����V�eC������>��{b�� �T��/�$�0�8�)�1��[Xm�-� 	%dp�m�eO1��Ef��׵��5CB�a#�Mb�wn�'\}��� �:U+$FZQ�Ԧ-Ο����R�#�tga�Yfد��}�*�������D�����6azƖ�.�]�a�Lp"��Aɞ~��3��#�#s��2 X"��A����w�'X"��D\�����z��gC]Sx�k�p/X�#����ר�C���C�"z�ٸ�R;�?��Y�I~9a��e&��}�lQm�.��D_a_�#����Jj�l���
�0��2����s�� ��T���߈�E�{bHES��C�	o$��L5��orQ��?��^��M~(�b�y)v9�)*a���,#%iS&�}����_7"c�{k���n��_���������6������2�$z��aWl�h��f�Q��v9����a���iQ\Ǎ��@3c�T��&�{ny�6u}�3����(�t=���q�ҵX��X��'z�}KWғ��/A�C=�	���{	�D�����q�|"mظP�GM�b�?C6jA վ�0)���wH��-*�sE��ZΉT�CQX@R��j0|�I~�5
��e�.�!cȩi��7�����Q�J����[u寏�����R%8Gsʞ�L�_�k����nT�G����ݚ�겷g����{��C��4���t�g`�Q��~�GT�w�"���&&
�ˮ�7�|Xe%g[	�������mǥσ�?���W�z9}n�i�w�ۻ�d���P@����@�"�v:��J�jF�f���B�� Y5=v�� ��O�Frn?��R��Vz����)���ﲶI�? (������tp�0�������yy,�P Vg�mx��z��x0d�iV�I�/.�c�)5!�1( G=X���1l��}�4���T׸Cҷ����� -�b��1�ץ�D��uc���(r�=SW�*B(q���l����#�i��>?�� s�K�Z�I7Z��M�ϻ���5j��Om�٥{*����U�=�ڍ/��U����a��l���y��R:�CX�ФKzl��]Z��qѳN0g1T{���{�ca���@��>g���Ye$�	��Ҧ3������zL�����p`u9��?����Z%�bf��b����O�1r'�⛯.�n[7j2����L�N��w�n�x�z�X*�%}���#������_���/*)�b��:0]�4�����P�&ho��>{ ��B&�����׹�{l�VC�G��4_��S��?1KO�=��O&��vd���9�폺hRfwY���9ܝ7�`�?�MP0�|��O�3���*�!Xq�.1TPՓ�F��t�쯂V�� E7�j�
_)<�"3��r����y0\�VT�1�����7��Q��!4neh��%�"�������Z���S�f��<��tE�Í唾����*�=�w;���N2������T�wZ�;Fۄ����e��ó���(�4ժp�v�ll:.03�<��f�I����pm��M�)��R}tT�
�����K��2B�"+���X3X50��ZE��s�Zcw���'�)�k�a���6w�	p��V�.I�ȑ䭵���Kbg�|[���9">E���4KU>T�C6v �틷M�~��;a������ T��Щǌ�I��?�(�R�#eY[y+H�� �YA�5:O�t*��̻��v>��,,X�1�"��-�5$�x��ՇE?����P�ב��;W�$~zTZ��/��(pR�+2F)���|�tb$Q��(X+7��q�
gz�V@��ub�ŀw�\t�ղX��4w��4��q/�p�S0?% ��i��m���!ל�c�W�җ?���HA��[%�+1��E�6�Ey0�9�:�G�f��Aȸ�o#܍��$��:�(�2ƻI�b?`0�`Ԉ-fo¿�qah�˴�ș�k�-\�4>�������(c�ilM��5��_�d7����8�iN�����+\�Wl��j1g�ғ��+er=��i�V^��[��%�,)#̪��7���O�B^-Tb��'j��6*�E�(C��c���@�W�H;��T�����B���� �!�U2~^g�}fS�_����B�p{+��_vN�DI%sl�fO���F�H���{�T�@t�&E�s��)m�yiT$�jbyhk��x�
�0RF�a���q������]��]U��B���so�vU5��`M;��;$���?�<�(1a��I \K�_�6�X��߻�XᘷŘ����iG�!<��&ES�=Q�Va��rSh� �#��BO8{I�z��P��4T�jM$ܼb��=�(�[������Q�Ҭ��tWͨ��y���?�!H��F;_>�����aԠ����~�i6�wk��L�J�|"���d��^঻>�S@�f~�Ļ��k|)�v�
�*��H��2�:��l$P�~i�Y�e? 3��{�^r��LVeqVeN���T���XW�{�ē.�	�J>=κ����W�5	piK��ЄZ��J�V5xLt���[O"�,)DL_e_~_7����� �ge��H.���es���ؖt���y<��� |���h�oW,|�bPP
�,�����&� !0"�$�˙��l �'�~�秿2�^�R��F^ia^���'C�Պ�
MC}����Zj� �~?�����̋Q���:��t��(�ۃo���h��D<�@\>T��O��p`�e9ᓄ�����/�6xa[��ǴaG������k���z5xhz1���]��뤤k�||���T�rE���b�����@�i𗳐�m�Y`�"_��JJ�y�)�ê�l*�Ԙ㵮�^��$9�KW�R$��̲λ�k�#��S�
��%����mPd�/�@~�\�N��1ўV�5o��]���FHW��z��NF��'�ʝ�пcH����W"���qϤ~��`�y���[��P�Я��"��~��!��l�Υ(t\�P���Z�q�p��]���R��H!����g��k�v�G~: �4��F0@�D՟I}�i��g�q�w�؅(z��T,�MzC�f�c:����Dڒ���A�������d��P��"z6,��m����t��y*V��!?�����{�Bؖ�0O�%��-8���l�6�UR�����Us�D`��>�xg췩��$�q�A���	�2^�}�P� ^q<�0;�UK�/���%<^� �z �'�� erR��:�aT3J˲=�����h)�\�}�l�em�/�� $�v�P(E�/6CfԸ��"���̓z�=�?m1p������I�T��$W��O 8������b똯ͦ�����4��h��@����L;��u��]#�k��K�!�.:���86�'uls�d^D�j�lI��c�o��2�AJǎ�j�}6@���)U���s;Z�gk�V-�_�T%���4?�d��'#}aa��C68S@p�q��D��������3��%��{�QR�v�����Fo���V`9���
���2X���/���$3Zɵ���ȫ���O�Q��� Ђl?�k@���c9[o��-u��^�`�!��[�GW���ۏ\u�FXB7{�6� �zP���k�O)�ރ�4z>d���B�{�~�����6+
F��g3����h�Q�|Կ� E�Kfp�@�SSY���8�ΫF�+�0jC�Wp#� 0;�e'_��P��12f²����	�)1�����QA�k��8��Nq-�b�8�.�K솎��q.�m�+�ȇ�gA񾰈F+�w���B��8���xr(J�+Y(����3y\��0��y4�?$8Kgk}ݱ���9h* nJ����,��ŗ�5g�*^4�{���9`Rb�!��x.~�)��Ȧ�W�� �9���-U~���Z����+-G�����Ǳ�0��F:���R�L��bUV1�ƹ�`�f��o�zhs!��l�Ri�����`;`W;�P�s�+N>6���hDi�Zyg�KYJ��R�#��q�Κ+5jYW��{�.���^�����*P�f<��H��9�3ƨ�9�d������c���Q��\�2�_�t1G/i8:�0��Ж����(���di�k�GPK�����zl׸�(<a����7�K/!Pưk?¸�H�BL�w�Hd��#$��'��O��i��U��+�G�U�T�a�UnX)��N٠ބ/}?�s�[�=EN�"w�áηY�Z�>�A���ߛ#*DZ�d`���w���:ji����$��{�W lG���r��w��m�1��l>�i�>E`m��K���ֶ��1�@�^z������k����%ӏ�L��
�ōL
���[��I7qPGR>cݚ�j�ת&�-b{��=���)8���]���6�6�R�f��Ů2�{�]������	�%}9��L��x6�wB����G:��i&�#��#9��z^wYjϕ{TJjH:�u�˿o.��L�?R��CĜ�_��+�%93t�e	�j�(��Z��]i�A��[�r����ă�>t$��S�:z��-W�62$>'�- ��[L�yec�"-�zN���S:�7�~w���$�/��6B����n}�H�5�@����>X�4=��P�n��^]r���0{��^��>�e\�,�ndCn����㼗���B���\TX�2��A��
ՙ�����S��{�1��~�;SUi���[�Y[���@/n��r�4% i�'k�:�)�
�SJ������A�:j��� %!Nx��Y�W ��cUI��e�Cz�?��`������+�����e_�G���.����)�}{��k!����?f���*6�:��
����G�nI�1S������N��+�b��&�/����ѻP,��n�:ƀY�E��*Z�k��2���uC-Zӈ��i��d����f7�� 9[�F��)�O��!���'Pû��.Ib]݄$i
Q-q�SUp����-��>�����ѕ0)�aƓ��3��o��Y�S28�VyXҫ�o�$'��;
|�n��Z�O��U?>@D1�ͱ;wD�Cucݠ.�؏�*��Ejj&�KJӻ��ڜ�Bף�]V�9��2�`�ج�o8Ys>�X���snmgY�����
]?paěu�0^PA��=�	��g�L�tf�~�y�v9��p�3u����3�-�<
�W���֎9�֨�`�(`6�3Ywk.��j;w�-�d�ɦ!1[-���d,ݩ��B�|���&�Fe��+N����/[?l���DQM9|�2����;��d7D �k�N��n�EQͯ���8�3�#�VE[��j����D&F�{+���~��+V��3L�۪��3i����</Zʺ.*�WQ)�Of��sa�d�$��9#Ԫ��W-��je�q����Մ&���8�ׄ/	6����y���^b=F��hj; ʶ�$�h��wi�y�q}y�]�^u�n@닎S����r/.v���\�(3V��Y`E����_���4������(øE��p$����t@��W3��e��+��<�\$���Qn��uy�,Y �4)E�:�'�T�w�M�N���k��h�V�H�)��b����PDU.�^RO�gVT�Ի�cUd��=g�*]��Z���z��U��O�-s'g�*iVTL�l@��gj�p0r.ENS/�+͵9_;��yq��D��M�B�T\E9�F���*4}�髌kH�w�ƙ��K�9����̵�$�T��J��a���� k�����A�g@a�1�X�M0��y`��fVtR���� ��k`U.|=	���vm��n�������I��g�CM���S���J��W\8�'/�k1z^�'���aQO�YV1K�0u�\q���o�|��*���Ge*Q���`����ƳC�8�AS� ��^��|��ga%2�n��x�^���YmMmѢ���ژ^�RJ�`�����5���Or۪�$�
��6���=�=+{ezHڎ�eȣ<�ǣ�m��jds�ՠK2_�A�wC�;�_��{�f:�͔����m�2��عs~�}�L��1p��}�@��0NE�N������8�-[F�>�$�b�?����c��r!2��$)�C�<{���\���7��^U�/�jv>.+�M�Z˟؇J�*�"�_���x����f����9�ry��wgp�ی~�k�Vh�i`�� �C^2��D.y���F:,�&�O�W@H�}H0
[V+�e�ΣH��B��(Z��:�]�;R�u�f!U�R�P���9�B���%T���ç~��CB��n�Ȱ��I0Ơ������ԥ�A|yc��T�ׯ ���E�O
?D�i����$����@�����+%l�|x��SN���y}~J�=�L�]��*�LQ䆃#�����б�l�y�^Ī w
U pRz(��3R5R^�#F�������G�01C�銡�x����N#[;�bؒ��:("9�8�ܰ}�"E�U��m�!��f�8�r*JR^�@"�{})úǇT��u[��^�w1�$����e�虀��Y�&bTy"`q���E�R�7�_4�9����b��7��u$��ؕe}�{���5k*S�;�җ�&��akڜ�S��Ur�	�B�P�������F
r�*�@kH1	��� ^��z�g���C�<���b&���2�}���o$斿��:��
*�R7���Vf���=�!����z�����lLKM�?Y�����{��O�)�z�s��oͷ�䓵2o�/��z��hk�ؾ��<���R&�mO�Ȋ*����� ���E����*�%~��JoV���s1|J�z��Ľ����֮6(Y�÷��U%�^G��'`�y�R[��bo�9�л�t4[�Y��%�9vTE�[v�|�������^�ܥ��h����k��)E/�����!���j���WJ�UR��M�t�]6 b�:�궯��! *�Wn\A_;�*9�D�f��No�{�įz���s1t`��#�l��}K��H�O,à�.
��������Z�ȇ{�R��I�B�9�Nq�?�R~D$K�Ip�h4���%���0@���9h0�[�U�?���bKjR���f}��5���>@D?ـ�~J�=�ǹ|�J-�5u���gC��R�h.`GrH�U�pG��@3ĵ՜�Za:��tS]�/&6g4��wJ�D������R$[Z�VN�k|GNL���iZ �)zߗ#��	\A�XH�$j�4ݘh?Uy�vG��YU��� W��4���`ض��2ym� hրc?�gb�:8�:��~<�#�j	���M1�	�az�7RN�1&�X>'ّ(�Γ5����6�����)-��ė%g���*�X8��ʋ�.VS㥟��,�}�H�%��������,����X6���y��r�Yu�ER��W���l!G���r��%n�o�l�>���OQƜo���Od���>���u�Wϫ�?���I�@��;�"N]��E�a{5�䇘-�9֯�ov\���K��7�9���VԒF�@���r?i(֠�֕��߱0��p/�w@ȇdq��D͎�Rq��}q��;��М:w˗�M���U���w&���z\��G�n���Z�f/o��3��f:I%zs��YQ|�5�B�1���ŮW�6G]�M�j���}7J@��U�:*	=ds	����ǐJ�J��Ƥ������HM��s�eL"㓍�f ����5�u]-��t��n�f��ғ=@�컞;J4��I���F<_F�ɺ[��A��oM�MR�D )�X�O"�]�A/z,�D��"���Zm�$}��Dϓ#��+�4v�d᭨����%�,���֐;Ƌ>�,{���?����r<�[,�N�*���Ȏ{l;���ڮ_Zn,�@�H`����-�U?�>"=h�H��.��Iq�0Inn�h�a��O/��^RA����ܶ�$ځy�	�pN�D�U-H����; �C��ȜR=Ā����m�{"<�y�d�w5G��Q�].�Ѷ�wň%��2Zގ:3�A���{�:��/t�S����Cq�j}�>��c�Jז,����ݵ\�l$h�R��;�=�é����4�R��ܥ����q?M#K�� +�ā
�}
�|�!�լtA�A�ȳ��.�5M�+k�6l�g)�X(R�]��9W��ɒ�3�z�F��������]����.e��˳��Buۧ�)$Y(�Q�|�Ea|٢���=�\]�����,v��F��U�Um��с��l���$��d���ǆN�}J����:J]���h�xrֵTT��@���6�^T�cc���������È���~k	dL���.� �`��Ɵ�a���`X@x^t�@��Æ焭�.��[8<��f���+�;K���L�ے�Ҵ���`L�L��tNp:1�Bz�8���G�!�Ž!=B�9ũ&��3�� �\�D�2� �/�FY�i�0�Gb�Ҡ5�����F9���ۀ��C�'�eb�;فn��ޖ�*?�*���`�Qu���Y�_����]�%�R��J��g@��?�=��-��}�2u����S�R�;蔄JMa�!�Ͽ���si��]�鬟����L+�B_O~,r�6��y9�V�?��K�2R���]�kk*cH��8L��h�ٗ�3fG,nM�C)�G�RYY��C��_e|<���*\�`���E\�OG���J����9OA$E�\x';fx �e�ۡ����6�V����e��*ٚ$Eg����޹�X�.���� <���2T���y��r!.k�}&Qԉ��۽�����r�����n�^���*�x�L�y���C��f߬�����@��E�5�����-�?�۬;����Ȱ���.��I2� uҡxW���lm?��G����~�GZN���3p�7��wO����(�F�t�`ĸ#��1:�c�zŒ���[�IY����[��dZۼ����čP�i��R��;�G����t���oh�TS����`Hұ�=��.���us�"��`�MQf\0����j�V~_����'ՌHp��Mv�3V$�a�K5	ں��/�MF���9a��lh��%�F�
�D�]��[f�i��,p7�pJh�˗�S+J���o�Z��g��N������ߖM+ubc�ɕGc�(r���D7��WV�,v|f
/�Rt�r����V�З4}�܁\ a��� �jЊ#e+=c
��,Q �Ak�*��� vv$�1ǎ�������vS���;��I��]w�Q�r :6=�P>����˄T�t�`��Yx��a`��`8�묚%�ܶ�2à}�cm<\���JaKFt�#3m^zqf/��ԁ8O!�z���B�`	��Dh�����cE	� o��>&D���E/�`�k�;R�qR�h>'�M��>_'���Q�4_].y�{���� э-�^k3�
�	�����ݞ�p^�y�$<zD�?�W�.���Xh�6��j`�� �  �e^��}���|�h��7�s��ཻ9,��`FR`A�97�3&�9g)�H�F.4?~rP�XEj�O�C�Әo.�t(?c��v1B����&��^�r�>� ��bx����r�|��|1�Q_�xk����"���#$���H� 6��<�޺���j��{�x��@��'&��ڨ�b�J�S�p�e/ۍ�Ϻ�<�*���|^���U������;��&�n{T)�G�"�X���YT�7⹜�d �XNRe����	`&�F�M��o��b������|8�ӧ_r���,�Nx&~�d.��$�9�}NQ�_�S�/z{�W9"�	���L� �?�2�����<%��_�a5_��{���DV>�[��v���ҤBwG�̶W[�aH�/2O@V�q��{ڡ�f-�����������9��� ��X��v�P*��E�Cw�:�Z�:o&[&���d��k���bKM�o@��������M\��K�Ss��v�	n��~Ҭn�1+% :Y6ZφK�ZKſ��4R[����� �/����z2˄��� ��4{��]�m����)µ�*�A��w�O�+���I߄ ���[1WV%|���#�	ؠ`�ђ[���� h����H2œ�擽�d�S����d/��v�;#�d�g߉��r�iv��W>�c��py�R#���Z
[�4�������ڱ��53��������7�-- ��&��V�`��Y�4�G����A��HS�ZL���KVةP�r��3N��,�^��I�z�#��r��wA*n��g[��s�?�k<���g�t���d�U��&�Y�p5��2����$P���[���"@��*3����[��O���Ikl]��B�-�w�<��!DB�-�9��:�Ur���HHYþF%��Ps�b�C�uj``g���:����1��?3j�Ji��B�,:��ns&�&���֜�I����z�DX�8��z��{ѥ֝��IP�>��$���B�'��lu�uQ+���:|(�	c7-���2#P�2�[�+�c4���q�&�Pb�;����"R}�2Ĉ�[%�gٴ)���|�Ntbp[�;����(�G*z���j�޾�}G\�0^�XÑ��v���w�/�c�Mu��a�
�}g9�PTOK؀~��5����><e��y�$�
��4��<�
:�^���	=�zy:9��f��^��*};��w��=�z����ay�ۊ(b'J�5��ĵ�{��͖3��(����kk�̹=���74��[�DM�GG�����p�F���L�Q�:|R�H�?�ZXL��n�lH&�������HS>TMF��g*p��E��F�c�ֻ���E$)�X�%:8��|�Y�CjS*�z��b%"`����_B�!=���)iD�Q�Ś�ܝ���23����e:P������������4��>��/�La��C�����I(��2$%�R�<@f�	�,C��7�%?�=5Z�����?�K�!��@)��`�(Ai�����L)vkF�xD��Q?�[��#[%��4VU��B*���x�;Z,�R�T�G��f�m�(�Z�&L�4v�n�9/=v�pa 4u/�l�w�r�J38
ms�U�W����@���(�88=����G^�4��?�/BA'zȆ>�{��䠒(�J�C�ҞX�D���vM�A
��J裻���zh��7�,U	
�O�!t�?#I�	-��0�������G���r� o��䏒=6�x��i3�۸��O�A]����b̌�Rx&�˨` viy�=��JE�>��<($�ǐ5pY��N�K/٬F��`M#��ۓ'�*�y��t�!�K� }�FYа�<��ɶ;b T�vU*�؜�D����v�C������p�e�@,�܆Υ$���̎?�a�hIK6��&h[�)�L)�Xոg�Ω��T�n+͗��O�����/ ����d�a�K@��u-?���(�,	��@FQ��mU*��{ix�Q�'�W�n�Q<�y�ͪ��e�\NC����,�He-`��R��Kt�<�Վ�f�e�+����B`G9g��L��S�Ri-!D6&�*�������xX�Qf�����5�NX�3n��,��)N�ſl%�	��y��WB�T%L��Cq���zm7������o�Mr��@�Eb�o�;Q�`x��P͟fW��]Q��=!㾔N�1 ^e㛈����e1�#,�"{��8�D�g��%�&���9Q-%k�\m�̗�e�4s�����׫
�#��s3�ڤ8��M�=��(rB剎3��W�t��r�ȣ�͘�n$���毮�Ї#���G;�#�.����c��c̤�
Mע��?HRѦ]d��f&�ǧ�v�iD�R��J~xTn�8�>��2qhp�Ƚk�͍�]���~����D^0�����&��)wV��R@�1�^f�k[��[����g��q�e�����z������kq�%�����?wrC�FaQ-�9�fJ���v�AuN՞1�x_W��H��b�����,�eUp-~��g����F��tDK��/ZNňU����3�?,�c�O�jw/!Ue����-�w��Z[)Cx��� ofن!$�"M��������j�my��ѯ���]6�O��M�H�e��(��x�k��������(� ߈�oJmj_��o������_�T�og)�O��U!��*j�>-m�o~�!ImIӦ��V�e��c����5�咙����k*�L�2��)���*�8 ��e���T��{SEeO������ag�Ǘ��"Dk��#�]������!a"�$4T�/�&k���D1��5ۿ���b~$�zQL����`�ޱ�����˥����+Z6a�t,���$�� �O����N:�uD�?'�y-�3I>� s��"���.3��ڀ�L��//͑�����ij�7/��M�1l�6�K���\�=�[\����F��467�*
��z� t���cZT|u>�c�CGϻ�$_ޠ�/O���^62F�o'z|z������M��g[��|�A�H���*���L��r6���EH�F=��o�rq�nfU�XP�F��XT.{%fr�D`�JatL�%d���%�ݻ¢}�U���5��|Je����"�۲3�j��O����fZ����̨�D�{e>��s��]j�B�yK�U���-ⶰ�~)y����ݢ:;�H��/��S:�^������K{�}l�3����zy(|N�d�5k���[�OVϛ�����K]�G��zG9�@��i\�I<qr�5pA3�R������F�����������6{W�X,��za_S?��x�Pz����V�gb}�T�p�2�����{r�H��7��l��FF�"/V� A�]��l�=�������W��fHG2+0���lq�O<e��s���&R���!F܊�a�r�.&�%%�I�����ɃX��q��~���Dw�]�ʀ������lca�6.0"��Uo
��^�&�'�������Q61�J�\E�Ʈ������x�:Z5��I���pjAͭ�4����#�⼻f{��å�l��f�0�`a�����
 �m�u&�]1���P�I��
�����{W�e�քS��O6�o~eh��UH�m����L,i��DN��.j���VTF��nk�Sڿb�}U���	�\%W��䣍=��Dz��e	d6�NǛD�EA��}�q/��7;nV�;������W�z�f����Z���̖3#_��T}hu�fcojYUl=-��n�v�]����R0�ֲ�{�!����&���4�\.{/^�kz�b��F.�C�}���D���kE�ǒ���]`��e��}LW�)��/��6��9��nl�Y�ɀ��"��D`��gJ$^"��z��n�❤g��~/���q��v�%����5[�k�){[�T�U�h�z0ʟvh#�{}g��=���("P��4�܇y�
!��� �P�RP�8�
ǔq&o&6~�
|c�{_gO��sP<��a�&Dj.��A�����d6Y�Z�����CA�W��V�{F����̑Rv`��͟��ܻ�=:��R�=��: ڷp=jJ��HnY,�g㪜bܻ`�Eq0E��`��k���E����%d#�AГF�ծ��ߵ��v���,F���;\=�e<1��l�!��u3V�T�e�R��ǯb_[�:��]��[���S��
Ցg�����������$:�c2�d�]$�7�:��:d�VE���9t�쁍K��YK+ͩ_�e�N&\:��_��U�xU_#�?��k:��ў�+|��N�H<���O�FV��;Э��2���!�J5v����d��#"T�N�ϼ���fKb�� �>/���=�0�5�+�a���|�f��$5:zʺ*�@V�0��=߹����4�<���i#��sa\��s�������U��z��*��p3�J��(*��X�n�I���bC/��^��\���Ib�"�~H� ޮzn��=�-����\����ރs2���!��+�Q"�;�$Ŗ��x�����g��V�A�C��3��B�M�
��I���{�4V���R�wB0a���}m��I����>�qp��0$R5�t�ɗQ�MnB�ۢO�|��j�<�=��ը�t���\��Dц��b��p�Ov�۷d��_�T�	V�U�yL���(�����+2Tàb�&���9�<3vVi��e�Aq=TK����ۘV$6��+#ߴ��k5�]g
a���8w~��,3�&L�	�,A�+j"7�K��z`��x72�а�#�m�����:���~@�]Ѝ/?�x%q/P�w�+�8�?�k����L��'�Xs�a����R��02��L��<��ӹ1ڗ�_o��.���V��E7hRFc���cEPEY#�(F�ɘG6GQ�u黎�?�V�n���T��=3�ë��;*�Y[��I�s`��_�SĪu�?e��������۩V�s�9���F�i�p|���"8ӷ2ӭP�N���O����Ido*�t��E��L���\�6����4WW�͑{��BF3�K��پ����4=*\*�
:(B�N�ss�C���
�1K�f�*��KKF�0�_��%eau����@������b$�R�c$��z'���e+�c�����9K|lynV��#��iG����-�oPF�T��)?�c�w�i�3���YE�"0�&�(t4:6_/9�DZ�J�����fSU���^p1�0M���O����z8���>����������QTЛ61`�b����Ъ���'3J�t��Ԗ��,2���p`�X�#4N�_^�r
m��A&6Y���K��Ц[kk{]B�����g��^u��YY�.��[�%�k5�B����7<�����f�O�{��'[;��nl�}wY�M�� �$Q&r0�D"kN�C�ZϛF�I�2�at�8�l��n��&�dH��49���m15t�~���9_�:�%;��/�@���'-�٥���A:uV�V�j�5Qd�C���nݾ�9�$�Y�S`�ap���21�"i�z_x�����0j�δ�X�ȴ��SP��;�>�M>�5�`v���6��L1�<��0�H%&�9|g!�F��&��h�����d�WC@��" ���b^Xg<�ޭ��E��Lބj|Z2�I|cXǟ��*`d�[����cG_�8��>��g��E�y�d ��$Q�`6��^�H���7Km�x�C^è�{����ٵ�S�~�XF�rIX��d�/	j&���撾1����%�W�J�G`Ȋ�����k,�� }�;mj��@gG�`���8cѾe5�ekj�F���Ȃ��Ix�����)�$��L��t'����~n�>�RU�#�M?)��yȵr�4�m�x��e���k5��OSa�͢��b���Rբp�ee�����o������*��7hM�� �l{�����m��)��9fh8R�W	�?��i����<`���5�P�7�C	379Czv�R�) ��~�&ſ2]t6j�e������X�) F	�ԛp��	�X�~����~�A�B
�]�vD�X�l�ST�ݟ"3�k)[?��+�}�eՊ7v�A��6w6x^d�����8�/ϱ�:�W�74���7�Ȩ��\+Th��"��-t�����4�������AŸ�y>����Ez�_g��E�jH;����ɶh�����3i��3uL�{�g�7'�S���d�yOv.Ȁd�������v�#�WօΖI�����ds��jlk�{�F�����J5��V�#�{�*jR��_���q���q{���S3~�h�枾��W��H�l��(rP�| �n-	oY4{�4�-3�q�y�)I�z�٧ܘ���|L�ZMw�V>X��l�m`���K�-�#�e6��9����$�\9堕MgDz1���{J�dXz�����X�I���]�!s~�@��as@XNW �e�w.��Y$0�ɰma!�$k����� ���z�f(ʔ�u���S�L{k�f�#r?F��+x<�'J>�8%	�ʱ���$	pS�&Qϛ���:AVP��^�PpP���(����)ezn�@��8D�Ա�N�R��y-���~���<Κk��;��`���VR��J�ꫪ2��M��@�nb�]9��j.�|��d�M��Te����i�iSc�-%��8=���ӋԻ��� �l�ͭHw`�li2M��A=�1T�ldr�b�6�l>�դ���W�΂����~��Cǻ�1�=E��Y���=��R�X=�(��Du\Ó�7���!��W=���>U4;h��({�"�B�${+�(�:�8E�qfH�G�p��R��.q'�
�?�����LO��j�@h��O}�bf�U�t;�N+�'�I���5���7v6hq�>��蒘s�3]�R�LT����M���n����$) ��-�՟?��r<yLL`�{[�!��%���6
Ѷ��TZ&�/���)!2ÿA�+�FU�|H:�D�m��ʗ����PJ�7���pè�4k�#�R�����G��;\�Ifar�r F4K(�n��g3'��E��-v����/�=}��cY�b[�i��I��@�S�r���ȐG᡻3@�z�B��� �9$����f�s���w}�(X�Ad-.�
�?�}�x������4�E�U�/Ь~�Q����S*5��s����Z�m?�l�9��75O�ڴ5ߠ�i�$�ڳ%:ל�Թ��ܼ�TZ�-2�;Q��*���Ū9��?b����9|��E�9���V�Aړ�u��\	�Y��h!p�h1e������сLye�HRDBy����ж��NdU3��i:��i���$���;GG�qVNO%%�2�z2�ӳ�%��B4|���zfY�j&g$������}�x��u�p�>��7el4s|]���-T-_	T���P��&-G�?~��`��i�m��Z2!�]G)���KF.�@u���K�Z�H|_��‾��;���C���Y	����*�>y��(�%��{�x�}�����;�*ղ��!�аZ��=60��!��NtE�)f���K5m�iऎw;��!Xj����R�)��M�oj�GK:s��o�XXy��¹��F��,�0W���d@3�a:�9�������� ������n�ԁ�`"��E߹|?�>��Z�4�Ӳ�����!�����ɧ���u�@��ԍ�F34NY�ú���������	�|^�}1����H҉7�d�?�Ӗ�*~�A�� 3^VX�*kJ`��x�i+��Q��Q�����_�ܵ�Αx�'睳���#*��I�l�m�oڟD�o���p*A:�-e���5dtEa'�1R�;P���y����}��/��˿)s�d���yPV(�uJ/���ii�UzI���h�e���v���*�*��+����l�?
�Qk���x4�	|�{	J>˾S}�Z���i�ŗ��*�j��o2*t|-v����9ܝgC⵼��\9]��~���HWО��Y�`�b������P{�D'd��H>��p�b�Z�xGccY��R�v��~r���l��VT�ڀ���J�H���S��F1"��,"i�׼[(����@�@�}�9l4������]��t�ϋ��(5]�����º� 1���� h��������[BK�����b��VJCo��m�X�~�@n���T�*�s|�F�7��_KK;�a��n�~��aŘ�ѹ�*�Ĺ�:�65s�)'g�c�ME����O��;��K}�D4�U��]��S���<���쪧��Gz7�K@7�:K�-]�@��w�i��,j��%6L	�H���Epr>-BvQ�G����6�T�u��U���b��Q�~�U��O(]
�uɁ�k���X��\�$������s&7V)Of��ņ�I���\i=�	�1D�Ò�sZ�ؾ�i��m�7@C��2c�S;���b�hN��GHn�����r"�*���9[+ץϽU��4ʜ�TBv�2F��������Zԃ&k������9���c�"m&s������9�O����uo=�o�-�����eA\���+�(�4����h����l� ������~{d/�E1\[Ŷ��H�Si���?*4�${�l�V<�@���#�o�w�E���>�Q�yۇU���i���j��b�y_�o׮`�Oy6n� f��6�h�����;�,@�ün�oN�bZ&f �ʈȢ�/�Gv��s��db�Ó�T>;\yzQ���s���x!c���Rխ����u�=�ѥ��� ��E��8t�x��VU3Ԡ�o��)���7�͗��2@�s�%�^�6r�hW�>}=Ӌ��k��΂�6��(I٭N�s���CM���;\?'Nvم����D�,�/5|P��U큄�֐��BT��� �[C2��9?�f����!>@z21�U'P~^���h�՚��J#K&��;�4*|��΋�s8҅c�|	�\MRoY9&������'�u!J�N�OzH��b)9`���D��l?ɿo�� KB�n?��.V3���VK�!�O&��RA��l�0�;D��Sj�rz��9oZ�9��R����<E��7����1)���xNշ�ՂU�YŃ�+���9{���\+I�/���i{��۴� ����A�?��L��'�4��ySX'���/m������y�S���(��;pٯą_P�6A�6��JLq��G��\&���sd�ݬ����i{}������Q�\4:Tª�A��H~ɐ'V:q�d\���P���^^�Ϲ_��p�~վ�eR���a��(aA�M�4Q�NV�ۈç�nb�,i�}�`�6L��ؾ<u�-EH���G�g��JU�Hd�NR������Fs��ߘJ��?��#C���2�!��`!����ש>���_�`�����)���@���kಯ�ҝ/�#�m=�*B��/qSΪ���8�� K���[o߇�v�Q��`�ʉ4��~�
vA��X3�r�o	�ڊWM� =�d�ߩ���u��ty����t^Z�e��
{Ggڑx�?ͽu#HQ�r�Z��يE�m�͐0D���
2�O{q���ڭ���x�b����	��p�����YM��̓w�{��������9'�������<�ο��᷺݀�W�%�U��an����\��ֿ�B��=Y�h-����o�����fi���TK�j���c���4C������iS��&�q�`[0H�e����{����'�u��IZ�S�h�0�8#� $�]�W)�La5�8��kG�e��b׀�H�6=��������e!7�=�wS�wEG�z����s����i�>�������#�����.F4�8�xha�5ȏ�6�f���j��S����k�����tܰ	kZ�S���n|��b��o��v! ��"�x�!��O�v 5����?%	��!=����Pg9������:�D��d�He�� ���#�ٗ��{2�#�"��<�B'��qV�?A�������Ҝ�3ԏ�/-R�`:�����
�=)�U�2����C�.����,X���XM�zj03��Ҳ�	� � ޒ�GE�na���1���h��h�/o�I5���
�)���W�!�/����6y���>�M���;�fD������R�m1U�
9=7��~��ʶ�S!�HT���gdq���pBێ>6P�t�_%FD�Y����VD������/�/� �����a���p�p������&�EfX�)>�R�^x\x'(7Ad�5u9V��=���tӰr�L��M��{��?0�ڵ��d���a9��^��ԁ�´��3)�!�&Q��<&ˊ�S�\$����Z��*�l���]?���8��43��ҾAtpi�;�]U��9!����~��݆��~ϮZ�\��vG�0-�����{\,3&�C(���"$�sS�oc�xgkA�3?7���ʬ�i��v��CFo_L���h�s�b�C��y�+*s��/I4I�׺��cP�4?��K�yhZ<j�����.�R�\B�J�*��P��v�m�G����I S�+��#M�<��"����>��3L��W��-}�%#�rF*�b�G���نd����g�.&�I�v�_!�_s+�K΃��c7,<�tN�V��!pUr�;�`my��Vq|���n�Y+�P'���9&�+��;�9�Sh��ITd�d�7Жc�RTo����?�CX���^-�_E)���A�rWb�.��j`��r�ֆO=��M�ӱ�EO'�A)T����ւ-g�w�y{�%z��Un������k0U'�p��s�dFg�)�����O�+1:��2	�p8-�h��Ư�1*@��މ�s������y����i��_��Mcخ��dh'�1�H�pvV��Y�ꦔn�sS$օ����w}�Y�;�}7bX�f���*��*d�N��q`1/ȷ�/%�4��XQ.�U)Ƅ'6�E����0�������n;�`^�.�T��Q�?�#pM�v�n�V�+��چ����$s����7��.��O�]�M�y�dhً�>0EF��A�M�}Wd�g���n�To���;���+fC�|F}�-
I�����������;��EBIB�/���Ќ��?NF�(z��<t��������~[~�=��~r6k�z��t���Ņ�:Ƿ�j��<��>����D�-���t�:D�3L3�|��/��r������7��j_�7�gqU�ћ�'[�O���P�@�Mp�"��S����W�X��0�)��°$k�Nn^�o�N�)����`i}5!���t�³z^uǝ��cVTg�~l]�	��6ű������I+�U�����Z[w�H��A����2��,E�%��B��riy9�q�� 40�ܱē�[#�8	������f�jp�Ә��â�~�L�(� e�tKKm�:1ɦG�>��}�sI���z��V�*W.~P��%|�<<~��)$�4�F/?m��R���iܠ�Q���:OI�2ft�I����_��[�G�w^�Qje�?ԓ��|
6��\� e��������X5� ��#��U�u'T&W�4����g�$%�����~��"�뼧���-�H�e&���tH�wf[O,�y�6*WZl�!y���?b��!�c�p��7�IQ�f/P�L?�Z3�0�Q�&h�M�l#a
���f1L��e�(�
����hvq�0�c�#Xͽ�̺}$�{ɎT�+'�(N�q����'睂?�=�0{xP�R��ܮN5ڂ΄�Ӣ�oN�zfVS�6Ȩ7�P���#b����ߐ�$-^�9T�V�ꠉ�N<@�k'g����:4(=�� a�+8�9��v j"V�Y�3�)k��ϙ�O���:e�)=;nVA�Q�9V�d�Hjeue��/�=�P����n�|]�0lO�Q�1(�*t��w��6A5�B�I;S�Q�F����We��E7I���G�CNq�#�U	5���*Q�h!�9e�~�C�h[o~�Q�vL{�`(Dr��8��O�w{��m8'��Z.�<�H���������Y�S�[����V��x�co��$|���o�>?��%�[�Z$S]�?�;��: ��
%2����h��"�Ӕd̤�?P��VP�4�=!j�n�(�e�I�YIa��Jl��n�c:���L�0�_"�� /��nAv�0t�R�r�.i��[�T:�yP�$<�F&�-�v5�L�Y�W:G�o?�1�ce?�{d�|�c@�C�h�_�Ǟ��#�쵰F��3֮�Q�����ČJQ�?��ð���'w�O���os#>�WN��GW"p%c(@7���'G�KtD&����'�ɒ�\�ءU��&��{As���mk��l�*A����|�Hd{y�o���!�_���;w�=�ݙ9�6 j��&ˉ+�ٝ��ESp,�Wͦ��;RȈt'%��zF35�3Q��.�Z <��I!%0t�Q���F�+����T��'I�����z�L���sPn��90��ݜӌ�}.���-Ŵ��_�j�е�Dz���c��R�^A�.ͧ���sX1��\��O}^�qc�T��j�"I�ճ։��Y.�{�o-1�M��;�l��F1��43�ʅ�6N�
��x�<uu��E ����q08�*�������B����fa�&��3�$��,�f��ȫ]�Gg�"�w������ldX�.�/�]��r�����M�p�Y��iym��abQ7�u�|������i=��ME1�q��뒏�yW�Kڝ��ϡmm���:rQj F�3�V�z��ƕl��$����_AzV�� ��"�v�����3��t�1��������kX�Gč�A|,#3d{��e�{���+�ڭ!U9��"Ѝ��1�%
H�K,���$���f�!xMni'�p��!����Ua�k�����H5W�q��
�`!I+����?�]��ۆ�ȡl�(6�WQc�Qi*�7M�[�_d��9b@��O��/�
��I��y�9t�9�I�z�*�_
Ҿ_V�r�ȕp���o{!�0�pr|�L�i��i>��Gx��xI�ga�����e4�ĺ}{���e�	��L�C��|QJ�=�\<@O-ӳT����i��E�Zy�o<��!j��WT0'1����N�S2.cFG`�����r�?ׇ~��o��{,���R�z?�9�g�٣5/�5-����P�~�3n��l�xi�
�X�j
�4�m�����M�8ZcHc)�A�װCI�:TJ�u�p�^R�{q�	PM��T�����Z�InJ�L�U�Ȫ n��Z5�̽&����V��&f�m6���g�3�8(���D�'�>���M���y����"�����H�+�؊'Y���N���׻3894 �=S���޸�����=ײ�mLc'�n&�F�2�q9m�F6�3�C�����k6H%������ǁ���J��~��Q�]B�a��5����[AR��M{��Æ�Y&>��v����&�S;���q$b���y��q9�E������2 %@��W�,l��p.�L��2=��&7�*$wL�B�ϼ�烼V����<!���lN��RA���t�
Wy3�ɸ�X���Z�B]�@Hɜ��8sِ��(jn��O�����6�Ar���@�HD��>Ϣ�����vH��Buf�Ol�*+�J�XUO"@�,����U�rC.��/�@X��+6Un���M�]M����Q%��+���;�1�L�8����>Z�t\&��;�! �ƭuC��AmR�A��	���[���o�,��Y:&(>��뚤�3����!\��Pv��z����g�
�3��6a�k�<X_�L)�U���;�J?(v,�Ï�3�^��ܢ&a_����v������ �.A�bK
���f��@a6(L(�؞�n�,��K���3��K�n��k�e��`��G�n�*�1�BR�|%}�{Ԩ����4*�G+��E&��7R�k�[��HC^L��-Hej��)�;i��m��]gT�s�,��#�����Ek���/�e��|H��ͅ��Y�<�73��
"��
m�GL'X����]��hp���
Y��n���Z`s���8�Δ��H��:j���_KyU��'��pӠ�yMsT�h0��jp��0�c��t-��`L���iF+>�r��V��RE#ꨮ�:k����_'N�@�wI�����M��z��]��<�̔������	E��;�|���J��i��	�m�#�/�5�#�f�`���1����,�{k����~�ns����5QY}-J�|D`8+�{і@@��8%�B�V�-9�Qj��m�tm��N�a�,a�2W�v~�Ga��PtG&��T�O4�S�X����LVR�z�5(��1$甬��q�ft
lu}��ܠ��]m�)�i�����{B8��3ޖN8�^P%�}�L׶�t/�^2I<?�pLpT��B�-�%rh����ߺ���v����L�����]�XӪ,o%�Q�Z�4x�}�i���
0'^պEb����^����/+��h�ӅE��sc7s�6jWǆ����5�҅I켥C?���������}0NǨc��*��ҕ�3�2�ra,�>����C�(�-�6�����nBSS"�7�����^)Lg:t��Td�K��o����d��Z�Lu������@˨c�0�r�l��}QIFB�&�Β��b���G��S���`�9���e�.pB�Y!?(��bkߥ�8�����z�(�����3{}���i��ԋ����T퍎�\��[��.���ܢ��ыjo�S�N���U\�׆3~?=	��0B) �G��;���S�rk�?lR��A�Lr(&�S�֖h�&��&9ގ�~;Y����U�,`���mB��L(t�z�Ԁn��瀂�y����/e{��i='�_|�R�ŇԣS���1h
�x�Aq?9����HS�,��E��_3��^U�� 3TY�mՂJ]d��	02K�K�R�O=���&<	K��}�c"Ƶ�(�06����f��&m�tL �j����H�ܧ��ξ�i�m1�t@0�E�cI����D�]�5��Y � �� �W,+�r�lmb�F�.G��ͣ���!K�3-����Z_���z�M1 �.�;8@*0?eXpu�U��N?Yϙ�}'ewD����@��vQ�Y�)v87���b؆��Mv:u2�}�T�<t���+�x��M#6�&\�Z��|;sq�w}�D\ZvX�9�X�5��H��R�
ʏ�����r�!:�v釶��^grOk*��%-��n �S���H�t="��jps�ɱ��L1g�4h��[�W�S�i�%������Q}N@e���H4��]DÇ������W�ӝA���k��L�j�A�$O�`.�}�u�̍Q��(���X^�$bԿ��T�\�g ���,7����8%ˑB��i����JID� �sEd��j֜��d\8��޾�&�`��Q2W?h",!Po� P�$6Q���:8���?H�nA�4�3�ǌ��r��Z���ޥ�6o��M�a�
\WR�d���'�%�6��-^�O��m7FO�m�:�흥)<�{$4�����0����mO�5����M�]5�����"s+¹���̼�%�`h�2:>a���ZwG�gNs5�Q�����2��j!�_`*<u#���M{+^0c	��#њ�\��/�l�G�D�w�E? �����飧|�t���ȭ��Qz܈wxU/�tW|���U�jA�&\�j�|��"7��|�s5AjFDMq3 �	@~���s���:��
8B�(��Y^��2���@;+�*�X庖jo"Ƥ� �Z`h�!���ݭ޷u�'��<F!�̋i�JO��4{I\v�5+h7��KP'.|)�;t���3�Jڰ�֍24=iˏ��v���׈a3`"�kɞ��93�w|�x�o8d�ob��;�-s�2���a�q���
>���l�I��S{yC�^}�B���4G	G��}|�}tǸaR��@{��#�=k��	���j����`�t���*EN*68Y�R�A:.tDK ��@j���-3���MU%��ک��U2Ԕ�0�6�ַ~=���* 7����n�c��*'��W2�r�P�P H�a�'��aT)�J��2u�v'����{n\d�R��=	SR���h��2=�dɔå4�SCt��o^�+/i�[�u� �8$����jW�j�g��ڄ�no?��-�_}k�ѡ��:�~���?{��.�U��((�l�m�#�jd�eȾ"�"G외�ұ�s��o绾q��O���G؆�u1yO���S$,$�9q�! %�P�tEv���J�sϾ�S�����^}YuA�l�V�e!9{����*�*\;|M���G �r��h�|� �&�X���(mT������,J+���vg�cCvI HK����ٰ����2[�ݐ�QBD���<���hE���=���r;��#sTǬ�-�o���auSG�LL����L_���ed��An!/>o��)�0�g�.g�4�o3q\��K������)�,M]x	}���Y��	8:�*܋+�d���"6>�f��؎;O0�x�G�? b�p���� �Ê)@�@(���!^	O(I;��G�񱭢YF�3�V���w_���k��c���'��'R���Y,s�;I[x��
�'���	E�CE�u>?,K��,�*ő����u�V�����	PKf�a�Z�������踓}do���D\&>�jN>�F؞�ǆ�=U���;Rf�[�j[������EZ� r���!_ԇV���	�~?@6��
���;Sז�#�Z�k��ݹ$��vb`�R�M�������}�K���K�L���{C��y��Bɑ����ˬ�Oմ
ʉ�W�AlN$3E��U��\z��'�>k[e^�dء�k9�����p���g�3��z}�A��3�����=�DP�.*@e���~����G�wh�.lOm���`Xd�����C9x�e[�����j7J��"x����5N���m�u2�y�Ղ�O��:�����3-a5��O���z����G��Jd��ҥ�*��$5	���̈�E� H�20i������#^������?*@R�qjR�Ӳ�n%IZ�Ň��hD�y7*5�}_��4�v�O �y�TՁ�e���A쯢
��7�n����?0���.:WZ������I�<�a�[�Z~�Y+$�J�	֝LCY����a5�<�o	���A�7fw�H������u��WU)1f�i���~	�t�{o�Oɨ|y�76�F�愙ƪ�\�� -�������#"ᢼEn�8K�l1(�yҥe�8�"x�'%}^�?���kG��u����r�Z���l�Xf���� �K=W�,L㰘@R�BP�O�"F���Ψ�C��LŢ��.�Y��K�.M�e[7��d��i�7��t��LZ[���UA�6�/��T�ٱ{J�h��>;�;}bo�ZDK�)tms�|1 ��y�#��AyqŚp`{0�i��W�{jd$l̢.�J6��jcB��.3���~�L?��
��7�e�a*�� �M%�"�y#���S[h��S!T����gt#53�m�??C;:���V�V���cNr�B��u���){�Oj� ��� צ(�o�X�7@�82���L���4N�Ĵ��ÚGI@�K���X.�aLI��h?G�Ċ���<�Pb��Tؙ�;ֆ�G��Pc�q�6Ĥ����L_�����D>�X�<�s]-�Q
&�=ա~�ޔ) �$0`�쇄X���"W�^��Q��️���|U���is��qe���.�*B	ޡ��i���k/��]  �¸����oÿ�P�K�f�(�_�r���5�#������>P��������0�aB�d%D��Sԝ
�;qJ��UE��Ŧ=���7ќ���	�������@�7m��	�lJ���_ȩ�mz6�Jk9�YL�*g~���|��*h����}��g���?�����!*�F��R'�4�0����2��,ӳޑ!U>W�Sϛt-��LN��i2��g�7�N@��~��v�{�.�ٕ����{Q�tkf8�5�4��8��J��z����G؁�lj�
�
�?H�o�j��{�p;x��~_X�!�I�es��>�,�=�����쳶` �V
�wt���x9�5c#�X�Y�����v
��ɭ.�ц�x�/���v��p%ˇ<�5t2���2�;x3]��e�Qk�ӝI~�w���Cygj%���q)����ia#�<���	�d5}�Vy��x�b���܆��5oX{X�4��ut� y���b؆}������L��{�"�t�����&��R�N����L��NIm��+J<�P:~ྎ�K��!q�f�M�-�����FjM<h���Ob�̵.ĩ�"�*4��!͙Dmo��Y�8ahy�ZP���+˔��L �V�?�=h�7�DՃ�!�W����uUE��Q��rQ�$bʎ{&�C�q����`��6b� ��$����"�������ox���莾�M�u6����5h�&���?���� ��Rz�!8�!�D�ń�����a����K«\������S��Ӻ�Pl��φ��iY߬��v�aLNP`7x�b���Ұ(�j�����_������(����:�
kL÷m��0���ꁠ��Ճ�u�͑�t,��_�8B�x���9n�R��tBq�5|��kS�y-:��ت�S�Ӹ�~ݝ��[$e���3X�7l�|~�.:���U|cC#��B9*&���l�r13�"ӳoz���4Bo._k�&�^�-s�e�D}e�%J�����A��ݑ�œT0�z����	�;�;>�b��B�E+cNb����5߃���y���j<6&���_�D�\$E��C1f�6S<�~���D�����,��� �������5��3�@I�E5(����-�H��A�:�>M���6x(;NDUp�@#��m5��G`��8;V��	�c䋶��9��A�#�bg +�2��0��s���7/�o9y!����D�y��41����)��9����%F{��Tң�o�g.�{݈]����>�y�鮏�'Z����ڍ�-H)c$x>�C��ݍ`V����R��0_��N�m�jC�o�+��d$�v��+��������)e�&B��1b��RbFE� �T��vW�~А�J.�!nL�lK��T���"�`b��Y�J杏�<51�j�^�� fѶC�N�m6�d� T����Ŭ̍�Aޔ��>Z�ʰzеF6�^�N E-� ����%�ޘ�C���m�hK��T��!�g�N�v���Ɛ{�vJ���9ſ�SM���n�g_�[�	4yi��[_��q�����G	�3�91��K@&K����o�3D�*$��,A�����a�:(;�	�ˀwn^_M��i�ʒ�  ����.^x�c���x[��(�x穅~j�k�_�H���@2o�[���� 1���O۫�;&�#`:�p��[W�4j_��o�u-�u7x��,�����FK���T��g�;��7�|�cu��0C%(	Y0��+Х���w0'X�W�l$� ,����h�9s3%��%8����;���&�}:�ﶏH{>���Sم�+��&Ą:��j9ݺ�5�����9�>�r�u��(�����n{<M�祣�yS9Nor�o�j���������s>g`ƅ��\nf�Y�1��-9T�7jȟz�ퟶ0[��Ϗ��K�uZ���a&"���`�E919�`ju��@!�x�A�����Q����@oF>�zY����Û��~8&����z���z�^= l��	��TB=�(���;ͤ��hB�^X�G��,��^y����T]�� I倥r�o�(!�n �a�Rc�2vO�j�� ��^aٯI��/�w?v(�x�$/܏����F�C�2=1|!v�f֕��ǘ���+���:��
4��E5���%t�\�Q�ZF�*mҦ�*@w��n4����Ed�71넀5ɬ��I0��ᚨ(����A����9t��}D��I%���\Ҥ��$i-iT�
���ad���
K�d*oʻG>�]�� �S,cM�R�(z[͖�K��B7hj+��gE����?�$6f��A�$��n�!�u�q�"e�l��m?���4b���Q�������"� P��?Z1%֓]���1���|�>c�<����뮇Ύz���REN�[�K�(��W��ƅݺ����#�BL�\��Yր*A)�TYH�]�U$�7��p~Z&xSI��(��++��p��Ғ��ʹr�i���G��כ�'�9�b �C�b#G��A�#' �NԫQh��E�`��'�({���,d��L|n�J�"�����x=�r��i�?_�~e(@��Q{�e#����I�t�_�*�9���w�Oo�=u ?A��C�9�+F� 9��笏��e�d�DA���_��� ��y��Ĭ��>��$~�oֻ��Q�67�âk����o�Q���X�]��6�_HSw`��m1�/���V�ˮ�Ի����CN�m�0%7+]�.E8K7�t�v׹9�>�9�3����]2�W�mS�y:eI�n�����R�ރ�[�QP۔~#�u��UYL�iL	� ��W52Z�ah��Y8�����,]fY�����Qrύ����a��c��m�uO�U��_Lv�0���`�BԐ��N}g$o	���o *�M��s�����R��[s 6�DW���2����p���)Ǐ�����P��ת����ׯ&��E���qg.�#y�4΍Fw��߸��SB��ք�l܇Ex��Vn;J��f�ʤ�"�Q�Q9={w`��74!�p`��c�7g��}"VZ5cpA"+*$Z�iF������}B,��J�hF��u��V��	?�$d#t�3�ၡc�O|p@˙�w�f�C�a;K� �����s�8�GA��)V[���?uB�U5��,�xC�o:)q��M�.�-�b�ޢ&7�*�+�+�F������I%{�UN}�x���͡J"��sߠ�/��+`�Ԇ�d�V3{@��RFh�wu�-���]
��?D��ؔփ5�b�eKfm)]+�<�-(4�:��e�L�RIw-����
&�y�=�-���]r|ǵV��*X�6�}1l ��d%����oC�1h	�r/H��S;�y.'w
.m�6�c#D&z����_[���!�%շ� ���V4;���8��c����?v-�(�sk>�Ｆ�B`�y��9Kl�z��)^b��&��I+���2/��~̨�!c����~�2y����^�]��a�eCdV�j"�ꄔQ4 �Ӆ�Qv��:R�e�w���q�F�8Z]����6����q���.F��-z�O[��e3���0:C/��@r��ԍ�SM���,(>S:]�P�Ab���)��)A01��B)G����.Q�f7���G�$�S{�1��T��x�R�3p+�(�������	7oyxf+�+�����ʯ����A���)j�
��F�]��[���jx�X���V����R_���i�<�L�e��$�vg��4ˋ#AL�s�/���Raݾ��E���'��d%B���>ŉ�1,N"�^A-���&�?���tպ]��+}�̑)O��9�'U:��BG*o´�R	�:Me��+2��d��:f�ì٥[�Q�����@�R��D�^�a-�Se
-�8(�r�J5n8X����dS��i�e����b��X1���<(�}�xH�a�ʠ�LE�Ĉ	����S�uh��@́���Z�����'�̛mݗ{�	(�7���!��g��h�h����~K٠=������xaki�+*8W0׾�u�QR�p�z];�����c�4��S���c��b�+w�٫^U�|�X��65�h�.���e�
��|J]׳l�?�~�Du�Q��ƬH�U��f�S�V2��
D$�ts��&��O��!w��n��.�P���qu�|���}�<�n}!�@
�$��M)n��h��1>�콺#�R{�3�+!Y ���^��Z_�O�ȼZ���2��L�IU����QCi��çu*_�R�J�F�Hʣ��޴�l�%��b)׊	����s+P���o�+��֡;�n��tZb7�+l�E/V�˽���i�:6 ����J9�gZ�܌p�N#{�Z������-�:���w߁8�o��{�"��C��D��f�w�L�7d��kq������%{G�j&�L�Bt>O�k�?����J)��yi���f�	u���5z���!��XQ�A/�g��m�"$�ݝL%Q<n�֪����\�Pa	��K7���z�Ƚ�zR*r"wůB�RRπ�_m��J��+1�8�V�T2���w?��c7�guzj&:�cClK����g�!�TT�;؉�9�������9 K*�P1��n[�ah^¼�P�*gC��*=(GO��X�-eY���A��.�[y��M��'��/$���7Tn4�p$�%gu.�=J{EU�oއR�+sO��oϥ0Hqqk���6��A��/LM\�iLb��	+a箝��1��.N���`�6R@c%�o�VkY�3%zE���ߥ��2W�+�T�������&�/Ǽ!�e�?�c4��#JD�+Vᫀ����*)�� 17�tr�{�����{&��1Ǆ�|�YP����13O��r�.� �&�� �u�n_�D�|tK����|Z��I^(B9	$V"�v��^ɧ���U��s��]���$���)q��Cܭ�ds�;ײ�Ҷ��&�4�4��rw$E�
<�|���ɗX������/�����iޗ���51=d]C�8=��� ���V��e�� �e1a�,V�]+�Ԭ�����~'B]��5��u���:�%W���ך�}��>O������ʠ\���U��0J��Y;J��V���Naz-��1�Mm.X-�וª/j4�p�2���A�H�=�m�&�[1�
�Zj�=�5tHp�ز"N۩ #U���'��RWv��1��<�s<>�	
������IQp�\h└�oGڢ&�Aè���ٹ���	���[ ���wM�l�Im��s<m؞Ã�����ณ�J�W�Ld�o���8����C��ܨz���MN�(��I3t�,w�Q�'�E�$oY͉�f�j�s\�g�bZy �/�޴�?�:q�v,u��Pu���P�}��29B�N����?4��e���\�\�������uJ99|U��G��$���,-�[����Y� P�T�m��:+BBZ�>̐�ZHT��{#���v������6V��M��՞���N��5)j|{A�*��B��RƎc�j�������m	�%���zf�?��h#�`-D�I%���;�"�Eo7@��3�oX���
"�P��ǏUÂ���tt����X�->C�Z�.EO��IH1�;,p�4~8��+��h9�m����DA.�[0d/?��k A�+,�)����ʱ!�7����o��D�8�v�X��IJD�PI�}�W"��6X�eyK�3��P��7����_ȉ��&��'��ɡv�sݺ	���u+�3b�עcf R C�҄X,��b�ړW]����*������6齅����5��1=��-���~ �kBVNM��4νnWs����w�=�Ҩ�1o��r��E���Kk�Sr�
<��di�8�Z�|�H<"|ɮ{�cѦ)�k����V��|�b+�T�Ǵ�M��x�
���΀8��Ga�����G��_\�%�����j�8�g⋱���#/4D�I���������9Q\�����@r�e����|��-2��pCLQH#N���{�J��琞v�lA��u_���q8����TI$f)�˿�g|�q�;��2�4δ�I K�cY������Amب�Ь1I9Vf ��3>�"����2?=I���I�w�Q���1˼��� >B540��~���GR��L�Nts�/$���Ｂ����>h���(cDl*�2��1"oe֒^�� ��m�FǪ�j�~Gp���������Fc��h��jn�b���<�	`�Y-5�^~��SD���'=v!s>�A:�[/�;,���=*���j��C�茧�C�e�ip�ZÌ@uEg�Eƒ�\���Ǆ��jLǛ|�$��-	DE�U�c6���3!��n8��eY
v�x�g?^�٠�P�!Uz��b�p��d�q�	���(�Q�=�Y�bxKώޯ�F��WA+�c�����?�l$��[��|]O�m�IW����NګNE5cƏ�)*'��{�*ͥx5���Q��|�.�"sÆ�k��x�HV�/I��Y)Ālʫ����/Ey��.����}�����jMλ%�,�I3��hn~�Q2�ce匇	 ���.���2-�$��+���ʴCx:e���/��f3��{��7���{O��W�a:a����VM\��Z�w�
��S:U>*�x�˿�AQ6^[�M���HvP�����.!Y94 ĵ��{��	�2�Ĥ�F>�L��-E�o֎��1�uG�4ߺ��E7}��+ۛ�a��Tt)��}�l�����_kkUԴx2��Ua����3�zz�׃��0Yr7٧R��l/���"c�����rU��0zQ�[��6����. ex��x���R�D��w ���zĎ������4��"f�Z�5�t�xТK�ެ7�f�1:/Q��N�Q!���Z�֏̣ޝ�e��/t�]���3�������W���!�@׼���r!�,r� H��ud�l�_m9�|����J�f	���J��q*�箟������,�WuRL��r��	�
�N-���>n��!�|��O�F>;YFٻ	l"�^׈Ms���$�hȹoj=r�O�兖6I�����k�Hv?�t���g�v��_5��u4���s�oB��cA���9�{�A�re��U:8`�z*Y���f.:u�e*�`ù[m- �.� �����ƪ��e)
$���sE�`���%���ͺ�ʸ���$����;{�ra��ePE�>]gN�}H�|����~G�y��C���B���ww*Tv���C���k���B��<�j7���6��� ]�}�n*Tg�@�A��f,ף��
R7��kE	A�w�O�^:_s|4��Ƌ ���K��ʂ��O\_lo,;3�1 ��B%0���2N�"��ws����N5ej�,�\�qޯ})�ļ�9�֣���X��0�ݞ�=L��(r�����O�*հ4_�����ev+��_�u+���20y��k���ե^��/S/�E9̄�ms�3%�H���Hj%b�m�� �`��n�z��鯙c�ghU�\�[�o�r�ab5����i�L��3�28@n9?��5�͠��2$<�2��1؂�9=������gD���C�f6t����rh�#p���ic��A�iv�����s��ٟ\ ]�[ML�?�s��?r�t�NR��9�,�-���x6hxɔj�[���9%��HjF�
nw�lPz���	�x��5w��=��s�<� ���������DH��HX�����g�V�0�U�u">�b7���;HH%�$#E�+�Gra�{n�zD�.�@���P�*�c��E�����C&�5�t���^�/-��N��@�~�QrzȻ*e�,�[�����F�#g�K����e��O���m[��bWD�8'��}<vQ��\8����^�&��Ca6��*i��W1.�8{���M�)�ʠ�Z��Г��Y%ꤊ�عst���©
(_��t/�Iz,p�e�
�R���Nhi�N���^Vǅ�?�F���-Oٹ��^�uT+s�N��9/�!PWR]�����+��Z1�^. Kl�r���Qݺ���&� �>a0n��?;3��%g׆(�aC��Ĩ������4�Vn�H����-��(#M�T���d�wyl�|�����D?�p2�O9��6oO�]���6.���U2��"&*���vac��<��P��[*7����]-4��} (�(?Ԃ-n�,��<������Z��XG��`*�{��4t����`d݀���D�g�YF��Ԋ{/��8��pKs{9}�c��C�a��.�_�"F�;Q����e�N�-�jp\�����2y"W�ɭ��x��u��;V��}�A(�/����F���Mry�M�F��w��1�_�^'W�d$��O��Ș[N���=�o�>?�B�,�KN�9�Ga8�'�D�J�ۤg�C�kU���"o`��x��^Ӝns�Y�<�s.g{+�y��-y�R�KDA��f�d�-�.�����?8=�(Z���+l���]]��d�Q�30u0��w�gi�Yܷ���ᵝE��*`2�U$�V��H$�̈�ҩ�{��5�7l���&�Xi����(-x�G9?>�e����=Tr��5�#��w�^)~k���`Ϯ6qc�ǀ<	;���a�F���~�
i@�o)���SK02RԻ������8m���n�Ǌp�."�4��9�����eE�HL�L�⡺jr�����ȫg1�a8��\A���=�t��I=���E�߇�vW��J<͖��Öm`�r1��LKQ�*�p3r�<-7:��� !�9���|Ԋ˴wW�럟M�1�K�p���Ky�F�0��| ���5|��|Yf}�����ѐ|��{���I�a�+lo�N\�C�m�5�k�C�ꔈ�o�*��Ξ�ŉ�e��t��-��`釓k������DJ�%q�L��ދ0����^"�:��u����m��t�v�4��4��ՙ�l4d�7��~�p�1ۙߧ]ʦy1g��t�]f�<w�T�O(�@H���)�/��!b/v����[a����O|+l c�G��h]�ڿK��*���?����,v��h��o�����x�����&��̨x���g}y \�kE[n뼪�>�%����zh� \˗��=��RFxP]Ev4!�htt�Т��0w����y󯖉�P��n���=�1k*��u�o��ȹ袩��E�I��E�%3w��m��G<F*���;��\����W�&�\�f/hjW�R���]��)
W����H�h�]�۫���һ� f�ڼ����:X���|�r��2^Sx�s��ْ:��]Q�Ŏ�2���SH��ݞ����KPF�B2�>A��ƈ��u>U�o|S?�r��@ ո�9o�p�X��D>��˫�2Dԍ���j0:멽^k���*�p=!��z��,��ѪC.�fc�)?�3���etq2��HSSB���G
�6[��dǦ��� �w������ޘU"��g�0~��^J�F?���k��sYyӴ4{��1��7rP�Q��ern�1d����dL��v&6�!G���W����ΏA�-�%[�������M�_L/�1�5f?� �1�����a+������&h����"�Ϥ2�B�.�;��?ie�ް�?,�� �Z�Eb����*:f�S��G���G��ph��|y���f#?��9�y:<���H'�)X
>N�5��O�K��>Z���i��7�!*�В�ԭ���͇��r������f�n��7A�+��?6@��.fe$��UI�2+L玖��$�gIp��и��<<_��&�9���K�9KLl�;S�d�CL7�u��PFi�<[�{���S�ޗ8�=��&<_W��[���`  �����ݦA4��WÜ�P!�ba���X7 h|պ@��o�>,�+���vQ�D�,A�iT���7�pE�2p��_ND���iC�Ҧc&sd�/�Ei)q����xC��tTY~�\߼��f��ݪ��^��c�Ӗ�,��E���A����#7\[���p�����C~U[F�P���=�p^"p�����	��%�
bq�$J/x�?�Kr�p��Dc�ՇȆ1��n��=@��ƙj�"���)���Gf!��9�62�|ot�b��N��{���{e����]G۾��9��a���}��*���d&�Mg\����ψ�a�#Iy����8̯c���إ.<n�6�q��v���}�i'�"�,�nY�bw1&��̘Z�\9�F���DJ��#(gt���0���e���r]Ap�qTϝ��FqJ��͡@n�
�I���M'LT�`����e����s�BV] ^HTHcyhl�e��I{�0�3AA�K���v���X�:�.US[�`�_\p,}�\�`l�x�[���r�,}�(���^goJځ�l�.�����Ki�qv�s�0j���sR��n�U"�*b*8p#���F��n���N���ދ�����r����JY��$=qв��!����T���Os}*G�ש����g��Q����h��������I?��L���&�JZ�9�^z8D��T��
Up�Y��hn�*F�Z�JZe�Teu�g�B*5���ĥO��#�_�nZ1�����Pi/Y� �h�����֝.�]�|�����KGn�����v��!�H��O<���94��k�Pz�w��ۙ������-J|3�WϦ��Q1X=���s~t���LB��h�B���=䂆n)N�n|AS9M��aRć�+�	l ��y+�٠�&Z��Qؔ���B������?�1�.w"Gh�@��yW�$7�@mr�j����_UcN3r�{i	zR��ğ\�ޛ��'u(势�U��j���@���H���[7��,۞�+ˌ&��<'/�=��ś�*�'i�w�7m��P�~��M(h�&���Fuغ?�Q�BT��7fJ�և��]
�S	kϴ����n�� ���B�64�I�,�Ƽ�t�q�Ǡa�����.#��mmb�W%�5-�W+�lڥR��w��؇�^�򘯨��<����`����h�҃��aT%~=Ǣu6����߭_���L��t�xM��,f�}p7�R�/�E}�m��j(���e}��H8��PqO���5�l��2���ƺw�L?�2�	, ����媓s�$�(I�Z��Lɧ���;�q �gX�qf���#m��9ҞF`j����%S�u���]���2-D;j���6� 2wD�C6I�l�9�G-�+�{�vY��2%nO��J�f��	{�����m�"�3�2�o����1�CI���_f��~\�����{K�LA�7N�7/B�f��5+MqZ �٪^8�~��hV'��ĬD|5�?�����&���,���R�D��.N$�>q����&�����a@�Hd�2�{vk�K�l[h��?���~c5
ň�z��N����������q�И��>V͏�
����+�г!�.lA���V�IW�LX����.�����P9Du|N-D��ڣ��ɲ�R��8�a����	/��qn=4[��Fz�Iy�*�p������47N�"��l�=b= 8�ѳ�ʋ�Zh�<�֕�\ػ��s����i7�$��?��D�|����fG�dB06�	P<1e'��+�Mf"��b����D7�:tO:��)�:�A�� ������_�A�	�L��T3\1����<��ˑ4��]��S^7��r:q�B����Ŷwg�+��Bbaܾ�,��~��x�����Fq��Z���V��dܵ��zC0����CE��>�B8E��o��(�A4�٪���ª�(�9�J}B�*xuL���91��9J�
�&����g�<�:�(��*h�0�x��E�
ɩ����
�?S���+�-�#�� ����s�Y˅��4���d��¿
�8ۯ�F�@���	u^S��\�LV�+V���R9@W����]Ԣ�:��G�WR(.@'%�8�p�V]y�ѝ{t
]r�.�6�u"�D3�,�2ԑ;�"L�w�#��/�ϓ�wwU�* ���e��+9�}���"y~ź0r���O�S����!���L�b�U���f�� ���0�D�e�������w�$2�\��Ƅ��&��g�/�u�`�5g��jr��ʸl���oʔ���Gm~7��y�&a��:l��(C�L&���h���\����L����B��a�d�L��P����|��W�"[��N0d��2��u��t^0_��`6�kC#�`��^!n�R1�/��>����f/�K���ԋ*3F���pV^�eo��s��k7ˬ� CƵ�k���FS�
�2��5��eH��9�pP�a��]�#����'���R'��5�-d"�z��v�q��*?�P��WKa��3��)�r����h�BY̤l!�T@٧�k7�7�F��ÃP�r`��:`=���+rn��p��Ӫ�=(A��u$<	�����a~�WK��C���d�[����[�]I��w~��e���I��Y?����<�H�g��ML6��fW�ӕ�^�bf 4�| )ڡ� �ᵴÐIl��[�C��]��"h�U������
�0Ur}~������N8vPq>G�PZ%ʰr,{�#~���e��ا�Ϟ�N���R�
X���q�z�Y��S.d��c�\�bE�'�e��ER�/�Y��9�0��c�g6�0Q��Y��A�ص)��I~�hi����S��ogۤ�]�1�.@�;p�d�)$@C�*J�H�oM�I�Ǔ�}�����%huM�gտ�IbH��S�Y-
&��T/�� �*~�Uj�r	��?��#��]�q�r̓(�l`.�,V.E�z-��G�[���O�B���A��[��@��'8�<�l��y�S�2�7��U"W�ikM���}�;���D�����|���8��D�������P��qa�wd�bAvh`�����FH`�u����P�ʝ}�ots�Y��NpS.4A���Ri�/F��#�z����@�������l�ܓ����V�?�<B٩���c��7S��tP;�>CvK��h���q�5N����:hP� ���EC �S�tkNp�l������[6�m��A�Hi:�T};��ggK��
u�օ��Q��S��g��|1_����N&�J�k#��8#~X��.��,�B�sM~�>��� 3� @�)��<��Yɓ�l�=]�i���9O�[��d�@���. ���킦\���#$�X��ksn?���C	wWm�W囩4;�����1���Jhp @��:"�����!��1u�,�'�P�?a����K=!1^�@R�Ό��B�/+��y+��˶8��2��5�^�����]z��>�T\�T�N��Q����P��Q�����˖�zM�_=|�r�8n����p�:z*Im��L2��4�4e$
KsJ�.B�'�+I'�-^�dR̎=6S�^����c�� G@m~�G�{C������܄���,N��30C�c� $�|�#�RLK���H9��3��]��d��X�B��$�'�t�R<8^�=W�~��cy���l�����E7Y�Ӌ6��}��I�v�'��F��-�,�wPЭ��g�����sQ�7
�7s�(�Fi��h�~�쐝���y�Bãԙ����&��_s�m9��w����AyJE#��7" [��� �5��p��@�3���\�0�!}x5����Do�oG'�P�Ӌ�8��� �9XO�@���� �s;x�'Pr�4K�1Ӛe�bmC>�?����8J����,[�$��dتX��)z"�s,�2�G�Ut�x]F�OXF{�WOͶ+�.����
��T6m~��x��g�&IioT�Ұ����T�^���
����|"m���{2��:U3V�60�)��W)	��v��բ+@�R�G��S~֌6NϹ�����ƒ�)���j�F�ז�S^d�)Ts��w�L6�U��SQ���bP1��c�$�a= �~�`_b��GU4�s�P��rZD3�7F�)i/�ic��{wK(G�@�"�RdN� ��g(###�B(���)��nc�i�S�À༹�?h��ԡ�׷+�Z5�Ka���F��X�̠T�,�ՈF�Nߤ�}��/�8P�6���_xA�Y��F��_γ��U������٪��j�f!�)0DO!���8�Wt�-���t���d{*6�|X�v��Vm�GxG��0L#V/�A�/�@TVY�J�-;_5pM+��R�Z'A�;��5>e��ٶ�r�T{�,���k���ғ��A��q������JM�@�w?�,��o8;��)��/mk�KyFlHG{�X��m#�C3�����E@�ɏ�Y�7h��R7�U��1L�E�ds%�_��s�٫���h��< Z�C0�����Ͻ�'Bk���ZrcT�K�K��hW�cA+�.V���R��##�"x2����h)�4��Rx�̡Q����@�"��IS���qKw��[H2���hl`�`&�e��pb��e�h�3��Lh�5	��+�Ă�jU?��Z�9e2<�W���nd����ǒ0�g�Pb�<p��s�^���:S~�JN��^/͗[&�֢G|-� Py�vƔ�����bk�����:�T|HMH28�e3�o:���.o�)&$���2ٽ�\��پ7�ġ��NMb�����ԯ��'!���q���r9N�S��,���F�ϴ{��51�v�u1�ʒ|��'����K3V}��T�������<����'�<���(O��VZ�ַ8
��HW���/���wC������H�yI!ډ�v� �F���H]C=��Y�O7�O�����8<�����Fgy�]8V��*T`;�b{���<�+�/�<��`(b�{���Ӧ�D��m�}��_KM������P�4�8Lpz��� �Dl���S���o��ɓ5�xs;$C=W���5�qA;��x���-r*��)�6� ��ɲ���ˉ׼o����A�=R �hN�h��C�+�,w<ֻ�Z6&�����]�S�N{��V����&�frݡFxR��~���$�&x3o%%�����8\�����P��JV#��W�n"�h�D�kD��L��)����:E�Z�Mu�kG@h�S�?;|T�.��U���2�Z�:���W�2�jڍ�W���MO�k�C�Ol��L�7��$25��'�$�`�������)�����"��ih0)�������%�Qn����
� ��]Z�Q9%1��!��%wɎ( ����ސ�<7��Y���{�zSP�8@��K���ٿ� �\�
J�@����rAq�{�
���W��#�i�ç�3N�p-;����D�	d�'$2NӦų(O�܈�p�p���SW���N'ɾ�+�RyV�V+hM�U�@w~)�c�mR �TQ�3/KT�*6ݯ��8`�+�ɰC��� L�5��0�Y�M�»�0[�}��!㲨� �Ș��Nlj�P�J�f��wb�HKm#�;�V�4q�֬�iX�C�v�o^��axNJ5��|��6��^Eh]}W˨��Uu;����ǋD����2c�\��<�1L�E���	櫥��#ɶ���Y+��1>����?wu��N+��ݛ����.r��V�'V\f���U\j�F�E���U)�b'FU��	�c?����GL�ޣ�T{w��24�~�������cl#����χƈ�Dp~FO��AK-h�#W�
�a~��� ��qb�;C��_:��:�ƎA�~�������Z���R2:���r�<�Y�s+1#�'��	_o�%ĿB�א�7�;�n���CD1�?~iuq^m�x�d =�ſ��K"�/�.Ư��뇜�9A�ԅ���N3;3�F�X,:�<���PP�Ռ�ucO�O}����,9�f�D�_�U'�@�:�� A&fR�v��w@#� �\e��Ӫi���Y~�=��?��?|�P#�� 3��ՂE И�~����Vab��9n|	'���MF���|�e���$A�#ؿ���`�><;<�Ij�9�P��hR�S��^�O�1�%FS>�Q�=x��"�!�q8�psJ�<L��#�RM����ס�/��VvUq�I�̤(�l��bJ�)��Io?��.�!�L%��b��}�/{d�~x��3Б�^��\%��U�c"�yE��;@�ݤ�&�=�*8״^������p"��F�wrGJց��R-����*S��3)n��A'&�a�p�W&�|���%JhF�Ya)���f�j��1��q$C���G��vV(�=Gh�W 7/�����ݫeh=ԩ,�]@�&L|�l��Ū�^Z�ɣ��F*�s(�C�Y��6H
&r�m۠�I��� k��7ܵ1�(,�>u�����g��*:�Z(��{�PKki�?)��<�1���s���yO�����З��lz	%Kh%�i�����b�C�R�%Ztd{Q�c��v��� �X�J�GN�+�ɧsx��+oS.'�=�"�Ώ�%�?����QB���zm
|
�$~>��U���i�Sl��f��^�v��9z!��6�?@�G.W�F�sC�DA��AB��{M��I&G�9���l�hǩn��G�6@�C�V�?�	���2�E0��*;>d1�?�
����i�c��Ÿ�cP-����������s��H�Y���5����k>��\�W��Iͧk�j�yA���^��S �u@y�Tk���k���VP���ILY���Ɓ
��G�����{?F"�b $��)a��d3*��_>_�ݭ��E�[�y���IDg6���#�9�����Ծ(���f���T������ѡ'���3�/n�u֮���v��6l`�LH嶉oN��9�����F�:�p�c�� �eD�$Y�qU�f�����X�?��a���Ib�:0~U�'�<A�Eů-ø�L#H#O\�� �t�4��Lk9��0g�Mz�
�)�x���'��0���k���\ݼpr�{����I�Yx����+��������h>��M;��� �}��4lхB�������G4�h�%JMH����T�����۫y��LB�m?),NAa)UM���qj�E�kpp16�x���[��XX����dn��֬�W�����pJ�Wsá{��+f�rS(i��r�*�%b��ldk���<PAs��D�i��"Pb���p��0���?�Q������Ym<��1�9M��>ڊA�ק8q���W偻j��M�������m��_�|4�-+�-�|���Њ�$�δ8��C7���e6�bf\g�����\Zu��ap�
T~j��$�����5�l
����fi0Il�'3�?��q�4��e3
�/C�!�;���K�E��w�ĸ1��O��ɽ|���9*�_��ad�@E�y��L�{ȅ#�;rrȚ�B��z~	�஖�T	�~X���]\�A�������Ae�l�D�L2\��FO�e�,��ЉLz����(��1���,��{940��2u�F/
��+��q�.�����&y�E���iM�=�P	5k��Nif���h��۔�4�FjU�);������]QgX��}y�rp�^6^����0!ǹ�?���P��GkR�;��e��?��
����<�Ep�'x|�H���~5��/��$�/�1�nL�n���; ����R.5s������ �Z�;q�CLU�]�@�UN��[�Ғ�BL �D�N��۩�s�,S�Ω�l�&��o�­A�ll:oىT�"c������������KF�&�τ߮��uq�:��s��Lj
]tw8G�eܱ���{>wW�"<���� �O�Ԕ�
�Eif{�;�⍵O+й�maq���� }��O�5�S�K����m��a�Kc^�����d�Ixy�>����S�7�Z���v'�H~�˽!7�W>8Jj����7*VI�;#��c��Z�����ӆBG(i@j��'5+����"����I�/V����((ӊ�*�4G��nX"�xT2���A���P}(O0�>��<?:u��2zc���1w�V�υ�g<����
�~ϐ��Q��9.=��f96��a��F��넻��W�Ue�,��rV��ۑ�
q~]Ph��4�c7��-�s�#�������V���c��bD����If�j����,���:�p����h�Zr�t���g�r�Q������ ���x��[�ѡ��ы�6�?��ϴp� �!�p*}���Q�Q<EE﫽V�V1��̃�@��9��(��x�H5�-\��d'��6��< �	��;V������uW�f�(A(�,6��O��C���$�Yj)7�23rp֭���� �-i�yH��{ϩ��}�Gp1{��W "�
5���]�=EcY��٘��g�#�S�[�>/�ౙ�-�{/�8�W�JnI4}ɒ�LzzӋ'��n�S��3_���u��H&pi,�΅9��Է��9U^�T��������!G-�^���ho��7����e��0Ek��1���l'n�Coε"0[e������[��b��?4��=IYU#�}��U�j�^�=�XwIz�u��5��Dw���M���n�P~���d	!p�=�S�����Ma7øV��&S�����5�q�B^O|˯ih�*���(y
�>����d\i@z��V�m�*D@c�;�E���zM�ÿ�5�j�'�2�P�<D3R���oU�˴��_�SI
��K�}ǈ&�)��>JvW?N>[!;���߂5x҄��!��x|}��q�6(�����$�E�����r��%��Ӌ�rN���~ǹ��a�"�� {�'�weFƇ��o���|.f��?�v¶u&���g`��P��N���A �<�E��-�5o�ah�SkOwHI�c�*�<f��^][�&���`0�S�IL�B, ��@U'p&�#o�R�����(Q9駭{1ղ�?S����g��E��{]-�*���tϖ�W�+ee�v>@ɽ���bg�z��2����'p��*Ԍ�-���}(X<a���=��R
&9눍��9<����"7<�j��E;Sl�&�0�e��jp�������T�K�׮Ok�Ѭ��_O^�}��@-N�U(A���s!UT`� x�k�E-��t�YV��&�L���ُI��R%���y!m�Lk���U�C�Lv��(�7σհj6�F�X?%��|��e�P���P���_��덵��[���mbC�#sa�Cf7]��W��!`�ߊYn^Vk����J̍󈗂�0,p�b�*�ǱT��Hk"��j��l��_|M�%�y���3�QYt�]f� 0{ľF��>����������;�� ���j`Wfp�>�=�36u�HF,���������w�抐��� !����EP����yX^�K�� 'p�����3�B�H�������+�D�\*�p8�AGVyU�	�S��p�� ���Ж�R�}�0����$�x���:pKT���'�1�E^GС~d�Nfp�����ǟ{�.;����6ћ��H���ڔW�C"��&M�z�jє�f���
;���d�;؄��l"���3��Ȋ�J�(�-b��"R��ƤZ�����ۆ�i�!� �Ϡ����<�D+�L�e����^mfÂ�L�&Q��Yu�����!?�W��m���n�bY.iH����d�5�\R��Z}����B�� �yDr=�b�p���ԧ�[��Z��thl�Ho$6��ۺ>7z���ք�t�9I^�N�����i�]���|�Q�Vb� ?����YBv�={xn+���]�?t�<�!�S�ռ��ƫ�����
3�<�x$��9��</�\9���5.(>H���~_a����v�X��,MS�����?�[�n���(��R%����������l:$ԙ���ˌ���v�N�f�	T��x���H�^�x~<U�~VV10o�}�Iy)���y �	l��8�q���V�[(w^��!~�a_u�
v�D�f\g���>$1ۃڄ�Q��\�E��X$�u��B���I�=��P��!mz�[z�@�!K���_"���S�{!�6�94��^�q��$�ME~��q�l��f��)B��[e
���'�
­��.�3Z�#�N�v��]��|��A��A� ����eNԍ��p��~�)ce��C�r��G��MC��w��~)��&i�0t}k�*{� ���A.�0Ɗ���\�1����EYB�{��U����×���o���&x�����z��/�E=u�\���rs�?�H��.��΍��ȗ��]mեj�����4b/OmҶ��0hE���eZĚV::8�zi_����K�V�(�#�ݔ�2T:}O�!���8;s���ۖ�j�8��m	����.~øTU(�֧��,eěVn MD�(���gw���isQM&F��}#q�\�H���u��+IB��SvDgM%l���]����K�'����	���p�A�E~�1�9�(1?����
�	��d�c6�ʰ��9��h�"hdZ�M��˞z4�Թ��کbT:M��(�t_]X�P+�e�L�Rm}���|��������3�us�s����0�_)���c�ur�tG���5�~{{���|�<��J����?�Z���.�ڒeX���(�Lc��{'w��i���0�M:�����u)������W��ĺr�(P;�N������
x��Q_���$B��'s�-Ln�[͵Z_
ř�Y�h�5|C���/l�c�g�_����U�h�����`/Q#�H!"1��G����P�NͿ�5�0sC���x��1��>��/9S(ݧ�y�&d�3�q]��Vk�{č3�F�8�t	S�\�U�=��t��vk�o[^9kY����c] "Gu�/�u0��,�B��S.�WzG�3��~�E�x�dڶ$k�	N5s�$Ćf�/�V5�*��d���-7�c:u�pέ��}�ME���,,��aUW=��tɕԝ���s} �ľ��>+&) �ҡL<��t����0H�?Z2y�Y	�N�S�騺��T� _���5�߼W�h'c\j�A9ӓ֯%x-���!3�L�x�_VDm+���	m��<CVy/���0�ߝ�n���O6��z�� �����!i�8�N�'�
�t�"=�W&��#�;�W��dy��?5 +�19�k��4Oh�ju��sMUR#2�:�XJ�/������N���{^o�hu�*���1H%�9����׶X�_�"%tWFlC_\�x�M���N����ݪ�;)b܁��cdC!(.:�v-K�����G	���Wp╿z�y*��qL���ߏ���������X��Nr�>9{戅�d����k,�hrxy���k�+��A�3wpq�$G>F�f�Q�'�*�nS<��%�7wZ��~MM�y$����F��+��C�l��(����ˑ���z`�|�FUERs3�׾7��P��b-������:ݔ�d�Y���PT��xcu�)�����N���dV��z~:�E��_`�:���2;�LP;�;��ז��J��ұ#�K�	g�e��7��M���Z�D���~���(Z�+���WWf�s	�竂޵5����<=Jh�0ei��vJ�g�4�>�ji�993���m��ݻ������P+��h@����=a�<8�����X�G�� `�%Ƙj�C&��ƾ�
�&�P������l��}�I�;��̰*�-(<&�ߕ�U�aÿ��PCp�����S���"L�����c���v�Ӿ���O��wv�=�g�߉���}�"#�}_�+���j�N���O#���������~����X@�)s㠙ιû��\5z��s{��i����W���8�S��9J��?���<��9yioN�W����uP���Ή����hGpy�����?����&j�;���z)���J�C���?���.�6Ԡ��B�n4o�+?c��U>�r�FX '�������:���P���b0"�<�����D�"�ۗ슆��$��/4JfI:��Tr�BQ���ڙ@�f�c!V�$��+[ ���q�@�X<D���n�R[m<6��(���Y*�E���B'�,���S��k�Gx��&��~�$x��x�5ѓ#�d��a���1ӁdZ�������&k@��:>�I}�專��w;��u���_1�T���f�:��nLf.�N�SMX���i
ޙGy��fJth�Ձ[z��4�Tx��ǔP�sNl�{G�P��I�m��X�m}r�|�~�ܡĤud����g#o��N���P���'���=�2��@��$��>��)��o����n�������A>�:�k�K����/?
�~R��)-�*�!��	������B�d��Rz�~�^��ja׮�p 5=T7k�ͯ�8�O;��^��.7U���G)*����/�=�3Å~�	ʻQ�n؉8�AU�0��3�4�Y��J�(��KeHٍ(���Y�ɟ�QQ�a��	�Y)ao�(�{�N�-zN�Ґ{��;��D��L9��U�IR�B��I�L2��N/Q�*��l��
��]����z507k�L���x0w��l�����49�^���l�<����ѹ�K��-�G�!��jMԘ�.�TS��6��,����ϑ�d�j�ס��H�ڿ�
a�������E���xE�v��3�;{J�/�T[�?�吉=��f��5kU&��Xim0Dj&A���6#�y������-�[�wg���>���jx����<0j�����>	xǚ����W�-	,�������:K�EiHW�I2�� Aק,�<�ALb����a75���z����Dƽ��=u���vE��c�c�Z`c�[JCxa��K� ��h���ek0B�1� Dg>�ݐ?���E4�R�G��,�8gy/?*�=�S��T�8��(�>�7�Jur��J�#!�jŒi�{�"����\��h����%9���mU�,w1fx��ӊ;��V����4��aR߉��w�0���쾞�xIɐ[�M\ϳD�.�E����}U�SX?9U�( ���N�_�շ����>��kw�����v���?�yĭ>��� kH<���}�:hj���Zz��c9v�(qwJ-/ߒ��.�:� ����Jc��X"�_�fv�%�>PQ�����ȿ@րć�S%d�6�TG���Ƴ�G�Sxk�FI�r�F���-P�ɭ=�H�*y�G��i/�J|S�D=^��%6��
�{W$�L�dɨ����q���Z|�m��I��e��_�A[S���|+��~_��҄�GU13ˎ~Nkh�$��b��#7��k�7wR���TŅ@����3Ifũ�͘��� �wK�S�I顪M#���U󭤶�,*!/��/��C�}z��t魆�<�"���@��C,c.YS-�F���8f5k� 	����!����qL ���퉗��/j㰙?ē�K2�YLmsԙN.�2Щ�33d;�����H����F���>~g$SR���|� {{��?}?�+*��o�&��b�[��T�q+Zߣ)-�vQ�@dm/��%�<
f�ܖ<}�i"bЎ�2 �,1���@�} ��uZ��M$V���"��ތn��Ϙ�-�x}���~V���c�T#C��;')�Z���\�U�]²�F�!.9��p�[�S,�oW��'�w�tZi���",�Ӆ��-x��Q's��Wʽk卐�m�l�7��@�7�<ü�2�q�·ƑH�]�^y�	x �
��w�)�/f�`�~,7�5�@`�k���sTp�������+t֊����4h78&m� �u���;�
�k��m�h3��kys:a���;���1�[�X��K���xc�I%"S�A��O�Pr�����~�,�@$�:�BA�M2���iɣ�k���~��~j�Ui��JЊA���O3���<�n�}YݜKb��B�Fz�����D��v[ϵc�g"@�cO��2V<��Yn*�*tt��i?��SyO�E��\"Rρ=�ɪyq��KTh� �R{�Rr�ut�㩌�ӉY���F�ckp(�'y��L�C,OTأ\XB��U�����������WF�'<zd�U�W�Xw/�ƦP�(�>�6Ԇ��*��V�D�+1'��/�8G/��'4;rP�������������A}I+����X
� ������d�D�J�b�K�n��EN�tH�V����˃�:y>�?du;f�
�Ջ�=u�z�p��M��/�p�i;�-�O����!8�4g�g5��*ޞ�5�����n�bi��u+�� `i����b��<��"؅��s�G�����&�5����1;^Y\64��<*��(퐀���3Eh�8l<
vЌI`��7�Э��8�ѽ���������aB��(��}��ѠM�3"���e��!�h�2���2�'���È`��Q&�U�c�f�C����/a
�q2"a��L�!/�����q���̾(�鱆^w��!eS�{�:ə탤�?#@����U�.�Ty�?YT���G������K�<��@b��j�fRQ�	�ƥ`�S�s��Q'r�o���F\p�����΀���-ع԰5��&�Ν�X�ɀ������I�h2�T<�^m��)�h�����ԑ���J��$<���ۜ�:6ܑ�%�^��v��ʃ� �Ԯʖ��lE�h��:����`��b�̃�%�v���a��'MQ��m��N�.��������q.I�K��+E�1��Ì�k�T,�QJ�w�u�W�i�qjy�C:���,���֢��m�
a��{��P��_��u�Go��L�Xı�Q����u<&�<��n�����='��<o��a����4��ʄ������Jo+٦�����>���_oh���}��Sص°5^	}Q�"F̠��C�mզ�Yq ���n�6�o=_��J]���|��;*�bӓ
�;rF9�|�9� 1�[�(���9Tlʤ#Hl���T�o�A�A$ƹ�
�4��(%��[�2����?�sƺ9 xcb��3m���(�_�
�k*-I}�M=���%�[�0>�A�n�(�y=�t�Lwd/����>�IB��w�y�R�0�Sc�جc���l|(�~Ɔ��]uG���p�'�x.t��*S�-����k�6�P��<`xCf5Gs	�jƆ�T�v�vs�-׾�� �Ь
G����L�TX�&wM�(��!f��=sv��������h�Z~������~��AE�ISO�޶��Z�ҥLLDå+�53 �������o
⣌Ά�OR�t���=���������͂D��z��;�����B.�pt4��'�'ґ�T����^)�� ���M �5p�g��紦r��3�p�����v@weK��5y�.o"�9��(�2c�rEu���J;��#�����Ďς�l�:�5P����b%AN��LC �����#}-j)ޥUr*��4u̴��}��P����N �c��I��|���s��e�,t�zX������i-�_��Ɔ�$[/�b"�'pu&�Hu����zc�ei�C��������u�, ��(���ZCpgP��7�(��;�tvU�	�  ��i�vV���:Ա1	���dd�^U9$�ڰ�n�?����R��r�,D�C0?��q}G�΃t0�J9�*�f�d�����
���[��ʂ%3Wo��e�zm^c(�g���Nol��n:ʦ�ϗ2H�!x�D�;η!ğyb�D_����ϻ��3��܍��PC_�ֺ��l�����K����P9�,tG�[>Uv,��|�X*c�	S�3���zFz�t����pn��8kE;���h���n�����UX�f|na�����)*׫��#b�>%�0Wۻ|�N\-�N�S$O���
�;o�Ò	vo`�&u5�ϕ����cR��)�2�i������\��\e��a��E���4��ά$���Q
v���5}��gs��Z���ܞ�t��#.7Sn�7NUtDuk�iw	׉�W��Q�a$
���HcjFQ��g��=[�*����!J��x�I��,o'!q֥���~nq�!�(��`:�>k�mŎ�7�͵�d�m�����w?�f��fc�5dO�p7�ҵ���уVZF�.��17a�RF�:�W��r��Y�6m����'
87Ҕ��![7�~P�y�y��� s��R˖�3�z1�B��k����*k'�k, p�x�`D` RE�vb����?��)�IoZ��
��mY����/��B���'T B�萍�!b��KN¢u�H�:(�7箐�8���;�*P�G�5��q�}�;@��7�d\���K�-F�B�Y �g[�L�S��o�6���9a��Х�pjn����9�_�	7�Cȋ؏�X딣�N��ZϮ|���� P(t�+�eU�Ut��?�e�-nU��&�'����ڎ������AԜMԷ�����g��vZzY6�6��� �Y���g���m���N���$$䶣�~��5/�&V#�´th �)�ڀ�Ge6]
�}@D|HI�	�ʸ���!��2\�V�3q���5vW[4
}<�������z�����j�
I^���<>{�i��|���V�t/�VL=G�8۴	.����-��	����`6��2gi<�)׏	�	��.:0��(:�絕���_N��rɻ�>N�)��JTI_x�Z�O�/���1�u��.b˗b(��E�9��33\����ܸzJD&����G�_��JLf#��=鳀�5�"�+�)l���v���{��'�� �1�����#�8�l�JMh2�Q�Ts�nP�B#`��%$�Vΐ1.Hr�QTX�k
�HG[�B�Q��ɖ�'���3�tL�z6���ۖ����11�=����6�D���B���Ӂ�0Ȗ+�S�ʠ�[�g<%g�����7���ܙ��g���߯$�FlI< ��iU̿���e����h��f~Ps��Z=iȝ����|�Ƨ	L��hϺ�~z$��SV�b��W��VeA�r��xE�恷�]}�������8Չ�mP���n��>�"vfL�˹U	�|��l���F�&^j���d���������ڊ6�`������7�w�����0����ܖ����)���Gw]���gMH�f���\��V�)��aI������V�:0;~MP���t�{��%"7K z�����І<�d�5�2�F�nǍK*�u��ݡSd[��'��7�!�U�E�Q��� lʪ�߽�s�ͻb�޿F�6�_�FM;td����g�*�mh�$a��T	��e�Nl5�$Q{��Zw�9Ը�:���� �1�9�~4�k�%�a��Ԟ2Kj.��@�Zr��g/�|����+�JJ�mW�HF�׍��R#e�	���N��u�������zL��u�V��t
�ӵ*F�B폊��Vcd�߷����"kiH����p7��P���5��Br�L��%�������.<먉*�M���́������l��L��"�&}�K�b�,�yES��d�Ci�@�ω�Zq�Ѫ�?�X�f�Q<��g��.k�c� طFK둤W�P#��e�p-�a�^�^��e`��x�'9��s��ۂ��r��+g���2c�1"Zh���ôp����C��p���*�v划R��yq^� �R�
����Ðc���^ɇG�^7����4L5��XvQ�u�U96�-���a�.��
�в��|��w0��k�$��
����`@2��%�c3�!��1<]}�qh�Q���aD{wu^�_{4��:�.�����%/6P<���[��.�}��c1�V�9rǰ{��p¦���[�y��`�����\�Ů�ʞ7��L�`2'����0?�2����(�#�B�(�B.��>�b�%��C"��_�%�Sn�I��4��J��9��H?����G��D�]P����D��>HS\�TQҔ�V�[�Ȥ�M�͍ ZSX,N��e-���s$��cF�F?*����z^c����NL��� n.c�|P�^����[��5��fmARd�n�&ߡ4V���RCQ9�f/ �b����9v��=ح��4���d��ֳ�%���3�َl�l ���n�BgdxVۤИ5�����D���zvqQ^��'g-Fg�����"��Ӫ�淽MV����S���&��S��}i9|!m>ī���;���,(YOX.E�I�2Lv_C�K�pn|`�kq؋�!�	Zޞ�ۮȸs��8S�疱�߇��y�?,�Q�O�v^mB3o�O�L�f��o�6�]�8�F
���T|1=�L���Z�ܕ/jV�������Jx�0�L|��
)=C�9B��׫�u;ɓ5�KW�PΎ^�L�4k�y�	MԂ��I�7_RͫBߎ,���2��Vd������	��쿏�����AB��*r�G#�m�����9��z���;��t׏�k7�4�.p"�����q	i�I	6N�yþ &v+�1 r���������_��󪸠�8�#���eY�61g�{>Μ 5׳8��<WEH��jU����6�%/E�.x��p,��Y��7�^)�+��E�2������6��[~K:���?�m�xs�4�W�$��cX�������W
�?6����Ӗ|���7ٟ��P�Q�MGg�2pxu�«�bP�`W��>�]�N��5aͷ%�D���nt4`��*������;�N"���Ƴ�W�E	��kZ�5�~���j�7M(�����;����sXO��1r�`��FǠǺ��-Tq�(�T�ճ�|~�e��.uo�
5?��2V� �J>g�p =�p�h#�#ٗM=ln��7EV�ǁ�ذ�(}��I�c��PS:Z�W����x�ʿe�a��ў+�h��~�I#o\A�X����"2<w�D�#=�@P��B0�H�/��T:m}ޱН�x�y���0�=ms��J��-,a$�r�es���oS�@���tc�\����]��9��D���f��D�;�n)џb�-�#��}ɥ&���J#j{$��[)_�w��.	�Q�0ͬP%��[�\_.c�����m}L:�[�2\uŋ�(����\T��,��|\�A�B	w��Plb���tX<<��28h	�LQ��e�s{�M^CS��h�.SG�,��<>��x�BEι�㨚�)[��cU/��[J��Uj�`�A 
_�z˶|?�&!���z��˷S{%@[0��r�������a����Z։I\Zf����X��TY��j�#є�:Q9b�K~a�t][���z�3��k��:_m8gP�����Lbd�o-�jm8)0%>���Dڗ��~)y�?1`Y��.�Gt���n�m�LV7��*��Drj�(���F��S7������o��T�U�(8��⾅6��-.�
�7���h->�v���u��z���<$㜵�.K��2�j��p�>0)�⁗6F+1�"�n�82 |�m�ZR$���w�Y�f�?^ �M�y%�[/$�Y���ZL+c�J��t��AP�?7E����%��W�ɘ�����߲D� P7�����u7QQy�C� z�-��W���RU�´��!	eؾD���t�ҩ+� ��[D�� 5>BG�ҝ�d&�-�l�˧ ˳�=9">,�b$;�W�����_��:<���[x�I��k�O��Z ں�aw%k����b8,:�#��4���S2�<�����P�*�XL��	e� ��:]��^&��=�|�����T8������\�=:��	��مw$�����SQ������J���w+��$l��}����p8�>���觤�^ �~��^ n��bpԔ��JER	��� 8�����5�W�w]��C^�`��,sN��Y3�u�bDT����Ű�Y��@��J��BI�) 9w�°�[�@�~��P�E�:k��u����S��r��m��y�<�����7XQ0#�B�)��V��If�)�p0"k{��p��s#�ϘZ:��1Ov�|���j�N�=�wh5'<� �f��PFZS
tͽ� (�t%�� ����'_�� ����q��$�Z�],� W����{�ﹿ�O7@�Ɔ�f�`8\Lw�J���hyzc������&�`R�V#c�6�,��`��[=u��Ąf)X ��E+�7_�{������y�=a�
��e�Ơ
�	3؃��{'S%#�&�D$�ݨ�+N�\$
N�����nRR�õ%D��Ca�}CZ��+ߕ�ޏ���6\� J����I�����(1G�;��)�rJ[�~	�
_������ɾ���0��r;{+<gݕ���l���x-�2c&�[nvf,�t��F(� w����������u�O7�nl��0EUZ�z�8�r?&~�AT �H[)�X���m�e_�^���Q%|�L3#�=�1RZΎ�?������jS;�1������C�-�M{Mg�CR�ax���z�4�*½�J��'LT${��k�:a�Wa�����j�\u�����o�2��xߢ@x�W.�G�'y��y!\s�ۡ;q���=l{�I�2K���+H�F��^S��0�<�-��2F�v2U�{�޾�jO�Y�}D��?nF�e<.�{�f�O㒤]&��1Tm�%�ꤸq7a�z�W��ԇе�z�^L���_μ�y<���[c.�9j���Y���m�YЖ�E] ��]�������w�iI��~��a��b��=�V�0�*0a
]vE=1����=r�m�8Z/�;��,�Q�V���;�^׋���éF����n�6ӯ�Z�1�3,]^D�Wv9�����|`�Ӕ��:�Ux���wW� l� ��jy�f����o�E�SP���(#4'Y�-d��Pc�7�E[T��MɵLLy �-��:��i�٪H��h-#wi��%��@�L���7�����MA��w~��7��B[/�:�Sg�?x�p[)�U�G�us>g@�wc}��Ί�����ի� �B�1\� YAR�=�����G�΅hRE[=oΓ�e�Jh�ǜV�\Ϊ�"��B�%���f��&�P{�5߷��,]�,�J0�Cq2a�Ս��W�1�ܜ���K^5�Q	'=|]Z�����W��v�T��{����ŷj�1.�n���Ƴ@�z���Y�F� �#���i�dal���*��{�O�0r����L<��ԓ�WL�TRy;����\2Iw]�>;1�Y�|���QH11{��	�bW�����}+ۣ	y�B�C���1����� p���k?��L!��-�}�!��Lof�����u�,N�qi�'Ǎ��(���
'�����Smt,�����QsK��(rZ�]Q�[�E�>�>���2�h�ԫK#����ښE�.s�
�4+��y*)/I�S�iT;= �i�R��"�`B���A���(̆L�]��Py7�j"��$�|������R�Yb'63ƾh`��@���XP�H����(�T�6������a�Mv�L�n�2��g����l{���� ٛ���
�e�-�c�������2g
��#F���z��Q�!S����u��ɑիS *��&'��ř�I0ӕ�}� Rf��8��a~��9�C�~O(��w	V>1�s��� ovC�Ǒ�K�"F���~J%_�"��� L�R��iWi@�-���a7@eq	'�etGe�R`�����z��;_R	id�2۴P� ��R_ϥ߰�)�h��y!9*z
m�(�g�'���s1�x�DE!�,�8s��=I}o����1�����DT��޽
���zt4vwWn�'���9 ��X�%��"�;�o���K���
�!Z/F`����U�����7!��:V�!���݌4i��|����G��A�O~NM���O���G]��?��F�N���
��r@�V�b��h��3��}y6�0g���Xm�~R!�����	,9�����w�0�*�O�� h�a��o�+"	�W��d��O�X����2�p�訟���;ux�y�S�����R��]��g6B�_2��T�,�"g���t1Y�ZsO������C>'�ɚt�Un��[F�,��&T�@��-s1O�8\�׼��Zuɦ�\�+�\�⪔����>����'{x��x;� _ɚ�k���MKA��]z�/���l xA��c����I� x���O���<��+���p{�tW�G�mI��J �zvv����B�H��I���^��������
<���W�R�߻��p�C�֢ ݫ��ϖo�� A�.[O� :$����uZv���D)k��kwٶZ?�#�X� c�r��Y��1P���}��F���:��L�Tw�h<�����MC��.2-�����U�,����J���f����~�h~�?��؇���+z��H�B	�Ŧ��}E=��P�RM��=J�%��'��=�5-��J�n0�k�8{���\�ud���̞d.�E��m����e?�.$ 7ټ���>�)�Hm
qh�~�_7n-�l�w�hi&�g�Sb�Q�ЬP����d';��o�Q���X�R^t1��P�ȋGA��D{*�B]Rq�r�
"sG��_@?��]ܱS��/���H��|x%�c�4���&0;1n���z���e/º��w��Y���;�6�zM�o/��;~{La��f����P���f�� �?ߪ�/j��2���< 8���Ij@ f'	�ۧ��t�!8lZy��$mhgf���<b\���?����{b��#��9�S�^Lt��,�*��	>�籠���rƖ,����|�ЎB� h�!`�%��-�?���$���z�\k�E�=k�zx�d(9k����#TX�!�u�
��ɄU�>����B�1WԼ�Mj�q�J�#hw�2]	_VC��,�plw�� q�8��]<����@)y�@VQ�ȑ}t���0����;���<�d� �2P4	:k5�^�n�v�ݹ��"GN���� �O��n9*�d7_��=��F����X�+��v�\[#�TB���T�L03G����F�u���>>x�C4�HŞ��S ��]"�*�:�-D���0���L�7��x{U���
Z��5 h��s�)W��r�#D�t����h�2p���������;{d�E�x���A���!�;C��%����v��O�G�y:��lC���^�j�A$)܊�@>��9��R���p��Pnx��R}��0
�åA.����a
�����ȳ���m��@��[�]�u��w��. 6�i�6���A�.�=e\���ӌ�}&�< ��Ni�����t_A��ð�m0����@4������&��'�,��� �Smh��*�DzpM�e��
�G��`4h�%.l��q=  =v`�$���)چ��?�[��s�D+�0��H>����� (��� �U���;#��~�e����| ����Q���vL)\]j{�#��x,9��L=������	ä��{����w��Ci�����r��e5��k���;R�(�7��7/�̳�#u����P� �kq,㼝s��\B�����Gx\�5 �?2l2�L��֨P�1쮓Z�9c�lM�q�a)cE��r�;�M���le�F*e0i�,���=��1�+qϕ\�B/j;z��r�p+܄�A�O[-g!�2��!.�FB��L����mЎ���h�f�q�cց<��s��/����#Y6�D�-�Zw�8 L���x�cːL�)��)��2�-�.���'�E����ݣGlO���TD؁g֘S��1л
��qf�U��[O3�*4��4�+4N"|�L2瀥��L�l4#����_���AJq��1$�^k��D��1��G����`��:���1i���o�ِi���-�c��@���R!d��*��w�V�ك���܀a����/��`��-ꩾ���<HL* _­�j��u3���#
��F�]Pԏ�2��U�.����;�-Ĭ��4JH�������>$i\�5	�F�}��د��ZfaC-���a��ȢD"�nN�0���NWA�����O�G�Ԙ\M�K���Tv֓�#�٘�`�V����/sm�4Z�mK۲�7ɳ��S�w%ZI
������O�!
�J��Q�>��������ի�>��"������u0jd�j��v�=�{[[��I�zN���j����t�D5!Q ��h������W?L�(<��G�.��\��Y�M�ЮR����F�di�%�"p��5I�*�.P�1A���a�qК ��&	�Bi:��i����OI�a�:�z��g��v�����ե@�Z���%'�q��{d}�\ h�<�0Y#���XEm�����fbqy�;�0*���-�����m�iP�+��װf�:F����9a��RZQ\�jn� K���!����+bNs��f�I��dì�B�Z<8�!�h��(O���y��t���~ig�n��2�����ŧ�XE�����kA#�Or�9�Ϋ}%z��6�{�� �<B�{8�K���6n2�bg'[6�2okU�� [r��^���e��z,]l�i��u�V*(b��=�[�L�^)��[6�����+{`ޤX4ۻ���`��L'�E�U��3�1%����=E�$�PI.�z���%���תB�z���3��~&��S����?��O��I��Cc{�Z��r�=e+��cj0��u���ܹ9):�񧨃��CI*������GF�в��&�[�O*-(#�8\�4E��Xi}R���k��-���[5*���uQN�F�~ĥϩ߰��V��5F��5��rAGt�`�|��q�&�i?Sٛ�����u�����nUd{��p�I0_�c��)b��1}$_}i3�t��&B�*���ΪL06����h�sy��H�����}������SoS����6�c���,'QG#��1汋Ņ���{�f^ �lRp� � '4��y���T`R�b�|z���Y+DP�D��-�g2�-��㢑�mOr���Y�aa���F6MQ|mZ�/cΕ�fe��m&>w5��AI��"U�%��
	�Dx/�?�]�!���d֋�^�+���W:����VנuE0b_ʏ$��Ү�����8e�Waܾ��0����FÜUt�x3�e8�n�<�D�K�V_�H� >�9��Z�L��A����"#�{����		��z��W6܎v$W��Ƅ�����	׮ݠ'�x#�:�D/3���&C��=M�L+�{(�́o� ,Q�	&���?�{��4�^ZP�4���Z t�;�RšPZ*t��Cp���f��Mg�:s��œ���)^��U��i�R����W+7�ٷ��=v
�ip��f_�)MC���PB�zלߘ��&��<��Tp�>�Et���A;�T
���9��u�SG�T5V-xj(
W���Z���1�sCx@5&J�I3x��}���D��q%I�J�j��b�vx��E��L��I�����"7,G��������&��hk݃MI��P=�Nw�o<���L%�=a�OZ܎�*���6�Kh��Q(�|Ċ�yV��nւ�b���5�Y=Ѱ�m4����}���d���-����-��J�8B�\�J���~�˪�Lk��� ��u��6���Vk��Ee��B�)���с�,����.ј���cF��k/��/��=1�m�p(7О�pVB��A&B�gKP�#��:\587����&u���w0A@��~K
�$���L&K=�/P�V\9ߴǨ�rg���)qKm���3�4�` �ʖ3ks�_S@ܞo �����b^
�u��jy�؏Ko3Vl@VKp�lO�!6֝����ϧ�n�vfE����v	'�3]2$q����²�,���kq�/��n<[�\ս����������,��,t[K��_�p��#�J9�V���6L��'��EӶ��ޖ[^�uvc��L(7�Gc�<�c/}S�j����!<��&���Qg0I����@� E
�p'$*�h�ί�*�<� �6K�����VLv���4��R�EjA�,g��G���mg����i�.RT�z��y�ęf��'��*V)��mʸ�M7E 6��.�9����lP�M��/�������u����ѓ�Ϯ�KOa�5��m	�8��+���cJ�������,z8m���\%�T��ܑ��
|��`E�FJ1l9�_����J�in�����{��6�w f|İH<q�k���E������
�B:Oģ��n�E�-�����aKy��>��5?f����X���B�2;�(� C"]h�iTp�n��vZO)�}�hDWFs|� $����z�nnSWkYXe�	Kb�[
���O�i	&�7Xn�L��#<mN&���79��ɍ;x̶����ꔃa�(%���B�cR��W�A�ܜ%L���yI�^��D�R�Ѵw�Fa%����r�k�]�=G�]~?�k_n˞�a�D�<,�;���!Q�]`��3zx�W�������Qx�F=	���P���/�<�K�a�ka s�ih��_��|�����n��R��8_��L��5㭞�/`vxL��t����mG��N���HnJ��*�O?$L�ށ� ��WR�L�OY�f��3��{e0���'�^O�*�G2��@$_!�0�)Ns5�`����:��.�3��5ew5�zS��㾟R���tio2��'������z#����91`K�H��-RNji��R�#��؈���-|�xYa��ՈC�@����% ���їq/P��*RF��N�Mm�S����٨X^y��ǐ-����lݽ��ڻY]%VMG����+��v���vw��Y�Џ���iF��\�{�gf��E ���	���e��|o�/"��8�����W���ھ�X��es�HV��s�?�����K�e�M�(��&�R���]��;|��Ǐ'*�p|/+`�����z���A��}��33e�8���m���d��`f���IHg�T2�����Y*�� �����H1�z�4��ԝA��"}���j�N\DPpa�*>�|�ܕuF��(����/"�Q�,��@�x{8a�D O[Q���=���x�!f���C�H܌9�4�ub��=����x$��@4ѻ �|��j�I���6�ǒHp�~�.]c|snk���w��
Zs�,$m���|�Ľ_7�L9x�
�A*��n��XH���l��i?)��� �)��mNG���n�:���[>�������,�@�>�F�RuFd k��"�yW�X��>P
9�gl�͏��5%��k���o���R�'�-��:�'Y� ��Z�/��fBS���.�^MW?)Z��
\0�#��<������^mt1�.W������	l: bҊ��cۍ;=V���</�D]��I~� �/D�@����R�۳.���X����&���l�(��DY��[�V+<��C~����Th8�-H� -mbn����%s�B��L��M��"Ql&L��	��
$�w�ZF�A��_� �b@z4�g��VF,҂������2�~����~*�(�fť��?��/�����x��˿R����:<li�_��P2�����egb;�;��|�x���;B�GT"Ә��{�R1��(�Ni���(5���e���Y�J^�b��YK]�����uz�G|��3y=ԙ��A�RsiB�
�ڽ����?m��Ɠ�1j���T&ݻ⸩ m����E�����v8����f���ː%UƜ�	��+|k^�<����r��'�D����y 	b�9U�
��!\��+_K@�]xƜ�-A�.(���ă����N��Q�i�8�Ё���!�8µ��r���j���1�ȡ
�=(�:k�r�+pi������;���/r�rQ&%X j���3��8��ۿ)�,���ˆ���'K�f�H��4�(�J ���!k�����߸��o7OͰ<�쉥I��@���_.��G�g�i������H�b�����Ix�ؓ�7��)/1
��v��9�a�1��i��+e�`nq%�u��Ű�*y���y\K����;'�ceO�����{詺;�|���.�7�#�Z�zXLª�&�n�&{���a�\PF�P���5�^;� f�"�(�BϤ�:wہ���q.	��-�W��*/J�T�b0��E^�.)kW7�H��y`��l�Ԙ�W��ǟ���Je���N�vo!d���k�UT�N^���*N�H�щ�����da����7"D9��J��9�Kӗ5��E��n�<G��5������^$m���b�����d˽�M���/�u�HE��!�?�b{Q�#���z8�-vNA)�s��B��
��ʕz�ٝȺ�!��Ek�.�㯔F�,��?$jq�ZK��i���I�c��,f�u��!O���2�<ދS�0��=�#oW���PE��dn�윎��6(��[�L �ٴek3R�˗�q�Hj�8�}���y�&��}e��9�qC-�L2���ӌ�,?k��.��Z�����}
�E=y+j��qn�&&�܄�J��/ުBr�QP����u0����#?��X�>�!5����%�]��x��RB?�X��A��T�75���`տy��%)�h�K9��ig�V�b~5P9Ov�K�A��u�2�<��pO�%��{<@a{���F�4i���s������w�-J�b_�V��d_q��)�-G��Dc���#������3�D{N8a�D�-���G|�p-����Z����7y��Ls���}P��?L���,�  > ��p�4<Gt*�v[!���QAޡ居ޣ���1o�' ���w�a�yc�K���W��H)�����b#�C%��e�3���H�a_��F\�t��Ɛ�!{w���*���XQ_���#�0qO֜�8�J��k%�ʈ*���`�{�&��D��DܿÙ4[��8��,d��Fa;��Ͼ�=-@�t�$�1�&�tըiH2{'��A��(a��hnqT*t��0zjƱ�Y`lž�L��X����$�Aȧ�
_��4�}�%�B@L��2;�2�m��G߇��urߟz�!���G1�;�WA6�\�Sv����>hx+ jb�l��=��.v�a�r~C^3AA%F�^��X�S���r㪆��ebV�*,O���P�(�����ը-T��{;�0������j���Iѽ4���^����F0&�%R�}IsSЉ%�Ztm�L�EJk+�#�g O*�`	��g��z��c�X�*���H�{���O,�]u���|#�eK�@��lm��F���*�7<N�XJH���;g����t���K�iXT�={�T�ޯ�������,����=Z�64uб���Пqj��<����*Q>��rN����:�6=����Z�A�$6+�F�XPu��8�o���x��_ Q�+��J�M����p�A�|��e_�s�M�-E:��~A�F��S�m߈��j��E�\�;}��XI�\,�� ��d���=`ԧV��T_>�d�4\���&w �@h"��y�c�.��}��*�k�J�t7�C���[�	Έx����L�´+i� K{��Y���^ل�f�f����~�N�S��S_�k1k���7�S�Ƕ�/;u#Y���db��Z�c�啵��ϥJ���yn��դh�5.{�����^��y���!|xxr�8��|�MN���á޶9B&�lϣlf��r������q�&�.�F�u0A@pT�ߙ��{x\⑰0F6c�Ǐ�c�)ޯ��6;�� c⫼9�_��i�I#�n���.��(綛>Ju���c2߀���{������e��N���`Ñ��'8��ހD79D�v2Ym�zި]K7j=z��|�&{�B�Df# )�̴���o��SnZ����g�\0���QVߣ�At�jD�l8��خ�9�c������2+�|��\��E���?��v��(�H��As4/nV�b�X���ȇp���dFk�9�W��e�-�������S���ćz�b� �Ϡ;C*i!/���<�p ��n/�^~����u�θ��70��1��{�Rg�K�!��Y���e.i`�Կ�ƋLc���ƼL�2p��14���H]&�,�S��N�ȃ���26׶;�٬���u0W�X+��(�0��#K�1����xW��]G	�o�!�m̽v�����t�Lb�e�����kW%�m"�	~�*��x_�� �O,RW3�7hB?���P�1s}�CTB~����n�MrZ����"���c�a���Z�)��˷M*��K�=�_��j�7����J�Vr?,��O��\�m���qJ�>f�]�b'��3I���I��s�"��-�T��~�����Z����ZL�wu�c��
��D�������z������7Dv��Z�!~(�:���r6æ�*8�t�$���+��=�\M!�CT�U�WT�$��Є��8��rq�4rȮn5)�f�Y�f�GhZ~g���Y�,>�$g�<j5���m�		�(�:�/$�N3#��\���4-��S�1�ŭ��:��-�09!-�;�V+���#X�~�n��~���yd���\۸�VPJoop���qz%��p�L��2l�8�{lE3�T�����xY�+ʀ���5D֟���;m
�)��'ǒ�i��̥p��Dr� PF�4|��5�P�hwu!t��L�1j|Q��T�1��'�14%�ͭ�H��_鯭�h4[	���jUu�s�r�N��R,t�m�	��z#�t��^&�����!@���g��w+�<`��aQ�*�o)���5�s[����4�kb���v�$U�{�:q���F�
)]u��,0g��c�%����}���iC^�%Ȭ"肵C�;ͩ��B��=�ɞ��p���ڔ��y�뻁'�O���G��o��~�ڜ2拃^#�4bp������9y�V�EZ�=�T�@S,��
�%Q�"0dv���XH��H�\�ww�dCIA��	���Oз.���?�M�M4_���Y_6�8�Ekq���&aM�I��_.  ��0��tHCǠ*�ȕKI!k3�cr���� [<�|�/�g'��O�Z���7� �������:�����%C1�)4/V��R5N�"���Ց����������F�˯�����,�9kD��rH��Xg�����>��;m�>����T҉���ÿ�M[U�ī%��Z��gT�(w�.��};�o����v8gX.���D���pD&�#X\>�Y�n4ǚ9#�݅��} �%��L�pF�}i����cNUJR�vP�5n�鋋��E8�<�� D
�<�e���}Sb�a��S꧀f�-%���k"zz@	�_�.|�Z{<�d:m����I c�l������Ju�U���i��>bc+��s#0oTF�la:���)���.���^���G6p�����Zc_��9�(z�xa��{���T�����˪�"-�t�;����>?BВ:8&(���Ø�Z��AJi9�Qk���Yf��� c{�u�I�~hӄm��ڷ@�s�ӡ�"M�RV��;F1|E/e<^�T�LFg�䔾6J��ʏW��b�+L�¼άdk�[P ��
ڝn\q|��ϓ띗1
��Q7�L�-��v�B�S�>C�Z䠗�K�w}���4�.2r���
T~pq��;8�Q1����r�6�	����c�ո�(� �6��`��+�x���,�-}9[rz0v��5~G