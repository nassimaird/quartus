`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tzx32CzqVreTaBGymZjd4F51eCfDairVsCQHZJqx+c+y7MT5wTY9fOEWdYhmlfGv
5X/HBiZ8ZIrbpWqXOeFP8pfGaJVw2BC28ZcPcAT9Nb9IK5qQCgzhI6P7IYZjQifJ
USQjYUFeuSjjAOkAqOAN2GJIHKWQSg7EohBGKkVuRQM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6784)
VlBmFcYNWZSPiEOcU9YFphM1KhI0J8fWGLATT5k8Q8GgsJ9g7rTCUaOw+nHPTm47
JnIvu39uTzLDgNiiSMJwjQ7tNz5Z99wLDxA8mmL5KSSxTXjY1JdeuXD9Jl+e0mig
5pCQh6BOXiINDv09BJgXcKEROBnQI4qZGEiNQvCUbx5swc3PbTXaxlEb/EGVHJ7q
6HN0e2UKddHcLMSsAvTD0xbgwA/aVBGDhNMFD3ZOK5W2K4E/uozJrOZIIj5ptEnE
QS0D/H7RwnWCzsrHPr87Koy3KAylHyJpIptMVEa+99sIKfW6xdxANfUU7Fp72NrA
lsoXwoWRXK1zyY790zmT8g5YBhgVUYgAl89+8TT62OlFPUW43ktB3TOiC2JvYsSq
fqokPbGdrnn89IwBS2UNdVdiR0ewwssqKbTBV8otxRg5qwjtYBHX7CEOn2EFaQ2t
i14PzHisfu0ykRmGd7vbAak2xLRdldYAm/fN9tTHBpD0KCkpn+I75RNYehHaXGU+
gfdp02eCWFRBwWBJPi9n6EEYyx/oaK8+OZRQFeizsdMEpNMMEeBpKYX9oe5PYRLN
J3bhKfNRo6KWlAAo7eY2m39m+OV6Bs8iPZVgykrzg5ApQEtJ3pu9efbP2Syvyflb
0/aw3kuwpX8tz29Qx62sx+c+Y2Lm4F7hqsRtw3e9LrNdThdJXsG48/fvqvvImBoq
7BL83gjWdWzzbDa73pSjnI2XJH8DmeqEz4z6LBL/l+lnfa8DXySirEJ1hURojsci
HAsh04S4dEy5UTJbsZLD4ElknBZqmUQEW3L55Wo+SSdXsJ2FTatmVwPR7Vp7mSA4
FhmaT8I3AtqI4eqaBtAYIyeBSwLcFgFPc1DHVJ7PGuLnJkSCQwZyA8sLGxfv4YDt
SbMdzg/4SIVkrqELG8x87g89++E9NW38LxZkHsOyJxgMZnuFwOSNqWTiYESvon8N
BVn7CC0CP5FJysIaOlxCnM/wqjxc4csFHydg3MBx0c9bm5/iPaDws6qz1FR7Ht4n
e1l3RLH3yizFc01APNpiOw1LlaAbvjo2mcJ/Nfp/RTZ7fEGtfVFzomuBSVENcXh8
dCneZEqMfH/bB4bZmyvBKrvF3tJlUqLGLnVPXlt/RWCfDiwvae3hfD16e+UtY9+w
SYtCN/lkfxdIjGS70bttm4CL90p7fuHES2wZlR0NK60C2ilisX1OWGQgGCtHLDSp
87gXzQYsr7m//A1tOcPuee6JJFhXPSftHQU3dmANI0hJ3BE2n+DmeYZEqCRbg9Z9
pW51gu0FfMOSVkqpMcwF+aT4U2eno7KLl+wz2LvD9uRP1adqJ4ZkidDjPYjmS1QU
EXzNFBrx27ht45MMEOT4a6YkfjYrE9TrQDt3fJJ8hmdS33ZsgJ0xnh94dhw0Ine/
AGPzwh3cZMnJVwhQ+S4v+JVcdXe3Zv1Xe54KMLdNVot2DkVxJmQ8G++1jh4S3dUf
RrX9JEL9JqorWIQFpPWuf2Czxk2dmRrt2LHSJvkeuJQtCspFFHhH0mOMQD5JqF3P
gvhENNnu1sqFkPr4b52CeofGu7tdDgST5/eLYch7MfHch9zevM++rMBWu/i9upB+
P+4mZfDCbQj3sc3JDkZU4CqN3GOTaBTlTMFXOUD0rsd+SRd45YIvNrWN2AK1OhsE
6SlpZ8hVLklTgaS4uy4i9lvG5vnbK9oxqFyZpfkoz6biEBgj/gg+H95reEXb9DTR
fVRWjZJkNcLzFvNdHj0WlOima/LeqL1iDYpd89OISzIkgupeChQHiM7hWqXDZp+C
HBgT1oYi+P7pw3jM1/HnoVtAQnIkCOMMnJJ0ZSWnvLhKoX3sP7D1QbIBTQERlR/5
vqdQ33IlR9yLhPCaYVjGiP3koQnydS+X/fwXlNnw5+8obnJRscXyi2ZG3FTEO9EX
/rvX16MWClGpS9/fLUZEaWNz66N3GFpoNxxdNijhWyDaaSRL0RERuiO7magsnj9r
LQ/EndNQwdanVgZKVPE6Xni2Hru/a/+lFuJPOvYRLD7xWXJwNKprzY+Nkdy8Nl9x
8nmhlqhfv6Z9gk76UCWKh4n9tfMrzYrmsEHrASZp7jLicGqKln1qe7DTZGWYX0yk
z3i9wndQDSNAgSDz3glrISnJcyPhGrCq+Dmd9LBL2ShjBuBcajhbHKRPy5DrC3DC
uvhTUA0piVVna9yZzS7fM8/igM8R4+/4RdDpMwWNpA6yh4CuNQ3oaNbRKkon0niX
DGbRM4VNod7lNn/sp60Hlypqn5R7KHoBKk6SlYJlmnRuYhd9T0gDJ6mQdwoQ99gQ
kWz4XDV/0RUU+rZF4tmlcP32dEcIcvBMRgA7D6SO3xHl8mjN+TvEr2m7WxZRVO4+
FZ+i4GHjVZMJi7DZiqxiezoTAFmu2DyKsWmGp54nwacN2JcIRo8bC/kqOPYshwY4
eGtrEtoOrYhsNCvFkXhC8JCJbeJ87wWFiDEpUgj/t16VF9Ke/FbBnRW0vR/p3DrG
lVWZt9RDGFVjmGkIfv0IAAvjTL3T8WPPVkKA1TQJR49auuiKOD6pXQfTRbecpGB5
z9olkdqxAqn9+C3EF1PKG/4asDfdWwimE/xvKpHpMpKqeMKBJ7+TVNBur53WI04g
QiCyn4/bmAw/CkK7DuegKdeI7iXErU8hs/x4BgdKdBlTtkdLZ1yDmdHMa6ZJgR9Q
y0VejlQO9ZMwPTYB43wqJB9r+fYF1/n4AxZKpYgQu3aF4pzyhxzm96xiaESmJILT
TY1l/MAT50XXOvTn1bWbDRiodBDlMWh9QkuN5ph9QlqqC/pP3c6wiGJrGYocmSU6
viBs9fh0ISTeMXZwwdqrnu5FLlJoaS+6gwHyYWMWqfQUg7qM5yn99EdNtHxPHaTK
EquphPGIa7i3bdFZ6Y0YuSVRDGPii8wzBuDhFGIpKSG1v4FXcWtwbkNjyIVkeAXO
noBo1H37mvv6qvCpaDiPKsAuouMs9Q5sHv8Hn4rVRWs5nyweaDfXSm5S67cmEsAT
fk5er8NfPCQ+kUMqRgKKf3rpaA8q35YR/wmbGjnfn7d0GvB+V1cAt9+pbb3G/CQc
FrxFGl94D4/zG0wURaKEOjf1POnh8/YQB1RTHLkwFlswiFJh/Wpcb7ntsspQkRgL
wk1MZX8mpPyRysz7KaFLy0cq4++FJHkkRHUupKIZGxqrjdQz/En04NbzmS2hTvSc
YZuYELP+vayrcb6Ou8kfp3a1wxy0FQ4plk5l29AQVG0X6D62oANyJuqeoC3IfSHw
zSg0yp9ZenSG1RMC2E3ONIUVuRF3vfebU1SOAStkKGpwwmD/JaJKyQ6Qv6HZ4ZyX
J7lTWnNQvewIHVpVtxlv5OeZC6dP6940VgXw2PFGBrGKL+dbjarEwfl0SYjQAZPn
YMKTPWPQCOtmG/twAJdE6kO3uFHKyXjXaqj1iEyRNRwacP9PjNlxt62P8BQ2+PkI
yN/wZOJcFvZj/EaugjqqBFL2qHDwz3PPqoTO+9W/X0NffKsTOtxZjuKKIgmI8ZM+
AC5TqE5v0jqTN/4bGQfdh5uksXcAJs4i0KE7dYpj4bCGQid5RudGnreYSplbbCzL
KcxNkJQddsb2irviq4OsKlgcOi68XFvSF00a0Fbx6RPqzWLafG2swDGWg/dNb/7v
8ZUJzG0PZSeZJGSllOfr9mK6xaeJUpI7syvz7CLOdfwjtnGvXAkcxIJOpYbG74QC
h/YxJSW9qcng5/TeMx6Jkt5SSNIkzSiZS9DYItc+MFXHpJRLPLyn+DbmLN3kF4/H
vcuMa4DSlKm5ncEUacBXacVxLh6a23RAiRgpG3y+tJiW1kJrDQUhJRo+ZCDyGwWR
BWSdTFt6DO6uGqhbz8iID9aC8hSCcILnJtVmC43suX/EaiX82GzeGlaq52gPfRox
ClAzvxssdXEZ89vnjM/Gl4yPEDwmPeQV2ccQMRwlpRoLGoxKZBIqGuV8gz3IMthY
QLDWY68cYGjwv2Eqaj6VxOoEnlS5Y34M8IHjaLa9AElUj9h2KDVnschWQs/V+lfj
FYtQkqp2BOxG5AOfURnXJnG39zjB7Moigb5hLY0flwc0PEI/LXhhFzCkiXi9cF6g
HBDFACVOEYlyMOS2v6gel6wOGBrxs5iuzM9er9AmFRB3iq+fbx/MVsBo3H29nJ9J
rnomstxSWLxi0USQhWSZc0KwTGL09PIpTWxGIjUD74wAZnUFrGFIYmhrCp/NbXuY
dUvMCQL+k3tlk0m5tolDWmskRGDlvA9N8l8QzqU4Vn2Ple/UZSwxgm5XREV9E1NO
duc8wDQzCDkBGQIro3MqaqhkKg3Pu4rSNlu1L6GpSHH24n+tdAzt2+hkRRll4sNw
HVfRMCsMy7t1paaUMTghkUKlV6MvjYDYTpzaWMd4PjpXnyiklHWOSdnSI7mvFvhG
dZVy8mBOixHcH2jxgzKCf9fP7qgBti2XoI18iPyRNZSQvprSqKS83p9B7b7OyL9B
hTWSupGaYzkt6GwrNH61BQmQgrEz/uuYKMO+Nhey0KUKinVwvQq4Y1kCSiNJVr9W
63YRXHruicFFuyxGzcAmTJYZV0wqWDT0yHeMyh7+WDsk8TR+inQGvAReWUGX5Kft
O2DUALZ1eIe2p0R6Oqg+AJCbyR3xPN3w8DHDHoyqrgPyTHemQu8rMxL0iT3jPDrV
9rfCUuNmOHTaDGnuxHqlL8xkVbqauh2BL1PIoIn6Y47ZV4nEqzAwoPvX3It73tqu
JG/TxFMnAJMmuhdIiI1dIt88f5vYApATkHpf6NkeM46YFdKoIwcbIQmvwHJISNUH
4mloqA/43duXO5HUPfR+zKnkFddbi+jdx7qtshG9RivttVLC/dsAUZSVUwiH/x3y
bQZ4tlhg55LBRSAuyDcEBCNIJKyYnsUbtAwzFkAv5JC3tK3f7dmF/mRtGFH6aWSf
qFu1gbvOBMo5jePXfJGl2+Y0VC5Tg5zdzbpeFZy6AXSWO7BZ8KFenRKqdljWSR2u
jFRLIuEiaF5vfCpf1bLXUDBZOy2toJ52hPMFmVyKS6KFYAZ3qmqxg6MHn+A79ylb
8A2Na/mKfwLkx68PIVKsWemNUgrbPcJvCJQvek+M4s8NiaTecIxYKfEFxDNuK4+y
B9A/QLpZyCgf7w8Q/8mQms4MnGlqGzeMOUJmf1soxJZpM6dw4/x3mJq5uBRXnRcm
W6WnnT+1qbZAKxA19PDjEHo7X4kFVxsprwVi89MCJEdA1OgS4NUSyoETS/RJ+U/W
r7FiztG4dqENvSjwYGUYEmIigth1l8cHMyfz7OoAEk7jM38Xx0sLcbnqIfFF2Apw
3FQDSdFbFmfxRI2IuNQzQ3cl5rGgCxTR05+Q8iRBtNMiuGCvwhQv+C+gu51iE+8g
BuZTNbH+sGFsZ8YwZkouuFGjzUxDA+oeCOEACC2s916fV0kmLBmW+tuRVev9Ckba
CrJueAeNPULEvnUCrGQmL1I7e4OgG7OU24+ommrMDsR/Upl26lfSicmqcedq2jFc
PhuDMHYTZCOMderNP6QqSQKSHS86+gfrlT6PNCwzzj1vEnZQS6gsIY3lN44IB8y6
4AZw5trfzmRt1Rjq1MOFuD+4gjVEjdocAxDi2X42AKdgoHsyzeIHIyB8N73Ed74n
3yeQxvNH3HMuVYJS0jOhnuqe37oGf3UoYRspehcx3KAjAi2RJ2tiNQDXOL3Iy0kv
XBVFjJLec0SbVmGcDE4RioKFRSPAXkAPu+qCGY7Dmuprbc+hIAmUrUBRuw9/E91L
2O18FIKuvfQDnHwxxqczEn7O1ykjBwwVJARYbtLyh6eJgjQAlGBd0jzQZ0G1AI6D
pNd2ZVnuYXDLlRTgnOuW/rLSq9HLQU8hSKvdRTeepFQTnLx5QK+0kqgaCWspBRWA
siXLy4c12Zg4SR0JzK9xqHjZK0W4bfqgCy6ywnZCfZuxj+ZZYndZExumMf+vGK4T
70bw1aGNsWMMK54p2krprP115fa889256D42AhIALebQKIqsgI9ycN1QSiYmAvKk
VfxR0tWwiZJCkw2FYsZivHOQJB3OXa5JKcCGma8IlYle4SPrgZvAaNxMf+mQcM6w
LvZUq4B891J9lgHp0m5OGAxBCwuZ63Kp8PY4hHKdtvTyPiadNhysAsVC3Rmd9zPw
CvXle9qnB70O/Js4Lr4zL4M9MPKtIpm+83AD+x5iwgbbzFYXgjXyj/RP034HJLSZ
W30ZhQjUflYlrXI5N3JccrLkk4Sez3b99xr8fc4xxU5voaHDuvZyjH66IqtgXsf8
RDfbZL3Zp84HVaqyzvb38JT+nZ2xWgJJ/aFVgc1yDEolJ06IcwhOG+tsg3387Ps0
F1VAMihee5djcgYZ4I9i+SMzryLKZoqGsZ1+qYuq/jtxc7mGiVCfTuimQryiq/Df
Q2cufbiTVJ3hTCxRyF3ah/CcwIjZ+4h3Ke5+F6Gp9vEvi44NlaNj6U0QvVfATLXb
WlSuzzcKII4ouqfW+A8N58nms206/xVSJnrkG1VITqyrJE5wpzVsrGyVXpSfMHqK
JX2FOh5nKkX/c+yN4WjHpCXW1RmSoBQM8bK+CHNVMONzcVEIJQQJ9t2qnL897oua
zDVkiotkQuVjq1KfdC4wTSsEAhxdtDsfb/Zj+VSLmFOcqrYC2QLwS/p0rJcOZsur
pzgto21GTvR2XB+WYroVcFJTTu3VjVqnt8wkzd1YfhYFVXyCq4MO8UlfOJ+AilFd
HKIKYwPqUaOcFbcZJWXzyvZHZvr2lLwRSN0Y/B+TWss8BtdqLa0ccoAffF6VZ9Zk
B5WctUQFSjHH/Dqpt45WLGOgaPBm/08XfZqbPHUSFbcwz9mJy3FEAYC9tGkxuEf+
H2q9JBCD3xDz03zW6CTobMw5UqARzbtqT3frrz7NxWhno+UbeeGq+aSyF4wd6I+N
2PhzDk8/3RllHpMs9UaHejnkevLJ9J/1dEH9X058w6oCStkWfScwKlkHonar9Db2
dtNqTx1F+0pFhydVwLytrPGuXygiCxY5LOkZuvRwWR7HVHrvn2TLrDI1ryGnBjEZ
N4dh+FMZWcsdAaMtYFQyZfNxkLoPTn7wVZvMvkyVdsgjoUh6w4Z8lgjWDxjlQGXN
xOx/0wZ2xrpUqMFhR56lhfoKSTl+bZ9An6bXiT6ZEHYvo899SVCzlk3H6mGczQq9
ZB2jrmObh///THDCVgYC91A17o50d6GvxXMx4DTA1Qt8fjAI1KaR1etAg7Bb9ruE
CKsfPxfyhAB3ai2weDzaRCa5PRfTB6xloma9w4E471Lo68I86od8QiMRPc1sagmG
sdnThMH/cuwEsknZoFEy4HiWoJcavckpeFAyf3BxLIhojJ1gsMGszgB91ARH8hAu
cohctW/JkVh11SLA3EGU142oq3cFnf7nx57LE1FkZREIaYvWlhJSbDJ5pDubx0bp
7JM/mumk+z43N695AK0MRV+sp+bW5qvFO7dnxh0E7UB+qCUQ98j3tenMfYUY7yJ2
wlc+mF/fGk7E7DhAt7lFwZFmIaEG4k7mH1dn1KkHPtHDIOb3CcZmUfE6Bo0aYAUH
1HLiwMi3tMQVHONW5NO+tIMgAx/sCs+OtgkNMrY3acyFv/a0ntHQgscyND2A5A3N
Znwg0ksPoOF+GWpHDy+Z7GYC0sioaQRgO5cOzshFB03KjGTZS0nAf6TxvFPMeiI8
8h5lGIoCMjALArx55TqPYATfzSJVYwupOq/fHHPzk6+BwdXy8w1OJNg2erSR9NPb
Qoa7G/FZnqrZVdq5AEFZDTL05aiYYBCZyZCPtG3qfsoH8wG3mJEspeUAX4e5Ac4I
R/NZGiF9oKJM5GxZElUf9qN/mL3s5io33THsnpO9E4QsDEpJVMfNcgDNflqcyv1z
sPBRSoOoylwXHBr9+FH9Qgo0LEZg3ya5auUUZ5s/xU4S6D9WvObO9uvje8SSN1Za
qgK90QGZLsH/9sVEA5hj9g7Y8zxuA4yzL0xyxKbjpOhnmbreS/FWqypZRMRxWc4K
xF9RL3wTn20YD1clZ4Z6NBKt1EKUuQoKNwGM9YH/3gNtmV2HLg8Jm8D9hyF6KQcI
K1qXiZSzPidsC4bFKl5zz7QXr1fC2GzU1GqZaAxBILah5NYlisOIl+LyD2aaRsf/
Is9CdJAxnG2JA10yt8WRZma0aD0qCe9zk56sJQEKEMN/lg0s+EsLiS3i2h0ijrBZ
dtIbLvZjVHVQAdwS+4YVHkqqGn4IaBBpQbx7TfLKV/QxJ86MO7dlRE/g6J7SGIIL
ANFcRA6zoLX700tlVR8JB74nWxT6TzEwwZ9eDBphn1BTAN7i35/aDSAlsWEicxaR
E1xxD2X7dAKAtVN4g6PK8usvJbRifzDtV9uEZhPVosqar4fEoogTR6XVgQS0dAAO
mNW+l31jUhRpsbIhfE/T3Ip0zsN6iknPWAIF4xeag0DaAQmhTIHZGWcrz1uZaEKe
ZGvJINmhM055JI5ZyJp92Xxewz4Y6SxYjrYbI5oEhsjTnevnmdk4uoNJQZIIEE2+
nA5T0DfaUYy07w1lvFfqkbGxG1hC6fWy8rLwBGeppPZwoRPHlwbzxiDBs82e49gM
cZSOuS9YWBYnubv40RHEaklSCiGzxjQDl/Xf56NDZOFPukVYbSn7g0oGWq7I4FtU
vMe+9m4vxyni/9i0ToJgbW0ToMOoKxwU+ftX+fvXK7SU4HBhQSNehQqIynNtt+SX
1O4qPw7/TzOfC/uf75ieOYk1lMNRvmhEzncBa+L4mAa0Aad+Iau3ihrKkPxnRDF7
jZU2Tc7UuPDJEpFqJcMfESNbK98FtHfdf2FLKoP7BUkonu/up3rGoyZFC8Zcmw+U
1Daz96R6+3Xs+leSH5T1EoN3LMoylw0vp9XhuA3g19yyscF7UepWjCDc4psWWn7H
B9F4dtCZqY5G/Shy/gXEsStvdrYyFnqIgov+9LHWvmkUEvRzETmFQbFHfPtNRyR7
4HSZMQ1IOd/TZFQJRsPmHJt9K+Tbh+yUv7/e+opPsyaJH/3Dm5yHfndRntadClTR
RLF5mpgYgF65TI7zt2UJHg==
`pragma protect end_protected
