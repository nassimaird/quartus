`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZurojlXI2W1wrNllYIhkLmqW3rq8GtBoV3RYMR1yUR36NLGNtzQaMfxASCGoSU6q
/dm+w1GX8ZR6IdJiBu2E/qT2EDpqVwTlW/vORt8VF49kXABAvklO8ZKh4zi9ivaE
WuQT4Igvx8HrkpjFZx/ArYIlEYDfiB1GoHIZfYzyvXk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46768)
pbuL2UYfzjOb9nguAqLlcn9SuCRD0cuue6VTWYlMAvRWk78hOxfVntJDNX905Yhj
Puarvg5na+qsX5KXZheq9wj+JkekmoutFwa0peEBj2UEr6tSAWx1zF20K/rUVm7m
rAhCyDqIX/6geEC/Nd62W2zb+9/jmcdI3kujdRK+zsQWHyaIPPcCz2/k7wUw99Ke
vQmLrVfaimUPQGWNkqhQY0J35imBPIYEACf933VLxWHvCY6h/W2WPKLutIqQEgVb
xI2W79QLBZESjFjvrwnE3o186/ZGoT1gxr0ERgv4s6Xcg4SkMV0zAYyuDUE9fYXL
mqrqahNjqdakWVLm5Pq3oxbz14pcvK56TyIKJnRursVf+RtpCw8Xa9s5jns66UYX
ItS/4faJdc9+O1yGxgkOn6nezySDkRI67aSkcPNMrMsHm8OkkFD7hpDySjkzeVDm
i3iUKzLMA4+TxzbhY4CAXPzB67Tc0ZIcx3yME1NC3v+91N9jPDz9TqmubgRigdyK
GfyL+hFrlDF0Oeg9PC7ORFMaFbnuoifr+8iFvXQzWqF8RDUonEeq2DBJ/mUUc2un
ECNVhV53yO5YgNm5e+I1QkhvChBOfmLxOhGaqXCFMhrPE7zAt6KGfcCpD3OyDwi4
0U8+muJcpy6zoBuc1qI7SOoGljwpBOGeC6Vdk7nRvcNwvuS3X3uOcbTmdQOloSZI
IZdJNR6qdCRgRRHAVRMtFb9xQn1MfD+b7A5aqUEOtN99bJmuzsHvYgWwEZGDF5+q
Xiwg/dgtO0dLXVRc9WY9TEjNLqXZvm0VxpVos8H+sc7JN4UXRQIyw9zKnawXOx5K
HioM1PKss7U9WTnuf2hdu5voWA3oLcdcQo4ZF/EcuRjO/m1BpcxFkxvDAS5nGmTC
CC5DoekhZJflAHH147nvRrGZIl1MTAlZgi9W7/wOQVmA995PNs8u4cQROy4hevII
8IVjDRUPOMv4I4EYg/wfxQr/Jc/AzGlZ213Ok/CRsg9l6wx3uOhpeQJOySp7JfzK
AN5bzRldc07tp68MTtofLKdyalno6swX+JIb7g1hiHFct/+k+HTRxD3NDQBD03x1
V1Qn1XALJc+0QXvNCVFFbC9wVRcUopAn4WMvKjAQNnOJnhQ907h/FIvfifQGmG1e
dYdj3cvl5myN/xtFZ1BLzUfo1I+FxCf8E24T6+Fk3gwtAnecrkBjkPnWI1ZXRmYk
4wyve9OU3R7ArvHWlChx0bITcE5KvIGvX7c7tcoT4asfNH4Q2GZECysLiVaR9r1U
/GCyvapI+5OwtUNM797gYFdMtndb9h/e+sgKFleV4ShwSckUgUP5wxgkG0+t+x+M
Ql4p/lrd1eEAnGhGUDxz2tx0UMmnsYlzgpEgJp3PlBD8vCoJJZ3VmDzI1poALmCT
TKcs6fyp2wdNs5ehd0hA17CbJTZRJME7TiZwJhfBFbKrk+Hql0GXBKUAO8wffwnR
q1cYMVzWQMJ1EhSstacDQc3/UXNgQQNMpu6D+1k9/lwM4IZNkfRZKX/8SQkaZ1L/
/D8DoOsH5d8tHU1NyxxTTJfEnqkcR6ec3HwnXZLv0+x+BVmUvXcB41B1VLrT8f7A
n5qQo52IpeArttU0xemQ1vbLQJTsHFrmPqIdmdihhM0O6xfjB+t97R1fVV9AKDc6
EP3vTHbvgdkuY9Lo98ztlTAPxKEQKQk9DGrXDIo7gTnEfkiofZ7guVLbnXTu+ajP
cNDlUEiiRoGnYk6YHjRQP/jC5OLvtWGlC9bf+03qGw+8fa0xh/QJVT2us2mjcZ1h
Vep+oEgyxQ7zOfyfF0prTWVIB4UkA5SyuTsv2dSsup/d+epiwJm4lvY7BUFE1Azu
AaiiU0RQnXKb0kqFBIIwy8H8I8kzLvS0f9li5UeT/E91z4NNXfXV8/lod5yAP6Ys
rHsyu+a4wrhXC379gHDsVzv87H21Fq9IXT7VR+OtsG+MNXChB4TyvET9pUSL6I88
odZwU2ZywupokKGKSH+lnDTnPYbXCcPPLZvZSQYE3L9DP8C0IcXhmKw+4oPhZSQs
Q6LccJBC22losJnuhOzZTWmfZvazQLB0rSktC/if6zGSImfLmRk/WsHPoevD4IsN
pnGIng2+OiYh4oHnFPmieGgMNkWcy1JvfpBesdAutlniWEHKxqK2oS96PYsuaP5D
vlDh5SMH99EJOblExEDjuw+8Kj1IK0wUm7at5JjjmpvlUqlIWncQifGVbIht37CP
JOZdYDzhhsrEDLGPmX9z98sXvHd/iPXpy5B0WbQ05KyaQNrS1OKDxBL91Jqlmn5u
WRsMs4Fyea3vRBwVZgqCFvTqop/NFdfSP1xByRBm6P+/20NPABMsa3SJu+vWrGUQ
aeWkx24iMmQedkZXaiiJJ59Uz0fV9rXJndrlt4xBIx4H8KmvZvMNfvX8G4rtT0W+
ThMwlIPcjyBzN8OSd9yVSfxN//GBCyYt+EYbSPPjfaFI0lsisQegZy28C9LExF4F
i6V4Z5QZBC9w/JJV5Kx+DkLiAIumEJAdzNa45NDgltGKeURuhSvrhve8Tx8iqQMS
VHtUeY8f0F0TG4RV0fBRXdFJxM6QeeuQznFcVFPHV0I/3eTAUcLOf12kqd9XvgFp
PrgNq/fFIIo5NqGPecgrO/3F7MOzSBtv0Caqm0a/Ihn8zKKEdjzcddL5JPLgzqZx
g4EMOxK4jUdwHBd8O6UgMv1aHB4HFq8cEQg17YYtkwl8GOQHtreKjzlYBCUBVd0F
VyJas2GX2fmcmam0i7jXmtvZgPNLHl+aCU1b4fEFon3toAWzxZPAbAO42C4LOSdI
1H+zSX1ZeMaH5TwMSU64F1FxtbtwmS+G4ksdtDhWhNyAI+ztDksnNPQJEXb46jBN
bKajFz7UY02tN+VFPrLrEayA9Wfs9TEdsneyy2U20hkF7i8QtIXfKUNQbO8fb5J0
L9vPenpxzGoJGOuCX+1yDyV+9KoUTHDycIcwuJVEHHsJ7hIc9hKLmtRqQApwVtQx
Uz0kk2cQ1UsqZX92bcGrXo6ka95Y3SvaN3kaXCH4ldYBk+o0tMu+u1YRlWJlSSRi
df3ilQlR77Ge3YyqT0AxLzbGIFioYhGSghmdwSPUjzk3ZYa1SipY1sD6LpDNoWzq
2PKrkzYkQQFLmh4E+KKxCnRUc5Q3DNqj0rdAO/fWwI0MY9XSetsx91p+Oyosath+
LYEFehVaqkbtkbqNsw5Yx03mOsEUdyzNz2qqX7E2Tyfc/WphxDLN8Jj+/Ik60QK4
EXEOBayTf2UnXzw46PX6203t0HtrKAc8dbxv0/8dqwdCApwp/XF6Y8FAX2LX0t2g
03x0LMKaDMle8UQ+DA1gYM7KF05y/VcF3g0EKATOr1u2QALdNnFfLncv/A7n9SiU
tm3v1XFjdsvZfVK5PlPEH0ZruolT5rM8qiyF+W68P8Y54/6s1eXjmmAF/YmHbupu
HyfPWpUBGSQQWZz5VOhc4dSJM5IaH/Sc59uA5Ksjar8FyDSctKR0lJd9Za1G3uSb
PYWYpUaQoBWO0WlMWolvruZ2CD8tMMTrdkWbLpu8b4PT5+i9mlXw8oeQL6KHGoGg
daZSmytjufdERgZUo8L0/oQQwYYaTWeg0N981FmocZSF6QffvM9oIxeBsty76lrS
WvCFrtMMeBzA3p3qsc7F9CJPGayDwSZe/31ecP1P1GPQ2W9JR6duZ5mrWRmv9oYn
NXN6lk5/cDrWOs3FYY/UHf7+1PyqKGoXeZzHppAjGxDMjR3bo7sIL/2fMsQMEC7c
aV3VGj2ZU3/Zamql6YaIHf57yWNY7u9FgXh2zu9zwSYLCShw3Q1migdnggm2d1OF
Hge6QBZBQ/gvc8HTeSUtaZSmETOqeCKO0mhHoY8f0Vbsr1FI7fmKjkuFfS9KnoQU
XmtrfQ2AoixdBlGFA0KciAyplLwfpsKIOGftiJ04ze6jq1t2bPzG9NsbJqo9RuT5
Zcl64is1foEgYjCUNgEO7Eo3D0i2iP8TJQlLd1/CUaJSuMVhC3iAk00gI1rtYd3F
g4CmN3t7J8RZfwr9CjZZl/x9ts5tFbFJ8N2dqKbxXlTDAbmWY2YWvBT+Y2DgZjON
B68kA9yAbdX1zUYWLSInz3a4yNllCy0UtGGdvU9yNEyqsPLw78QAWHhh7Un+zaPz
YNaL1ht4tVu+aVIhoKKX4X8Sf2PK1oqxTh3p7Grt6B/uSxOQQNNOe65MPAqGpz5r
gwQwSzHimBk8jef2sbLIGtIC+8Jbz4q86BGhOZWY7Q3SbYBaVZ6525ZSsQ7OSsBm
5l7mnlDyI4WcCCrDqvZBFBiKzjZL3T7qD24S2B9AVkpKTHA7wGEidhvtZKMnpVlE
f8HLOL/nKAXRZSlz/3X60gVvigbKWrGgdQ2CDFL9rP9EK6fiC6GDGRM86VTMCowM
NCVNc74ldcQNJ1q34G9nxgzPB0JuoiDVKD+6cFxNXY8iYjbhrR1WP9EuuNGt0XmK
4HO27SHEOsZAiXbWlGfpyHP26boHymVp+lhVlCxCrKsoccx/4FaD3hU95IEg1N7L
XOFUdJY0wo79haJndsSBZal0vDzYIMV60g6MvfH5Eo3mA5VhBXKhRhmZlPjPVaLb
OtWl5y7qTYAcy/TT3DLsdg+AvQyztvM7PZ9Sb/hZkjLA1220S9CZwypB8HP3XDZ1
b06HfvKm31kahKtVuF/PWlhJ1c9z4HNfy0oHHaop+eDR8nRng2lso1L3rlAuzdYH
dQktPz/9TllFhuGo3B6gfUE7MoqpC4XRa3EMuECKpZnx1lYBnlnniHrLcBim8eKa
Na3+nchAKaG+6E6Tf/w+lRM6R8/cv/8FPU7za96OAeeYK0NVM/7MtgoRPi+VGuVw
56wnVKaAbQVjr+s93VUVIxAZPUBexBPPE+jEPYe2XbYHePSfnuqx996pLg8/P1mM
4sQ4XUVeGKkiNKw6Edfjx4fnQSw6MzfHimZz8gp13CL1TEwykYaUFTMbXDfNQOsR
tzO3Jmhb/jo1f7+iyxJjarB8mNn21z9s7HOYAz0ne/bP+QvxnlxEztqGoHneAUde
1VpNaMpsfEbjxJIyQi50dR5U4MkzWarb4OyHkDeTHxw1UPCDEiUWSAeIT9i5ohsU
yt3juw2kFzJoiF6TyJ8np6U34lPiXS6sKXsnV3yxBkNAoxY2scijwvvtYWTBRCu1
Wg52os/wcEiUT9cjMa75OK0aanlKtqI6W/ncjIdjcWZ5o+ZyjsN6QpBBjMy87fPo
1zBAPhQmfa7MF9eeQ7gpgM/C4X3WeyxwZLanJqkxzWva7cFjcy9l4KXcR/U3UX0Y
//hJQEQjfaTWcOfWlIzinz12A5za6BJhGQas0G/scUnqsh0w+9LCpTmJv0i78M5w
xs1eakvLrmYVEUCU/A9fUOh2SfrPj60/auAxxC1mYCVcxR3VpY/hFjF2bhhrda6a
GgobMGGnBk1GwXfYdmpUZfc5kxzZWjoU6Ya5VIR/JSCkSl2oXKNqnfjus01qnI4Q
TouTgFbsP8HtTX58A399DNM+0zFubriHT4sLgQ8lcDQ1W9HUNwT3gkw7NcEN1K4I
+5fzibMkQPRk29AZM5VS7mMzv6X8Ogc5l338ivDlHc8NZA5ycw8/xwpd1ZfWEN2V
eUzd+VDsR5CuvHXd1rPEGmEBl/ozxpx5VRAmphICq4CPhbTQHuh/+ibkge2N+8sq
ly/eCCyMSVD58UPLudcOtydLbpFq1rzMRHZS8+AeOVNTEp/XqRagqve2Q47+xg+J
guQzsyFbQD39bf3B8XtOr8lULlzo/BfJ25MjsRiQL1JKk9h5A7NVHPZ4B0ZJNxVn
z1b8EcOeGaCNAsrybPZx5RfXcsWBUUC8IVWxTPPcpZh5m5XFrjvBouiu/uL2cK4G
S4zBDW3WPlurDSdX2BZhqVxHInULxO5QhwPYAOUuU2e8BcnRbV/AGlyM8IgWlSri
7avbuviC+6lRSZdxR/tC92yp+0QCoYejCLJy7KqRoH/b1FaG1QrXlmCOtalVohAB
CIFWuTESNg3gNo8zuyhNO67rmDTipB6Ht+OUTNaE7lXT0e3JYlcQ2X8dKo1AkEBg
jNCi/K6QYSY383e9FnvwG5rJ6biY7ezGP+nyQJsmzstBeadEjPVV6lRIj/bR7b9b
hte5jcTTMD/7wkrC8wTdkO67dJN4m6wJKQ0oZXKdILlzPgQ8IIeXUP8dOXmQVfR7
wF47Kj3Pc5JP5X5QIUNnBNhObow2jj06U5QMyOitrf+q7A1aomDJ6KklLqwhy6bt
I8JdQxo/lVOwwdFduaV/+9dta3BCW6cW5lB2N4iERoeG0sIs1504xcx9TOTra5OS
WjQib7JapcC4pnJA/D3exndSSO0i/b9pP3nN7qqXiu2U9c7WWNoqAgyfVG76ubIX
aur+gWB1dER01oAh0y6Wg8HntFJN9IDg09PUdBl7SamNV+NJDWr/9C7Bhxyz22YB
COZoGJJCOTsCD8MeILvrqY7uA60LJbQqmf/2y3AAA2G4jXNP1PaoJISIp1HuQVDi
fzB7RDPU7YHeAAhjCBGUXgj9lhBsUxiYOJ4V4mItqOEOR4mVs0J2pHGjPn+DkKOJ
92YkvphAzc3AzxylTmCMSV7Ti+0KKk6a94qbTVHm30hywGSQFjCB0D5q197eYm6x
7s5hl2Di5+/TxA+ggxWkca/4JWsh13xi2PJMtfb8ThnXW/4TBCgzcOzEyZHHQmSJ
SsCgiyPX6u7rpaaB8Kpm2Oki+l6DK+EJjWTMVkeNb7omjy0qVY7ZEDIW0lDHyp8p
pkKOcnPbcR68vFXle9+yR1d7P1EpeCMC/YY5OTxJWII9zwukQAxKPGI3k1HNAEae
usT4uVq6NeuBIhhkTnLcBqjvCfuITQQ7reXejKNLjM3aKJ7NWRpXOVIpoHjlTEfb
KepO1Qv6MaSWXlVCLa1H3HtCYv0tHXIvZh29+uxox+8c+YPmiDcci2KPXR8sf+JA
TzShOFV/a4xItO4IRDt7eOcg6x1Fdl4G71Ira4KRp1bEs/KwXXr5zDAlUXu4TGji
aQWgQcuVRk8K3kLk6MYqWVbwauJyzinYb0jW+Z5nXlWkA/mWfZh9wmW+nGA6Z7gs
KbP6rox5QKXGTd/GdacZdsirzN2Wx/WBip9DDnpIIhAw/uw0OiB8lO2InnnS5fYr
NePvVDiB+XPfdV8zB7zEjmS+sTbMpf4O7AM6DqGgeQhX/f9F8qOMKCGxnU8CjqOY
ewzwleTE3jLRLfuRlOWTdr+hR7EMHDvAEMPH+/uNEcWq4nM8OE5kDjelo8AwUhz0
lvMdHVOcUC2kDpopcjytbQMxJepGMi4HD0tfPLdDsnFLqfS9qKBmUMgtzxpu0hNz
0Ka52kNGWz3C6LWZpAVPfG45r6TMfzRaw1L/8Gl0tVIwoWZOI4+rnWHFnymcNXO/
gzRgWSVu93erslOysmlYnxZy9DSa7Sc1YOp/vUSml7VF8UzS6UonVTKvi6Sk3RBz
1gh/NDg29hQ+yCbG/2QFXrFQp2xqGpsukI+y1I5QUTHN9C+2Z8XiRlPq1uOD/QVB
YnYRYBaSwjKv1TkqTHyn1UNaADHDYqIpgiVLPRcqim/scqNSNr9CD/eqqG12g1di
L5Gr66A6s0NDPSbH/1DeDErewU8nLolpjUvQ0TGc+XLD43LCH8FssUJ7dxMWZcLf
wNAGqpZA3Ruf7E0qjaYriwRuU+KYtlJUUIJCeNsJJOGQ9ZYKZ23wmKd0WykVDPLV
hp+k0Ehib4965RawG+b+DrlRrjJ6QIprT3pvXAD63Gh5Ln85ZXTS1eOlN8MCpqWn
BtGg9UOJgqhGZR1dFl9KOw+UqEqvFI/RcEA1i8uerhzqb62h4in1mwNbmTQNWsKw
CK4qtpdsY7jSdflfwCZG5UXsFolHQEmLNEwJA8V6iaJ5IRLyfzWZItSyBDyhtAbH
y47565v96b75g9QjYL6BY9v2F9I/o3xe1VgfKrrypsDxUZUpL15JezIV1SX4brxo
DpFcCNs3iTYtFZjGu+XSJ7di7pSMMLo6jCr+iOYhE1lKwTvdPrG+Qkbxj1tclF6s
l4zWTM9FcGka7dqTFsp6WlfVw9W9I04Q9IV6oCEGIXRLBUk2hTeA+XBFSmSqCiLc
r24m/TQpIwDf0ohGn56dtetSY0sNCEdL/pa5fOglGrbiFkWy4S24wHaAgS6oUk5e
lfz10074kO8w8AIAfoUtLYuTAE6CfaQU1cD8usZtIu7zqWQgTssl5dSqmMjdMyi7
j6SjOAlEwAYeKjzStoEYwFU+Qe/VSdegPzRemcAvDnpO/aBwL62eE9D2SFVFI9Vp
trw4aGcu1Vdh/V33tS0PojXsnsdVi2e1X7U5r4al9NG5z6e5fRhiBI6jSEPvQ/LY
WfbRwK5C3mNodp/Do5m5qEbTqanZnuHG5Tfa9Vs76KfLmVNuWb2M0pxOMWWo6lPl
RjRzXuUF5D9S7AgP5UJtd4FYnMeXnFKVKIH3z9fm9c01Ah3aGEm/gYjSt6gQGjdU
ufV+eU8cCCUTiwLwIIu2zFj41riBeeo7PmVTtO7PPkTBVejU4y/DSNrjDSk5/r3E
C8gynWh0tFWOWwUaEzI2KW/QpFUJ38LSRfEsANXvZmi/B1MTnMYU66HW2QSCfAeX
uQRcAq+5niMep4BZkzNhW78bHL4ID6LXijLVW/xPXy2rFkUyQE+Gr/HrOeWRIbl2
oqsiC6dT7b62flxG6NgrhDZx4Mko9EvA/KQ9O9HDgwJkptDFKBjjD5ovAhMXWHJA
7taiErv2D2PVsiQcqBcR1BH8W9PldiYuJ/wAIh95Um/mOUKU3sUP3AtV38dnOebq
NKrOkGZ+CdSViAmaueArjSk2SB+XsDg0RE76lFs5VzgAjBRUyxzXP1BnejEIl8w1
QJXqgo7/7hErXTEEpdtC/SsyWg76VgK14ShZDFZ/gh5clKEPEYS2DLrRNjBXvb6c
tSySS39s0yk1LLPTr9mxuVt0fo5RI/sZdJaeys+P0PCnw7xfyw0285CZJPbvlffW
4pGjQ2zzcYBrp6rwjyfztAWzhn12PnMVO1w3enGMFk+6HJZCGsFFVPcvt6MJRdGt
T4513MLTeBQbpGCBUORo4xRBU2xNii6THhDNxPlz5yuCtLKWjwt59dlhMJBPG3KC
Uc2NoE28nwD90Z/1TwBB7VXB9UyPzTfecHI40XnCaSjBF+e1tQVpwLFdr5NcE7cG
7Z1uoCYJBgRmtxqylPDTWhW2z8I4uUL7pPDwDQd2KJ0qAfOQl74KuWxFwGgsng7v
Ro2s4r8Ji3Cjdwbl/PJk0GkYYacVHbNwp1Ry541YNC/pUIaER2LIDB24wSba0Orr
rNsSOABb4HsE7nUrR45m339ffG9e7/WpbfxIMvmRCvZh+GykKikYRlxEy/2xEQqM
vQ7CgA9br/tjU03bEX6pKUINTDSQRiKpWSkhYL8UzIgoThueQkEuxMfg0CFS8Ar8
12miIrToSdgDrUEmODZ/QYZNC09Vvx09c39RqFGmd6bEnX7yVY2+dOEyKgd8CYn4
LdAezD2sCHKwIGswjJVxwZCIlm4wFs1vR6AG2Cld6ltVxHw6UWdObMP5FI2+KPVM
l2blOl2SWmeZLmpB+9bto4enf7decKaiKJQ8LimGdonVrpyo5+SfFkvimklyIl1P
uf8iCgnQboXJkt7gU4+XPEG4U9dXfivCRLMh9XwwDnYcZCwlfvd0679rMxOOXvjl
KayHx+UjHs6/IKY5/4nog/dosoCSf1Y2hQzBj5ruuP8YQHo/v3YIpIy09NUOngPu
x+BDW6Wbv5/Gdd41sElLVe5FyPXOP7AlI5JbvxaG7qm4VdsDxjzbFv8ta97BqhXf
3aHz9Zd8TPw9bFT54b2hu/FalAlNavmV2qpFrNWbMlbBzLGy3mYcitdaKveEyUZb
60bMJME3cKxML3Y3Z6BJkn5hYgLeu5AWznkZPIM1tl8mSWrdOZ4DFxq+Y0R8xoAL
txN+3MVAOCgTvCiNMjKIEg2HUV4NsnwyaHiPT9v2dk4lSTsOu94/YTvAMMz7Y2Vq
wlyLpsyqVefvIuES5fOMIGpVq5Dz/EymVq7Srjczen8QnMW1+kQiShRuBTtOgY/3
Px4ab0LsTEL0tepg4pgKXOwflRqP739IuA7vy0f9UuDWlWmNfl7QBv7dmltaPKa7
P2i1R4WkVq39tyGU+EsjvozD2GUUZe4sF1g34NO64JZ9BAfkOG3CUYhbxLD7yXr5
n5Ak014V0xGJ721Y+pIu5zcDroHK0qUiVOQPn3s0WVviZkIoTbM0P9/n0npslpnG
xeBl0jsJHLIdmu3XZVCWKu73KtgJ8F0DGDZNxJ/Jbu+Z+aoDXrUB6t14vIAN9IU1
EW+jeqxoOy6FsN/YGKzfdOeeJmHBsYcaQvIS9qDEbEjgv14V3yN+TNM2TxeFnZYu
BSV/xYOZhfyz3onzTlPGvra0riZgvp86oXRDNFrzmNUAcsBTJPeHP+cJInft8qv0
BCmWT5UWe5tnU0OPXKvBCBjV796eCw5C0wHjjIOBOuQvsUPJdpVqTEK4SwOlsWzn
W48cGpsFBDkl1qjcp8vjk250faUHf1T+FF/aUrKDqXkS2qFgZpFN0vLvKZFQC1fw
+ZNOie84XAlFojSK/fh7V/0fSqqMvEusGswOdVcvXiUpaMiuv1AvrLkSJrnMbOEV
q0rEopHI8OOS3RGfFcE4n6/5stSF+Aa/FfFdKMr1XAUZNWFA3tXnT/nqe8H0RX5/
JDFr3sNg4B+DzaqFlzkl1Fx5mDqu20HPV1sQB1L0S9tKQp8C3ldh/WzOK5bv8Psg
TCKlvMV4uiZIS6IUEp5+7q/ZqFoU6Ki+pYUXVZ7MyQPQa1CHpWFurd6KBNkwKnyl
QWJ5LAiiYMzlB4ur7zFJd2JxgDTditRiMuz1uc8QupT+oYINj6w8l6U93TBxVM9s
dYmJRNGsM9tvC71/3lx082Y5u7ZTAj2CW2QAEKBJR3jviOFQ8svsWTcErOaxN63t
Dd8VyRATLcGuVWYdO/x7rPc0vnixG9GYBzl80BAF522qWYTrZMXu89sT6IxmsfqG
Tz9Bbf0FZRoX3Uk+PSJs2PMnzPkQtPEAVp2l2808gLffznNooajVyCgt2m0M/V7G
D2/dHiQHr2FpE45IGGT68q68rWvBNdZLbz5zY1Jp3ckKz/PAshr4KWy1aL3oYLEc
5LKPdTFTfSH3/1JrD6kAe1wc/xEUzmk9jZFwACYUPcdx8QsEdFsLTADqLwX1dTtk
qeXw9GlaWSEBlYrSIKwzwC1dSpAXtfc1ypR0fZTY1HXkLL6JoA78WOV3QDfUmWyP
E7NmTzzU8zIO0yvy/gpGyFsYcbPsa4ryHpmLy8BZWQ8ibNItRfPHL6ag6b4dx79e
lDTGQLdvO3/t3eCH/a/gmeEN1SR6A4LwmozxFnOGyUhm4kryiXxxj1J/I/0FHeUm
qaSYWG4j4OVJ5aPG/Mia4inNI0Qhj1oVIGDPjOYt1HnNReMfL1+Cb6fiX0dNHPGC
1BL4xTJGr2C7eEpjCnishSz18eWCXIU7nkg7PFqzcuAriAJ6sdl0g3TTJjk9GpLs
pAUfP3lFA89Cve/TMkypNuZJsGimMJirP3YeJqIUmvLhxA3AyI4zOzIsoc/tQJr4
GGUYqfVA683E35AfrHu8TOELxo47tmeBP/RhvaAEpZghg9GZCXWnnrXagerRjF5s
AJsZMS+lyjJOZvrpRluXpy3l8eoC+Ato5nHlk2eiPXyfmp5ll4C5WF4bhUy0z/Ce
OIrvSMbwZQP9JO2S0gXeuryhqjeDOBIJsL2iINWm7OniCQHfGi0J1QfKI12FgF8P
O/7LpK5EIW5rciv7iu7qStZF1gx6083wC6U9ZdsCBwh7S9c26/C8/qoiMWQjRPlk
uSxOGY02pZpJbNzDWII9qd7/86Jfoxuk3wlX/kz7XwYRxsNbcdt1GPXSIRFjR9Qx
kAmAubxOCY9LpaikBI5f0ZKboyBlGBti/xhJgCve8JVSrRmCgxwD2lqhN3Vq4e6O
sa9xgOv+a6wYde7ZG6pkq9alUbJ6o9qMkxGt/q5YtWwBUJFVzUjd2Gx9dUX1ODSE
EKCmLQMu5wIBKWvCWjR1tONuM9zHmfuSwQvQtME089YA3Pm9q37Nr24EZXclBBo4
yIWGBIhlDUFhNb9LAgDjVc2G8c/sRZzGLn+GWM4TV57fRJT5tSCZlSocM7lfmuxq
cMiE+jfvpzIW1vWyhjBwtlz6uhxArhdXX0l4xMMqsMiM7IUkY+zyGup3RvfaCic2
KvCfWtA2JLMh4vBWbZM5RhQ/8S481p7KtBtuw6AXm7MzvL4DSOr4qmGuM6NC5qdu
SzFli0j+HQT+ErAoAs0Vlc0Id+wtcyWE+AXw2R7uQddV4B+ip/dWJfYQFQCbjPe8
eY2fwqdijkFLjipXZlyZbTKAj4Fwq61U4Lb6CEyaMXZMq8LjG2yxAjsdMefH95l/
YBisbQOqq+ULDeXxgp4xjSpgQU1YU2dTmmuYfFLZ6eWhNoNsN2tKBRBDqVWmtrSP
LJ1smJEFwr9VVYORlfEG4YmuIo2C9xgB5gO2gxdOcKaGp4PNTkt4C9u4DOSF55OL
Eezu2qUZwenUgij4lTUOoKEJMMCSkhJ8x3S06tHuQsIqx9aW6vZIITNpOoCTGR1j
nlIE7hXPuUwIQZjYgRnCmUmMuzJIh9tRJo6P9DplFX17dpJKqMB8PIkLBlhc1nY0
oNp3Uy37mpKYKF8GUn0n6bEqB6yzDRJLqT2mdw8+43CjAKJKPzDQEux/dU/JCZUK
t82b7yz9my8aFb8MsIRKJcJ7hBi5aebEZHChKxo+xhVjvDMN05tlvSRgNDX1dudi
9DKh/5WBQ/jyysFmMAKNsEImKQ+h5/5WeICnRzuNzpopbKTvqgF2rhpGdsGY0nuU
wtgCRTKPhRWVZQ8o8nNK/hBDKiyJSlzaWsZymG/aVsP24kOTK2k4LZ5cea096Avd
HKK4bDlhBZrB4uFXgovUjUUV5jIb6KA6KNdDAy4GHDhIgkTgKvjPv3zEWU3j5gI6
NPjgkyr3t2rtYwS2/3K27bV6ReQtkXNL5KQhG4CRXcqOSSo3g8zsV05Zr2pRklM1
lVN0jOwgjOAWjOiFN7MYkKehuosCEd66AMmszAguY/2TMRzjadq0VGhr9j4QAtYQ
onbZICvN6BALt2lU1C6n/vQHCEE9f0XN+iAiT0Gwd3VRNvzR1pj0z5/HPIOwb0j0
VAPZvkTQFiwFyoqsEoD2YLyyYs7+RngeTeSwYUDeEOMSjO0QDuxDaydvxFkLNhmx
UeA9FMsfE85BxsmYO6Q52IHR6EoHNawSCrALPpKduvOh4w7yfGTxtp7z8dElX6EQ
uHIm0HfZP811P3acozH4dWy6HJuamvz2BsVqLCqgw8625eTw+8/n3OAwIYP/a+JP
DGZZYwJWQfBI6z6M8T6RaBrbW33jumjA0S703yKYBKH7s65dfpwqMk3OuUm84wNm
hVntnf5XZaV2uqGm7LQkMhmHhOF6FQ1Hp3L5blitgM4HK+fyV1HgWlCRyN4I7RnU
MrBNZ6PvFSc1T5D4QixTlUOA3wIYsXn0qe7CSjNUxfDQgYeWvOtoKQAD+/qWdPoz
7W/7dleo/SGmBX8YW4ACO1I43PUv+DYg9ZDu1hAfwRTSLhAbs8QKyoPqctO15StS
TB3/AasJReA+xDHW5ZqLbiTKy2Pt01NRT8OZPPvD4DDEj/eFMpO4Q01sx6glavm3
tz3z/j1OH3cbLS/WmHlYXdz8D4VcPyMJuZOuDTT6plG4VZwkt5I0OBZR8VPTbz8K
cYnoNno90ocoo1UcG/X5gHFhIBtBoQFdAgH2LLc3jlkjgavsvtxcH49z6CZVaYT0
HD3JoTOyFKir0GLfozeoIuZseVM6/TFb0JZ/oGmK5/b7Ji//NkIYI1CFtwWd6YFh
PjUZrueVRKFZm0bJ1V11CmCdVEr7Ofs7BIQ0Q0MfHe+MyLiNKZplzjLPRW9zNOe3
9j+xLc+d9lmNA6t7CECI3yKOOcg02pIksJH7Q4hyZaRhdtk99EvSmBDte6KbCRS7
rvJVzFYKL7XhNA//c0pRW6RKgidRVIKOE4QlNiupHiZkfzbaRnMQYhMbhlBpDCi6
lhzViTZvqWPcQJppggX/ryKrgbasgQnRGA/6ER7LuUlOETYjLS1D6rlEO1DZOTx2
svVe7cwxJXB+1ecwrmRmWcGw4efCpTHZTPgJVzV2VvZ9oARijTTIrpTOqN6JaaMj
aC1hX+H0EO44wKus9j17tvI8qJBUmbEJk/J/Z/bvmIuvzNw//eCygfDLboHTyP78
A7mT7uPCf+PABKbbM6L8LFSVF9Y0JWEvAvxCbInRsqH2shxqRQigABGfmudHfRhB
4Jzg1F+goHKJixkQeoLSsY+9i/0X5m+pHaxYk5wGLGwUtHj+C0r6ixWtOH6n3b0O
Z20e0TOgPMSXBq1eWQ7+SMGA8vNQ0lNEyJccpw1cL1Q3twIQ78jJuSEw585WwN7K
0agB2+j5Kmy9FNvdonFnBdedYU/MYohmwGI+oP+oCZN8IgWCdT6Mn0qZrZp+4HSp
Y6igpz0Ag9VW8H10Rqwl6ZOGqEf9KEj60ZWNOWOukDUgp6vr2al1SGabAoZMxzI3
aLBmM9s6ww6RgUzJv2mJF7QwmvxN51R2Ojl+I5Ysnxd82s7ewL7DZqafUzFBB1W+
QmTLgWfuuOUU0avaRRSFM06zU28tWY91S+FPBXKHYYr7OEV81cjx+k2RUCsv71nx
LNYko0rDR+K8skcsdSPd5T+xQzsriUjCOmC/eweMHuC4zYaLzR01I47YM9/WzEMX
xIeWooZk7vCpXtAmCoKFxJKwYp3CL3wc3MLBQCE45nt9kq1fvK7xwIfMe9Zkived
JmywPOLeIbT1Ci5niE15r8/gQwk00VGRk8mdy+Pd3nwgxjeEt0DupdrR1/nRY2E8
eWIqFtklpJuvxOIx01Bop0NLz1oCO1AYGs/U9Fh7/k1cV+uK0zxlsCipyoC9hPDp
N39rPF/m3ZLCGKvqco0vh4Ihrzb0CczqogHwp2iXF6ZHb01cLFWiF0gVm4jIBft6
OD6pLHhuXH8VNo/nY0zhDthKTPG96QktofOrQQe/X3tpwvCmKqDjXr0FPYeIVVFf
RhBmiYSECW/Cc9hJXVtFVEOm2PqtGEZVjrM7gbLnFez9ngOeaMxLNDIC3pPcOIK5
CXshT45bsNnLO5ucp9FKKZU10Vz9kG0jL14t8N7Ny0iACyDxBrZ/cK2Ks2eqxn8f
10/DWsUDrd4y9aZ6ux+Ossfv2Qq0JLZ60p0ovqzDbzz6AqOhWnfUmsWKr9qphhuS
iPgpc2yEhEe0l8vPPMZfEF6fDc5nnkPa+Ro2yKGpeyl99fnTBumbeihnadg5IaGc
EWKRCpUF//ucJVqWKdyk/Gt7w9aX1Qctx3E3Xc9ZS5n/UgF2RYpoADhw7+Ycc98A
NaSeU5QSHyo1lGX9i6rl/bvPVfL+WENH+73DKDvOsHnEVJdemY/s9jY9axOieuiK
MUIY1IgcPsOKmsEfAkLrK6q2ADFDMZrMKkphfC7YkbEnO5k0dkqxjWF3cMD7FoNH
TDcozNucRdpiAgbZ0FoxrMU4HaaQKTbz+KIN5fEuF0L088g2DMta5ANAt07dqDsk
zYhjgWS3/Yh4J9OeZcvWMMUyoHZ5TCx6GmnqB0VZA8BEuft5+UG76mT5SIj/kegX
z2indQ16UKiVGLnnwC/fqbKENTRNgEye3Dkw8mh4i9QGTLxUTT7dloKYTjbWwBYN
0T6FZ+FYRBMGkPxwlE/RZdStAvOeegMwK9sGMYgnXmVf7xExfAxGgzgDzWfv/23y
bIW1qqUPyXVgfrhXgWC6VlTzfU3J6RzGfnxydzs+fmqYKp7uVCxT4NVnFKEPC23d
cbl/DZGZXduTcXdkZ3Bz83WB6d6IDe5xaZ9oLuUdM+iwkIlpZslOTbVeMRN3GFN3
t2WE/tbJ3QRSnfX5uThdXDJ5l1AkCLt2WjWh6OwdQPA/Hu/+2luoIG1wLOritxRC
m11eel9CbjBaTRle60RBeNftxIO3AWHwnQMYagQ0Xra1zmRcdRoo1Gz536jgp0t0
8uf9nnyoBfGqfDkANlbztONUDtv7kKS+htihm4dniCeEoOWbQVcw1Vuetim3Fqhy
vW3VoFgdbP/XjRr958Y84xzAIRafkAsL0a2pp6IoXaEmUi0qcqiNQTmied63g32C
QsDj6sREKUjhOOP4YT12nIKzmOYi3UZzzvRtWo5fG7SnnM4NIm6cC/d6Nctm3b3f
fzZPXsSOIxP/mu/+icxtG+qNKVaKsr7J7Ee/vzOxWeCgddvIPBPe2tPq6i7qNPPM
UDxPMSoBrXSW/j8wm1LesD4yRbYEKgpWWwTfW2mmvIsMHIUGTBs6HjING+foN7dN
LPA4WQ9cum9Xt2O9nS/JjM8rx6C5+C0jDdlf0EzFnRRLBQxf0JRApL5ipAyvp+En
VIHNLdUHY1N8k/mwVa75Dc89iUA87e7ZYT6ZGmtSyVtL2AoM3KdPu7Cua3ydpmYS
ESESilK09Pt5D9Ud6iokSqTLFokm21dof7/3tNakZx87pBxLeRXUwGoG6C+eogti
xGN1DIt3Jt2fMw6DFdpEcwhg4aAExdXsHIyrVw6tXaGJasv9kP4xV9GQA8JiAVP3
qasywCPp7hztF4tuXYMAToiQ8vJMsxJ8cBg84X8kfEywcvvTNlUniq6GfaYTvG7R
N5a1fydbHlHn0sjsplxUP9MGQzFHunsl5PKl9aVYUFhK4pyKXFaiR5ynfGiA6aSR
CEZSuuY53Xi/hz0cTFMJMEjmSVcLpgsWnqa08JjztDIv6Q/stcmjE+rPp9OkQ6yN
7TeJxivlkRPl7sbw9pF8HGs2VcnMVPhBxNglCZdXIKIxYFwRMHRA5CUgtC4M5pTw
dZj4tQgVjViLeygA8vhZUDcTcbbgGMOuC3GhmvizQUVvd1XM+SbmMbrEgd3P9jcX
JtSOYsVQyZgCftCKTYBTsSezYr1uJKvtRHZ+Xt3jpC0Qc+FGWKGedPTcOApYU/QZ
2WUNX0PowiCv0PG97InTk8xGAbIVEelTHC0OJPmb81Elp8nK6+/9uE/6zxQcTnc8
BTR4yjJhsxS0N7ZhQWr2dwCdk4Gk3wrtXqWCE7jKD9rdwwX3cg69US8NLqcbIO/j
juijICVB8A/sCKAkB2akL+0LYlDpjyYmbfz2u/YMeNk26fk4gxMtyaiTvp2Tarn5
pyxl4HyXg0d+6tmTrvQRbFRjbUpZKIfU2LwjgZ+C6hEz3rVrNG6xU4+/jLD//z6U
GH2viXYxe2Ab9Mcx4y+jAgIyimb43u+S8VUmbiZCPGap/XSBIqGtdNUYQd+EJ9Wf
XlHCHTlEYf3fK65fdr8LVDtTVEGDLv0KDxc987zbWj3Rl9QnRtntaeG4ZATbEFTo
EVj9qwmyup3cxAjczTlazGgKn5MqdTenSMD78ENQfuXPacF8y9TDjAPddBiLX05g
3GVFp37c5BSsRW4lFU3SoUbiBKLNe7GRtmvrDSNhwMUrO+MHnnUsSu9gRTScUNSy
YpLr4tRafTLIDl+vhMH18sa7C3hWKgQ3vj6MzreJUapsU7TNNAIh8XDQygZRl5lV
9BOPydejNzR1XpjaeL9n/23qBiwGNnKgiPWb5JT6rca9r6jMS0uoeolZ/aOqhZ8m
GD0HZxQbBNBmbfqve+l16GdyrtRWd4OYRTX3EeUEiFf4uYcHG+m/9D0j4mDQa0eG
AuPRlEJWvViLMx839UEMrR7AQf3rEVmoJnadfiT2ZHSyzNGLbI/QK+FAugWy4PdK
bJDvnnWWaw4ZSlHWWp0kiMyjZ8ZWkz5O/SIVAGq93gN7Owjm4IX+B8BUBIcMXQp6
kPYOGZvHpcMImFtgrjL5aJGZBF+694PDwJUdSKndrVnJ9A9BXf7vzb/qNXAYJGar
aJQZtb869+afzHZDB3x8xhEa+6fgt/QirK9A7MaxtUfE0P+sAJ20dNdxeHU5RBBP
y1HNmJ0aFSQnNZILjTuGcyj2yzwb6gPQqSqEAiYPn7x9Gl1wDTl5IP9eRtBy6Rn9
cL5BtB7sdYSttyPIG9x/qLMOGkcyHSfBhEfSQtlZF9OBRWHmawNlpYh4Zd4jsn9I
yVbXl9DQ7u29GyTzQRHqU8vanuhYfAe6JUnur1zVjKuflPgBxvhs8WTwziILwOUI
CUcammuwRJ7d0Za/lkb6Q0ZdjlBF8BvJztaKC/1Ap613kablPldKBpftQxwkXZ80
uU95TXrfnbxhhasTUZ4STm3FtgUaFNDD1J9ZLcwMdhrJCGdDRoGDCc95zEe/U3QT
BIXbolYVfnp6GJx2Uqn3LiR04AXaFfJZJX1MR0ciMBtyld5lbgK8OfnVHf3AZSzb
pDjX+tORYggI82P+d2H0X4mfB9oUDWsl2/H3wk51CcQonpYvzN/GsSyHebVzcojA
JQ5kTICP8bYeBMBPCJQSml9P1CfOWfCyhyn0C3CIoMpso8in78adZhJiSJ1crMz6
1KC0Cs/ty65g5yNec3gOZl1m8paXL175fh8HoHuE8TjvK5xEbAvHeHlqVDIyHj1l
Aoj4LpkrsKHcqADhS8e6cTBF7EfiumSJHtdDmRDP+ps8LCRdNx3s3uUmr22AhByp
jTezxJV6zRLWuhcXItQrCPQVyn8mGbaRGDQMOE2SE5GTXA74y9CVcaMUEEKUqymd
Wxp6uA4rjqIZuqLqUYvYxRBm69IDEGdTQjrFRyPYW4TZLQ368MHIFO0r+eRbBTwv
XjJ2cmQaTeOEUblRiP/mKCBPdZ/VQytkjLKbYjprGFGUQYVhSKHgF+VI9JpDwJoa
+EH7n+b/b0YBfRkf5sb63N9DKEB82yBAWehNJjZuG2P+Qm3NrAVqDLSpjdhXvtj0
mk3+NekL7Yb9BtGjOK9ueT+J0UsENBuO/OelkdQcsHH5xOKNdh8dYShUzFU3Pb/2
vdmnf/bdzrxAepIY+d6EYgzWsXc+NyBAoi7dDV12KOhcSBeejFomGYM40TAiZXAG
WQ216fubrJPt62SJHG7B3YFm1/R4Ufnsy78aucQ8nB/S+0yFHM+4QWfHwvcIy6IF
bGwVYcD51XVmDB0aLVa1MvmfwdJrEiOM+JHBx9iv68/AaO2GNF2Ly0dTQ2mdh4E2
qMw7tqyLuXdXqHPHaZQ97n2+n6Z8OtvAHiU/3gGAK71aflWe1h3m6lO6wqQKnc1R
Dphk2xxmBY+ESJD7nWgBwL6fSTGMAhhEMuy7SP4HV2RuhXIUn5+tgtZJ+i8y3g9e
ZbkwN+yv0LewVlAjXJ24RJg0xq5SDMD/mwAsPmcvdrIFelLVw2sa4K8WOkR8EvKE
52mwGbW3NBaNFAAYW3XL5bGgKm/HUtaodFOV9KJWjrihcjRVRzXaC5ZXU2AjsOzZ
msVZiAFHLSl1H2EULFo4dXbJxiUJGv4TVVcqni2axPrEHGX0F0mXwf+1xfB0KVDF
RSbyifLZX0euYSXrOdXaxSi0181vUWooDgpfMtvYotI3MpTlkpBJaJy+fNmoPr13
tZN6VD3OGAZ/ysbHOSCN+kPPDKWvuVyAyOy/nkcqkMim8Tkl+GIBkyis18mtWrND
PuoaB4unt3Zt6L9w4vAEd4ooeU315fiaEFxX8aULBLrdBzxoNyiga0UMnJhsQhDu
6Zh8X/qzK8dsafftOJyDTjTyC7kFcQipUAJTdw2SMaJaZEdbF3gukdmOZq9+El+9
vPfC57u81A8+c9nZFgbq9OEu+jLMbajmD3rAEWtMsMD99NHuXr0UUNBlRrUb++VI
Knci5PFY11a41DZv2+mlTqGhFJT5ElzWwIi3hWWlkalQ8GOkB7kS7a40kgrBhM0F
BTlD80DGmHkU8GGRrsNVvwCRw5eGbG0UXoAKNavjqRrUBD5H4Ri+m0qwKXmlPGRv
FdXuIyJeYyP5TL1HgEjywqHoLLtkJelwqORwPTc+X/rO3bMMVFGfHHqfG4hR47np
/iAVhwIM79PQ8aX2k8AbUZ9hU8S1wxag9FucgfKcRPOyrvvnybth7pe2V64STBRH
wvpGnIS8B3vPSq7xYaje2xs66x2nhdj5uNddX/GXypmA2bhBsUdT2fgU7EPeQm9H
n/D0Qz/Wc1fNMu7rsyTvsLDWX12F35EiQeG5HiYFvjwU5EUc4XUnstozRXOJ1Eqw
WFEuVGkdyZlbXB8SzlvRxDf+EeNlkxiWmZFaLbJf9p6S7QSPfhnJ8X/Yawj2MsPp
ZWd/UJ6voNEDEaQLjdiu5C88iyNKX1y0DMfObuuXWBfhJjuFvqRRQ3NBkpFKgFGR
npgaHpvTqd6nRqXaUr0ypYcpRCIFSSiAZlpSDioXRk0WfvYUQwJrN3VZqurcVHLA
XU6/7xuQ8B5gVSvmIXhV5ZOb5wbTTTVlxZH/EaDOaC/9iE6Vu+tCiICBsnEsplxH
20aS/yiap2++3A0oH/hYSNH4qV/Db33jarcD8/wVZyZaOEcBsm9bBfMbFrC4g/xF
hHcxJZLwezzrj1+oxJoWA7erQG93SElQ7aMueikwSXRHL7p3IEy6CT39NiNs1OeU
8pmTNzwUSZ5GKdG1Kkq7vrKZ/V/QeTtn6hpywN4wDgZ9n11zTEngKsHx9fPEi6gK
PJsTf7UgYItstVivo1uLKCLaWwJHNz63+dYR0ydo3bUk0pCzOCQd9aHw7UmKv5mk
+aE5JNq5cdYF4L1gfTQDZzQkpfn36W70LpEchUhWqU9S0SF8HkN7wxuTs++DbMSy
jPIDHPbyX1HVHK1QUZSQh860h+Cw10vLdRZIrygr2vCoKwDzZWttnrO6sBUGSf7U
tzGskT6FjGwHbttiW1Jyb3awG/rlFDs+NR3D4Z5Pq/Us31QDoCzzXihjV8T3PQnO
3AnnHi746/AFLy1UkZ75ttBrOWpbDNXFNzHyTZWBxES+DvcGJEyZ4TRyrSqCsOOY
qdabTAkEGwdBDBgZaTJ6f/0PEkqXrDlnvkVbY7Ujmi5UGImgayDl43JGPNls2sY9
z5zzijllH4n53tGNYXu2sxdvlKD5h53rrqKF32bIZFP6T/XzfDkoOEmUIljulu5f
fc0jYQTDsEnlnbVHTcGivYOo6K1PuYdK5YBcjrUYOho7g/XnNekIQuy+38sR9zb3
aBX+K1PnUGkfpx5ge0OgB0B04P5PPPHnwooaFVhztzqu8UC5Y0Qy3BDl8+fOCcbg
JGrGK8uFT2e49ZxG9vdlCZ/1a6dMyMUA8q4i5A5dvYvtodVuIQokEglml8UrkhY5
lNitZaKqcbxn6th06S947G+DMJo6/l4ZRp2s+apTl25p2d2p/+67hJXdO8Hdx483
xs3yPWftmdgDIwDcNDnm0GLi4LABJFk7HoEqAHQJu6Df7lZ+q02nM1GW1msGHV83
ML7UQOGUS1OOG13e4tuIQemo+Olc5PpmSKVxF3ebwV1w24xuzdLoB2jsSzJ8Nq18
GLwr/Nvwnh2Y2/D8Xy+9CNwCbbLChu2U++PZVQILzRktxklnCTehtl3HIIbrEDMh
3zF/BECBam3KjpB1QZuW0gDth+aRXvp2BhQ/ONmdI1cYKBMZZPWdWQ3hVW6l8v4k
ide4SVUYUPOj9/AkiQfbaake6SaCc3byKiip8bwjPXOirrld+1hDqJo65nNZhcxb
yiUPDOnAtitGdm4iliWL8pJXkqzDNFT2cDK51YO8MapaFPSvs06+UrPlGE5N017m
ruUhYi9Ifwn0jWnUqe40/BNUzzie1A7mla76lR1VvVxIOnclyu8uCXjQyp7Z2ufX
Ubkdqg9XPYEI3zDe9ymcf4EY+x5Sz2Ij7c+UlpfTb8RNvO1fWxnGmKEeSmv1c91k
XdoEGpL+RBPjmZdQXLogjWnjMKGht8nkg1D8DtpKXBlhlhBwnvd6EgwqS0pHZL3x
vvcjqCiritmB5zpOkTKUUYFCav2gMIgrogkTpavaGSSorXK6Rpl5uAJLQ3BjzKko
WLQPY4d37DAjgmpNFOc/Npq6PU+j1YlO5V2prpKYDd3BLkHTTP4SrjX15FBhwZNZ
BBaBSn3APYa8h4lsb517gBI1yk1rvQkCpbO6+oLtpPZ4vyG4kD7dI7EVO/11jOp9
aWqXy3Q54Uusb+lBzhL6H/wASZ9S7ZEGwp1TMdIDFk1CSF525ZMlD7BkmQ6mcPP2
Oa/teJak4XgrXmjg4AnB/+LVMxzidjQHu+xdTn9lI9/qMLRvoPLyIzrwZXF+fkVK
OdpIrvudvA7PClG9WVZBIBFhswaZFoQkig9vjg3oCb6e0qDskcrKa6fyk64IEEwR
I92Zrs9nFZRRG/fRm5QQgm3TF8VMlomPlnVhgNLiD5ONrUaE3V+/C4uk4siDfpom
yBNkq5fQK+ZbZw3mAU+gsfXHIh0BfqcUJ0E1U0F2BEhVNkZA9N/M1PcdUFvl2cHC
e9AmMAZaX1KogOvDPTE0anfwJ/E0uglv1BJJO4qZEJiqilfFgMPaJ3mIyF9QylAd
pI4vGhjT2SyPnel0vJPlI2RhGF1EpQOzlR6b7itzw3ZwT4i3Jo3W6Ye4Ex2ZJhJc
Ttgbe0xZKeVPyjSxbrhvDgfJFXVnTLsAWrNvj+R4uvHBC3YrHFHL0I6WOvcvwtaY
eM3lklnfkL6hs8mMjrmHGcEZZ6rLhuLCCOWYEn5kAA05zbkq3fOIEzilaqjS2oTN
Vt93YsLsq5bumADa42BoDshu9b3EL6HZTFL4EUsk1NWlJpoycwIM+9CeV0TZ+gu1
hRQxx3U+qVpbAfIi8kWiudzn7vomzwlhoUfh8SlbjThVVgklQEZ58QLjuVnOkohv
l6S5n0XP/2mRU3pG/vQbRKU07P7YdjySnO01mb8/XCj5GnX6VxKUS9yZnbno//4C
V6MmbbrjlZEHUYk5sSDsoiBrGalECKUF0A7QOPyElM8x+TARXPdUyYd9wWibTlt5
FeBPAn7dCIyp32Jxu+VmXZDj35lYwv52oJPFCsFVeFMwp8+pcCLMTWrbwl/yDVhP
1YhQR02LlQEfCVq1dzzdzAOouyIGQYL5+hWpRt5S987Yqpx1WpnxzECnG0PYqxfD
lW/qlwsWcoQlDKuuJhRnvUsLRBMY9flzsQi72HxCss45pFp1fPFbbFjkI3cO8vNE
6MDqu60UzyDkEa8Wvr47i01Ka/B0I0HM5Oq5H3nUaEufKOfBELtGesdYtUDB7p5d
c7Be726cGsuQtZWTdC/xVJZ7RyCuXGHwtA9ZzH0wtm7PJwbuYmzRH+0nvpzyiQPq
KWStMxa3jl1VOrRvWF0nm/FxqMmriGg30T4hIjf8wgR1/RWetxQMqj4V/e3ntd4o
Qs2S45HcljYGD0++GN2OXHArk/5ZPy0RUoLLtW/82I7618925zPCHMcTmj2brT1g
F/2VBAgbT8TBoYQKw//63Xq8FuB3enZW2bDcG3xMMnN3xish9Bjbt4qvZuY4JK0j
zxwEdUBvuRS9Kp2qsaRYeOEEBzS39gFUI6gABcJkSvPi+O8NDbw00XBRI4hFhEs2
Y/vccaaiQd2wbbqA7uQVHBdLE1o5qq1m5+8fGg7nzSyAwGcvpitx8IJnscl5Gpp9
5XSDlhH6halUFl2Ee1BtfHsKU6TOwTEj1SqQzrJdjM6l2I0VSFkI8Tezz3XILB+Z
nRkwfvlt7rD5yoRFjlF8zf4/GsrwTkygmo+OeOqA2dArJDCFA0oigyWiOSbLgZGZ
SF1aIBM0zMo9/5wNQjm+aX2SIX5V/mTGClC4jveOL1BWmNSJpriWCzbK12XjH3Ub
kWtTkq7fvJYXkL1hYF1KrIqZgUn2+deCtCzDTdrH3wXpbU+WIxsNFYZW2P8XAX8G
KjVTT7HCLdssXkgUweWAg53i+9JdAX5/E6OwMIG4Ba5YI+ofX96yPk8fRrtG+mQy
xGrw14pkEd86FLNYyd/bKjezOSK7BVL4iyeVf4wSZRdS1Q5FKdxZQ0JmiAFNgPBP
5yGW3WwpKvIDuYui92/Ozj7OA5TMktWauLZZFlmRnII0bijeMnhVybWLmEWAmZ6s
NFwvOgMuw39zA3PDLmsP1BGxrk1f57Ova0bDUlH+oQ17K4yW6IcN/chf2v4aQd4o
0cCvXatbSFzSRoDDm+hdgW8CuSPjVNVq7IoCZXl7nx+a3ey63RC6hPHOD1maHXlO
b983PzKBIRPzGTSCfUXTl0pXDOfJ5yS5swUjng2iXNUsd4e/QYfmcf3FSWb1WDd7
p4pxaZ6fI9cTpxYgSucxsweMUmVlwSliJ7nkebW/+3b0W8UnKGT6VJaR5Xh6fzeY
JOlUSFA77o+7Jzn+6XoxtyaXDX5R4UyIZKM9l3YoIOTfeQ2bqw7u2fYfIAJ2hxJI
Z1OpFTJPQt6zZAQKWdrZAxHgATsrAAtme6xdapNkVHjaD8JGsI8uxPkZZ1tN4vK8
9tNTZCOZw0zS8JXYllTgxHtF9MPWbvAyyZFnwiyB8XeOHcEsqVnk8ZGcjHyJOIoq
7EGz7M883XM/ge1mjSZXvuOLvLeuIanOJyA0Fwg2j0DyAuFMKp2rISqCeiUXCmv8
RslN84+qUqumkDi2ShD6JgZaH6C8SjTJIIq/SqFH+JVzGddGQm1wwybf7r3bLfx2
aUOablP4LSTV7ccTEfxWGXrTQwYcJJ3dAfcrPnxKuZVnCgFViNgmAdi4CF/mQBCt
SzHuNeHadHuGgmmxDsptgMGzKMLhURnPjamWEVvHHbHFW3e1xoHOqLINFr7yqF7G
aQCeUzCTT1IhB/r/wOWyNRVqRCzFNa511IMcU5qWCo7tsorMqGazf9JoC4WaYYhS
41c5ekWXynooyZoKNuSA1vg3WXRMs5yVDoWTyEJXIMmtlB7l2Sd7Fw6ONgvdZPsl
9jMb4lpkODA2MhbVhutTKWNHB7j/57e5VYd42md+DZ2C7xt1xqyHwc7tyLdShD1w
7Amyq4AiAC7440M0ycmOlDQh6OpXwLQUjBS+fcDXxrpG+bYiZw9ammwcA81QKvgC
9y9PznBup7HFrWFrQVISq5TLNAuLzuPRMuVtpny90HiNx+/3QaV9L1cLAA7ecHc9
S4a7KxFLhbKMeALp6InZgjzdTn5XeJUGonX8z74D8cuc2dAE9jaXjV4WcYEDHTJx
06+8KPwR9BNmMvomFk4/tLAFJENZLWhF0yTQUEjS8o2l8i+lU9V2qT3yZnbHYnSb
HkliBHNnBgrNbQVqkczvSU6BRIFGYsRsJ+xCZIUrwhvKjvKfHWYVRHjjLmj0xdZx
biKPZxCkc143+YMVEDiQ67XSXJmbxuMYVdT8WnPZjOySaW41jH9UWh3p0ltCJ5Ws
gtJO66zyF2i8+4F3Hkv9PJ0c4gUSesQfzDRlZP49GB8CSeDV3yKpnqgKEUXXL8cY
1LvyEoxTpQ51msMCknC4dHYRYYx8G+wamD5tTUMNNxI5MKjCpKDe1HfLJm3ub8Uv
Z0PxNInwnHuxNp8bjG6bz2fDuUaWfNETqOpOi7GaOJlsBSrIje4pSMgwgbpfmI69
Im4CU3decy0vbLJ8IIzOWVrDQnYNOlhXXIeiDnUkCjP8he09Iq4P1U+GdGguZbTe
3PRJ42wLri8oOiXs+LNqvaajFrj32tm/3laQ+PYFCHc6UTsVRzdljQsJopoip2aX
G+7qdd4a/INMVOsRnMAW9Gx5Y0wx20We7JBRkJkoM32qXtaS3joQgN+cpyu/UmJ8
e09lHfXtIvXdvTwuaUPU/Mbv4MANQ1miTRPfYcg62KsahTZ1Z/KipJmv3caV+z/a
lDrJ/+1J2bQb38s+59Yfh8SUGAjypgfs1+R3NGLOPK7RwzWZJHY6roma+N/0wAU7
0CJVvahav9IawwUh4538+ohQ3pceQuxJgAFrqNXAPv+zzqu0oQi+d8Bo6GCj7I7J
wqSyv65sfwnCtntm772mvXgJXhlonbhm9NNKh+BOfdsDzPJGy7ARgGcfcMcFVpIv
x9Xofh7Lflq7rQeTbAmlbFlO0P+YTLwwLE3ywfoVLRAqcXU4mfo75V8npZ2ak3AZ
tKQPmj1ADa3E77Zgw7wx5etvoVIrmjwEEnvHdkVjK9KbyISaJPI+GhY3El8QTl27
he7OG4d1VsLR1zTFrXYLuau8TbPJV5z29fR9m9o6qtT1vFOdIqIF9XCBioLwKKCl
iZmEvRNwKQB9ivcBEuFQ5rqJ3hWD2hTiCNTo9XrPuLFQ1Oy3H2EB9LLHwE/Gtw3R
j/3DBW4Ic2dUdZdylxMEl+/6PPwAId1VilCVK7zvf4hTDrvLJRabJzYkpBN8c9qv
UecgXFlDufKu+Ay1O2d0Uc0BQsYDNJFvRJOHiEVOdvMs2NT+qBpWUoAnYw58YGLO
2lmF716BCs2ibr57wWWfDaPSmigX8RhSmIctg86IKwzutY0JBKRZMWBATw4HOLE6
kJVcJedTpWLWA1eB9E0tUCQIVTlMIEWdjXtN7lWXJ6uI4Y/5JM1XV6UfMozrvs5j
e9Fl13Qz0dGB/5Hn+j7SZr5lrwjBnIPjLZtD7QDoJ3CUG51N4I7cz3oVMPHN/dxv
w9ckWBrOGW5Lfxzwz6yzdkBWGs+fzmpEc8NvjnMJG2ID7icxodCSfvKJh4mLDDaR
aggNABWO1y5lAJQvIdNYXUObYXMKGTsEZ85P/imrulB3X6RPFUgSiyS85HcEg9Gv
7s8RIl5EudEpcMu//KLvrPbd5LdLFejI2399gc6QK7TjHc95LsyLlibqzVAl0zaa
sFez1K4e9BEylR/AKGs44Em0jd3XFH3O2XXboSX4OtVh2xXVz9mt8zCfB1RZwz4b
zy8tTgvRoOUYFoqRiAZ03BM1I8RvSNWRFd7cIoeVAgaZDy8OyHKMfcEjErAKKKhh
6FqSlgR2HRAqyD9eVINCB035o8P2v9+szs8g1hkfEt5mRacSyj8fcfsiLpmd+Z7p
YCW7GTp96AnQwC/UDZi1zzCovmjWnTbG6TUqLc60Gw2Yp75HnMdOPHHWUWtiXzeq
zsbQ9ZdZuRUe12QcBS2joqJudMMhL1mhEw/IQdCZPbyvkEZYMY21SUJoz7Wia8S1
rzrfLn2TpnV6FwX7BS0rsVj1TK2dh5OHOguXcSS8VhYWDCb57hqSpBS822QuR9a8
jH10LN5UsDPvLfnC5diJQUlUFu2Mx/6lrCmV2fQw9KLxQtbzRVwCxTWY2mBUC6v3
WuHnjT4PtG7a9iEu4mTD9l5/ITeessXEm60ltTSw8Ekx6CBfL+NbKaz9n/zn1FRT
xf8yC5lbK3KlMOZqmdoFhofACI0FMY1jCH//mHcRgpVQE5KYLzSnEG6bJ3NtDrx2
GsR2vD7fhvETbF7fsemt7ORBo3uGMjkkUCFtkmNNBLlBCZGgxk67zTNmLqsXZuOZ
oGzcDZONDs5nbH8iKR3CyWoeM67BaaxblIOVnDtfVo7xryc9Br9gzzNR/nxybvjn
r6gpzpZbEpdWszjKXdmlDSu9GqwrxpqaPrko2O+0kR8kSk+zdcxJQtZ6YbC4XQps
Cr0Hwr5QC6OXUR415/R2767O6MyehrE4LeQB+LSvnh8rXOKM3pfbq8VzJB0b56dx
kWA4M1pTq6TJqxVEOAVT/S/12zRmSsgfP2+2frCS5+pv+0svcuNZOG1wOCsA9Ywt
Irej9/Jxfng6SXE9NlQ6R4x3/p8jN5d+9phQDLzrGG4la+yjzWqWsRVCdSzjcHjx
jmzLTFMzk5McYsTYSuaXotDNMNt7kRLndDb/RPGzqg8tp5pJFPw/vf/7F0lDPRVD
kHwDqGOQE/ya+OQU+9jybe5Q0DxtN7F2Rco2bHFAM93amirZd5lYM8RhLyLOB6M6
zM7+T9QLPNJYXQr59C1xUA03zoU+EvyfEX2JHPZV7W0+yeQwmUcqDDRjzmVEk9Bv
c9125zyrKPt7lfy/g9b5dMkxH50m+YF2f7HZFxaX9xJfiu0aNJ7ug0WKtR3v8Thn
YCh1+fjYD2+XuBUzaLWd7D7bIFQmv8NBTfEWkhHEQIeLMM+xhG4hs0fsAFWZnr5O
+T/GEmTRaJJAhEg/9DZ7Yj6RGZ80jB/z/GiAd7Rtaqybhr5auYEoadxm0aa3hAMr
j+IKa/5MUCTv+4VCT24DPNCT2WW8rIBRopcXlNTrYPRshVKlrzupyxTTzvCTa2SJ
vBJtra8QLWMPlOlVNjCcEje8kpe6pINNadv4ztmcmT4TJ+U6ArKrG7vdD6ClWRZ+
PEAeF1Gyn96moJ/SeHYnhpZlRqyiOqWJOp8F8DthDQ017HZq3pyYUj16nMIbxovM
vUY/mK9Phh3FknB7rGCb366xG38Puewm2trsfzVStMZ24MtlzyvOxBd7nISGHS+3
rdfyuZ43zy9U9licmnYJP3fshuzLJHpW7Cn2tRFznckBdMYgNlPcsAYibqsPSMND
sqkrNd+CZGxLiZKTPD3hGjDy6vdlidC4prlgmpze5kSgXriZI4Ql+XHzlMmHTfuf
Pry5WBi2Y8C6eyKxmzDCCfZZIVRxKE+zs85uASqeFxNa9acYXyWA3ZFSZAnClWwh
lyG5E4LZ5IXXGdXditH5oPRTDkrLcF5FKzfHufq5ayYnHCWvJj42M7QUBKZmdzJp
xjcc4pjBq7p8F0qvdbn+jNgR4DBX5CL4584QnNGWj+jkWeuQ4/ywQKRzWos6ESn3
i8OAgC6ttx53HUwnkppfCg5S0bhO96u1dik1Ej6JA8/iZA9BY6T1SU6Rur99Ssiv
VVJ+JddDJT5eAcOhar51KTR+102TCPoVUCGtOgwMYaR9rComHbmHWUpWurfsSadn
vK/wvSdOGR+BQnDEJuXf/dNVhqnG+LxFnsoKelEk5JpoR2XCtHxjKfoGTS2wZHzg
AFFVhT86BcSbpqkKt4VJAS+gIdgdQUrLzhtWqb7RvRrY2vHneGdbPq2Lru49MHcG
Och9/gt5Ocz21d4mViQBPMTOAMduUoixJ4AzSEyUsP92zDNWTbdYuvKPwWvVFrbg
qs8eoVV17R6uVpm36VSAI/4SY6WZ1k/RFF9R0qPbtBPFnx/LNHraPJdPj+QsVueM
rybU/Pvf9dYHs+ic1BfehHiaU1QTrln6Y9cTVF8zl51HVlvFj0PppPlId964lbD0
LBYhi21VJi//M0Hq9O7acRlAS+AViGEquHUVB8QaEFbAbFD23S/fjdHQWR6B51VB
20p484AinVuHJHXZs+Em52585+ERcGX8oXVMdSn28FQQiC0DzAWmAQLMuNZjYADx
JuOGXKDSihjnaq3Ex9nDmmvLakWBe67fI0FgjPzwRghAHWl6s9Xhluduo8OuzTHn
EA83TCeJY8PTUU0hZ4Bo3/xgmISp9n4z/2Itztdxw6a7ZjOOU22RolchjV13R6n6
H8fi1f6yVwTYvHKuA59tKxGsnAk+6sCFSqPqqjAmpNanhQstp97YPjGAySfbAXxO
Qqd1hepojZ+F+eCgqAp4XyCT7WcuOP25cbKHSMOdOdpmZ4HorHrLQRUx21dbTMPE
eYJUdNdoqmWeksjTA3Q9YWPWIS+v+jcV1GaWY6yMjajf0icqUWl3Z7zuI3r7Yy3E
Q4Nw5AOc1CrsyaIXRGXfFf+DwsztKThM4znwhf7VWMdBvGZ/CsBEp+S4XO3LwJ9s
LDm2lbp7aNOpuHF+bkwBWx4cnV0P/3uRhTD68x0qbNqtbm9dwVoWVEfDLizy+N32
YVMUQcTEY3r+zgXXbMqUmSBXB3cKIaWMtRnBl7XTHAx9Jvj/Jg/bjsU44j42bTwh
AqAGT3eBWaITluZ8Yegj6BTPiiqwLovTfn6h4kxhludphxycIooWxrT5o5/kJN7t
ZEhLU4AmSA1FopRVFhMRisQroluKUaIkDKy9BWYjw5QsVhtJkTaD91pGNdiIb1sT
lSL5qi9tGl4fRTd9vn8GY1qsrFWTs5k3x2Ty1xIjcnVhUo7jPdXGuyDH4HeZ8NsX
qT9GTp8hiEqi+VWXJuDPmhCQvDFSJbe3z1T58YHKiGqbAc400yi9/f2WolnIB1cM
3/QISf1KKZRW2JVWBkj124r/Pt22htX5ouiG8OGdhBdwzFMJPbOZ967LrVuv09Wz
zano6tvTuWAorE7wkkjsRydjfp9xyqGd3vpaYfhRt7IJ1sXm9WMcGwe8T5qTKQvx
XfXdfwHVR1W1AIUi/IDpq2RsO/V4OX+qTDFEfwd5De5n+pAKWKRn82SIhOWIToJE
bZTxUNr+8WFjWZaPVemGQ8svavk0g06eL6c4Xw4vOqKebsdZEIIU6BFW7pDRX4r/
amYzEN9PciygCWyVY3wDVws1QsNacsViiIqMWWsPLpa/hRwQB57NDJpsEQSnhQv9
yviIO//6yeuu+wXBrlno+AqnGYSAo8+4aEQVlPZI0lVduPiqQdz8ZFSWlEO3h++S
9vxeZJmUBhJn2DXwb6lweOZTVfDeg9Yq+nVGAZM+i50j1u5Nsh81NBhVsE0eoUyP
qnuEYMWDlI06n/y9R4hqJ/CcU33DmD0seMLgy6es7NrLZzMfmmtsiv1vnHps0z00
eOVle8tscJmJmgAugpetzYmhf1+uNsLm6cucurAecO+K6gVTdC4oMf2GtNUURUk7
tWamaDHeE7QPgosp67Hxxlhn0r39jBh9Vw3Y/5XZ568qs7ai70VziUxbQGlEZQ6j
t6HZu/3WCoVyVDEDPqQL7mHp17om7Ww1fXp4KxjkZCLa2jkl/uU06NUn9WjbG2ix
cMgcW4xJjuBayq+YvJ4LicCqIZG8+8NHMgsL4PTfO9cBNam8EOcSuDd9mZWodjrQ
QUHLRGWfi67IAY975JnpsHXGo3QlSp8pU0MKFqgl7ub/delLLUhvq0tiDBHgj263
bjqRVHqwJm0BcRiPcLf52vwzmy8xKsj5YFL98k1x2KEHNDMUobR0GELzv1WmNQ+E
UaZ+21Cs1tX06Uzn7i8Y4RHfdxo46y2aVDZReo5nKs9Mgjo/pHLNFiYeIDtoyE36
hVXfw6t0GV9fT4uTGKdHnooNC3eyVTxduf9YAHoonJnTWQnudHRqHhf9FDpRqQNo
KbDsxQRp7AfmQqH/D59S70OHAyA6YGRIPTRqAZq1yBuLA5+/2pERXn7hLAw6DwFQ
j4lQqOyt4J1jGHuCeEc7v/gcv4j0dDT0UUuLfLALTXBS9g1CdeU6gX1vQVXp/GT2
RgfuS/hhVFgsnokheGIOW57AQDVOeAxy9tVi50u24s1awCh/K6oyYZgFmw8ZNe4P
30IN5CuSJ8sisUzDsREJfmfNPGi8FqjkLCnUOegvVzm93r9dYHBU/TPg+8AujC8a
JZjZsTKIGBN6jBl3GUpJvZRhB5hEV5C9qNxwX5q8xEapbe+211aiMeix17jCjrO6
uSEOM5yvATy9YycpogLUx9rc+1X7cTiE/3/J9ueoPp/WVZGN6+zug5+M/ANsgXtj
uJ0Wyf/Hw2sNJ2Eu8r8GzkZQks3lYlMakPMYV2rPAuILqGZDg0v+D5ihftbpoyk4
OiVquFunCbTTtCN6AY40OFvTpavFJLGP3cKCXwC2VWlOCdD8S+0BUzDQyc+OpC7s
HeyIT8hPoBf8pbIorZrdMDGFaNN1UlnP14RqUEA4JKJ5i+dD8wxSGT0sDlRcp339
eXgQZAulU2ZJwF1fMmTVZZevAhBRVPLs2C90BFXNVbLV3DKzka7uznhanqSL9Mit
TOOTm36KeGGYBjClDGuLtoq1tVlXgLThWkQtkkZ1p7ez6DLF8zFCn6yFcCqh9jJI
ztXInmGG5zQvm4mlyU6mjDvjNPGNowpD0XOKELqTsBLSgJ8xzjWWs+zVegQh61Ex
GHCzUYoHemHwtFohXenxfzvcXI3cZ4Dwqq+tQhEtG5f8Ys9PnKdI2E8qu/2LFkfD
jO/nGKYlMbrdqEljuc4zzUWf5FDgfoem3xUCpVtbS9uaaImWh4PsFdZ2h5hSq41Q
ROS04Dkbo8DUsvVQ/Ne925yfir89+kznKRp8MDZFXPnM31+wGfqH1JGCT8skct5Q
/lKHOHoeCvSiAB1dfZxxHf5h8rmh3Jrp7Wny4m2S4/Neu/eWv+Vra94FLuJfPBsY
EvTOXUvkNKSmAwL50DOQErH8Di1d5FYwaTYMgaQlEcYwIYhnsIbcMps+aJIb6qYh
taEv/44yE1Z1Uj7fKSeokpuUrRzt1hB89NBpOLHS66HBd/1lV7NRhMgnLZtt7+By
RobbuaXNtnQwfHOSZx+aikrYbxeQyot0ihITGKIxcSA6B+00NS8WUfc2EoItmPus
/qHvV6F0nPS//ksN1P/6uUSgExUdZ3Tzmr85q2y2hIPQB1NKkM0nYmF6+oq7x5p8
kDj8iUOBtJWES3k24VYFtHu1nQv38OqzptJ+3YbC/AKzfVxjwpoVIcALQjsAobe+
FKNvy0MxRQtYkMGFZwsOMAi1Ktiy2bQDkCUclLL31sX5Av060Atap36yM5xCCdml
iPha7JOSoZ6/TXofrlj8wLr/Z4YbpubL+lWtanhQdMATkx2z1VY7k8/L6cBxETUQ
wMrz5sy6xUHYzlnAWUiEFu1zqpJSTvOJpYurjkkrEOTxMRu6zeffIiJMOQ2RCYLi
BGyRwTYobwd2DiojkXC9/GTFW5bVS5pAFBOYLk0kZ2HT3Aizi7dPO5Ij4irf44GI
P8AZmXJ0LNTuMsaLPMVpp5Vht3HQKXSvzmNEVFXJVNLH3s4UmSrsKq09Q8TcUwCG
VvgHO0cjRF+N2vFDYHnfRnAKijgpFQXJJ8hsoWoGICcpbyoZ6puMe/nhVKDOA/2e
v+A9tfhtVIyRytL7LKwLEVN5uxDkqNq4sXFGSWCovByQbuKeyBz7noEDuPFKEkCT
NoApgzniitBb+kdoMNSD6nbp81+ozqIbVrVEZXlOH4C/0R8+uUSqDPjGKTyev+cR
/FOE3ulIedTWJsb3Fpor6L6LJwHcIFACbmpurWnsntpngLFUZ/v6DMH3g2/Cjg4I
16sY19pZKPiCErQvCiz79WgArB+ocJOJHpy7sX15ShRmPlrD87vHcKMNO6Dat1Ri
IqmWj9sKtGMtioIaUa2j6z8XczhJ5S6rbkZc5Oi2yaDNNhTlcMX3hS9JkJYS8BjN
FRmIe2lYgO7Qb7nQdi2GN5V7YuCiULZJmjoyeCswKxS4MWqrcddMh/hQx6DNftIr
poIT2QbIDZuRbLVhGwGjDUnRbWdiNV6W4PTQ4vVStup3+CetKGhnfSeMYMhygFeP
KN1zuvO0zX3RKMy1EmcCVPTHGHFM8nXZ6IKqypfbrLCqrI8VGNhtWy5pw4hS/wCM
rgRDA95CwR0/bdqeJ8HUXVcsLnPAg907wKDy12ba8QARt6R/bHanzrQNE4LtxAsy
LpwLrubG4TucWYmVXVPPSPZ71NNnpntyvGzWXXPV3Nn8ga6jBbR09k2MmXQqC10p
6FtCAJrWUBV6k0t3WWufEpYoNrvIx+tqZgbf/IKy3nP93GGxhIrQK9/ha50WpaO9
eT9SDHHmShmMKe9Hr5+mpyqdasJzNDGgO6GO4EJQJ6Pbrtz2qhyT1ZOfui99nhuG
SojfMkO8a/eWWu46ogO/o6lsFbI+3+1ps7tN5txjTj00soI+ggyefWU5WF9nrqou
ZUobR48DEuexklIxAVt/v2rPxNOx5/3ccLhBHL1CxOdDJixLC8NtbKEKlIbphIb2
7MNEJNRa0JfgHbRvskdNSsYK3B+4u50w8rTYPFFeUkseQmUigDlUe4GeOBT0GmSC
KhNOnkMbEBu8qaBSBjs7WKPIqyP9Ffmk2Mu0CISfB4uJp0kSxKkXPX0f0EnStlh5
SiPQuWhJzno7QjKXC09D7ocFahtJle1HoEB2WoWsvHz+9eGxLAg+IVhPSK1NpAlV
B5/hBRmSsw/r5xCoGHKyXMXtiAVBY3KdAIv8b3qYjr/UgxByY/u79BwNHIVqbfl/
qnkxlMtz2dj/cZTTZCYrxhS4qL63SivXsmZWIdtd1LaNVJhimpnAO+LWHbjHH3Rm
HJh/XN+QcuJQ1SPIJ6S7mNK3aYQ/naMfZ9c6F/f8v5oPf/ZPy2oSy+h7Rdwyiv9y
0Ch6WINZmG8cRV0UXAZimIbGIJ8u6u+zSzKSg7lrXTbI4l2RbpXgzTE0YyTJgC2M
TveNnpGBlQGUXt6O8A8lf753BjIXZYW1bzaSlT3lplHB0Ia7DJ2IcatLJGnsNBnq
jNuQjaIMn/zrIGXVmjLhp2v1227E1qYwyCH1xpstY2kuicv0M+NEZfowZow4okuK
hRSkLYbMVmSFpb4Uejwf2/MAwEaWRe+LIJeNT+RHEsqlKwdUCF4wywaAxCEpmOr8
TF2ER+IGBB8TTqYBRz30hiJowKi3UWv8na8zLzBguLtftTOsABOcnVFJl5a89scm
6vpNjY48bqw4qDt0Cj9K3Dq6fUg1/1kxRdHGlwbbhiSu4KL2q9RVsvayhy/4NRBZ
nm5cKhZwwq//0gmFu/+UaNWZ97wXocF8+IrAHbfANNeLtAOj/VMrS4sM1n9Cv/Tb
Fb/CYX4J7WwI1+Wf+CA8zDRHs1A67q1NUKi3a1CYwoEps0ggYmjrGjp13GGCR9W+
mIlAMOWRBpnt/7bomNV0VR3LDK9ktArOyOBiXBUXODej5R2OFYgMNlzMvPIlczdJ
O8Dun4MSFHF5WAa/0yMIfcrcMbXIb3wFWixdYr/7ytd6CdtnWdBxSaDpwt90htjy
0Yg6g/IBgL5WzX68cNtMFdrLQsJrwwnDqSDSzQfNqnJ9ZvbaCaCGja6RUlgnYoiz
NeS3ZyzGJrudbvv3CyVWO2duzaEOfCkDh4J8Kx2tXZY8XYdCj6+W6WBEr7co+/Sq
q2gI5H7HHdYGsKh4wc/McPaGSYnbW1fJVa174Zmcr0pTZxYgoaCrsRyXx5mK+oxJ
ugcWrfldSaSoChbJekiVYWSmPn+6RyzCzOB3/J5PdXTjM78NuvS0wkY8k/zVCldF
v93IBUCcC9SAdibu3qsJLMBwp5wMIQSwdEcanWcO8GKRhyF1//cKl2q+l05ZfVKL
wf+Ws45E8/jDlNgC1YIM29xbB9jZI51SI6C3LQv3MXwKqwch6nsP4+t2QLtQTqfl
0Koe9f2jUwxPCRGDrH/rae8YA5jFlmiD5kDVJKuzy+RVuj/dUh0dAaZKKUBMmN7S
9U29lKydxDtdeuLwV3Q18oZO8l/57kYhxa4qfrCTPRf7EMXWe9761L9bceRkeecy
kOfkucNCD5iDmsBrslW/gXSaJOoQKp4TsVe6XwtmmDuILiVViRDQf5M2ILu81AYD
PlXMotLTAV5/tPxmnfB9rWpSNZj4TCqfjSeWez9FLUDpyvs7qMXg+O4DU0Dybp2k
iqMyshdcCeV9IyDnzK4ANPmLxbCA9QpNCqHzC5aV7VcMzd4AJW1PBS7bQgzIrhr3
n0Sn6iaL4OTxyGKA2o45wFgByxfCBMlKZyFfDaYWfcwwAL0f4ubZ/WGcxGyJInpb
RU9m7K7XfOTPiynNrPK6qJE4BEk+4Unu5d/foZ+DwzkhdMGSGnSiQrwbNrm0Dpee
Q6XZmUPLGOvB08IaYW3a/CgfwUlkZ0TdkUeP3Hpzt16OkIOsg8c1J0WP3d0rV1qM
CIDKQ3+YK1eBHVNw/n81npLFGlmGHFZtlPV/kUUwoRxoA2/rvCD3ZTXbe0qdS1pz
M/c8avF5TnY9Px+EJ4wkHPckx5+BRoM6fnUXKmOFxfdocaDa3xvgeLO6T6HNhKw6
gW0fVkooU8zw6j0cqLQSa+wEKT7FY9+sp/oMmTumpRP4K8LqtWXfH6jwTZ60NHo8
R3oxoulmsE+vfR7XziQnlqap9qPXpvNnW4V8H79UDJlK9tx2fRb+ONdPEI29e1am
h3GzTw8A0t1A96qHfHO2UXLQ17Ct+7Vi8V6zMWoEJfmRFwFRzV2M/NReSaTOR0WA
mfO6lW2JRXeq0bF3B2wPQsAHjDpyzlae5QkYPClh1bzrjyxS6W3RnuRm1ltP1ooT
04PzaYLt1fI7JxsGvVI3i18wuTU5uTWt47/th2qPiUPhdafBK2d4I/Pwtu+bMOCv
HnpvDfekRXJs7yUvSw+0d6znlOssfyaCwRDVGLJZsZdFMf7Z2e9ds1qiE0vnboIS
Z290aBcH8WG2V7O4kFX6XylEo0b4rjep0owf7vsa4AyX5DxqigSO1cuxA3YPJ0YD
BoVnjYDMBuB/dkN9wjsSZC2ojLHpopr+RJlcE4QRCgN0DwwDimTjad2OXFxPUdLM
l3QWz8JSC2TbofIiKZN+tbB1aYPWr8KyvfGUK7iIXTa8VHckrpjojojJWwQIjOOR
GykIbmNpejxCeZzSgloZVquEAbbAaehovANl3cJ1Nn3cQzQlPC7kJHnIQ5F6HX4W
dqRk/mtgAYtBAlQmvj2kCibGtVSdHMhOzQsI73ACIK0VvcRffPAO/9P1AQhblhAS
vFO+ChSmuwW1ZdaFQU810owtysRhqirKv7zb3Lv5L8ANcT4RefdMXFQRTvkpuOtq
My8mZ2CT8pjdkFFQRtUnvf36LI3k93YSOQU8H8rZiKHniPykSkv4Di+P2sjWhQwo
viguz8pEA6neU09sHOIefmubQsLR5NL/XraWrznLtuNUxzUghnzlk3v1mp1yhkVI
K/tEfdwOe4EYeWPbD3W8bkzCGZClAQWeVmolWrLk3myPtgB70RbH8/giB5EZtUQx
7kwVjiu1sqO+8VxNXPvd1w9Gbu4yODugm/gG4whfrnVBry8c6scjv4+To3N+gDzq
au+K9uY7GNXDs9VkT58Zs/h+faHPhXveSgsRIxyB93PNfyXnVDrpoM6I6o7d6WTW
vNV6vKl2Na9VWOVOGlZ/oXqQYU7A5ZLWWzN5J6PI9tubN5AGcK+DAe6lVI1p26AG
1imcqh5E0uNwcsE8pixlpKXlZlrTYkEZQNyrbGAspWwHdKwMoufCKpAEiBMex41J
S8hdVdPv8G7HH/4+r7XV6cLcaIcjNqX84tVRhrrXZCgy5gRQ8kEZxHeVeD69hVmd
uB1HRBDq7/VwV73qLvrcstVouNV53q+xaKRUZi42t/7hVHj/b00uLdiBpFT4TPj9
qw2XF3Dct3N2w2keuLKkH+va9XSg5hKWmalmKK8Vl3+H19XOQao6ubkAbCtiQ9kN
B+YptsXPWWZchEQnG/82sj/7PCsfoEIMdzDO4FwDP6U1I0kqWRNaXS/Cca1kRYjF
tbJtv2cgk1scs9n2vhkh4dGlCuVj3mT0v5PrpVYRctiX+WBBWT+UydczLfIzPClE
rLJamYli/WQ4Hjd8ZO6Udd3++Ty2pfYfZNM2GtxTXydnIQuETLGMXDHcRkBuNA2z
j//wlIRWAwaGrwf7EK91rUp4F3Wl0fUOhimMfvPv8hEPoGRSUn7ffhas683TDPGo
c4/RNrB3aGSCXzWfg33UUft8SGz8sg3HyHr6tWnODxA9zgBajzwR0k1mlLkSLc7E
gxWbEWQbP6M3yikXd/hHmhEjkaeu7pVq4tBtIohHjXSFDVyX4pa1Kfx4LoYpel/w
E03XHih20DreVngzPNEghYaZqydXFIjgtDbBrO4kJnM/2XqMgCrR37+KjpoGKmOR
7qDHM+XzWOmDVri9FdgXqkf7hOZ7rxIljwUwSXDbZMKTlbxLC+CJBXBARirWxxc3
rnA1/dfSAY+4Fz+ayw8HlL0T+WJMQPM3wyTGTsDL9H1boIasSocctNIoutYPrPTv
7h/BWoBULJQY/TTOZEGn9qF36kBx6ksglno7E6xqXftK1FbTnm9vSulBhzQyoCEy
lM9c9YwteQk0x7NWU1Nt68grQl7vbfPNkwaHQ5O0QVYeSythaf2K8dOd+SheWVUi
G2HplVFbGxRWSzq0p0AabnxjX82POyUXjLPnym+5pturrwqdHklCQSh0JTWe5ryT
LBVDI2HpZoAerOG3y+kI8QeXeq1JM1d/SlmnWKMmeOuX0I4YQwOkrKi8ClDBEwmu
sgtzGKsfrHjyp5SyaYtwk3+QO+kx8xRy8B53Xz73eK9RfYCYC5PBwHKhf2qO7FR9
zM8lyXUuBc2tgNlLpYM4esUztGUAXsNsIMCRV5vaa48okBEwPggE2uKObSZ2yuvX
yMvMalnJ6wk+SVrISGUo3OWk4KdPYizNbiAE9/4L3h3lR7Vn9QTMhOn/Z4PKZJfd
Ckf4HLIiYuEbzR6r4BLu80M7ozgDZKi/MUDN+rpJfoBB18hHZs58aXvIErtUVW3t
bQ+UudSiVMglZ2zl1b8e4XmZb3LQzjmmzWeTcZN6DyjTO6K3UVcR1leB2QE0vnrE
nhunTMOLqEXZ+kkeNqIpdnkbvfdEq1XyGo2pkAl5wAyH5+fEVzWJrVu7r5bwLKX3
0sPbCUTojajr2hMoZmuvX92k4kXu7+dbfSMTVBuqgPMRW6Z2BWhtx08VsweznCst
PZIA+SgJglvTW0N2Fsm1HKEIJEMZmWwraNutxqAWHm+NbXMJX5YtFvKPVVXEJm3C
6vC/QLbv5yrCUxEnqNebZ/Ut13dwLDF5YjhYhCF46a3XVVm02973bi3+8CpdRhgI
Mek62+6OjPbgdW1poq5egugUlDXkUROLXQfAU171iXoQKUP4VPZNR6DIgYWl00yK
kg9obJWITv5FckbA+e2hHGto/yQ0RNtpJOhikdoUaimVYGcHLxjaGP3v0CyRyAx0
MaQQ/p612HCf9J0h9x+OTEHTMCn3gI6Oqdb/1o8/okfhp9krm4Eibg8IgQiTDOgl
rRqAWbdZx859mqLC8LVdr4DQlWdmuHZ4FXZGKO3Vs1R/PtOv4zyYHNPS5WFwotB7
Gace1sRKhv0nrVRm0s0YAzAm3qnfHoQjDU+06urz4OLm+2/kIu5ZHw3xnz5sm0Wa
CrkReSAXY4u5NWtyqqjkq0oaRIJno3cyallfE6jSzNQLN3T+NVrrUVXQjMnyhG+V
V/wW7STgESLcVeUhwuciakRqbii3VpzLq6RB8+E+WSra5UWPKlz5cxMP7MlUrMgp
wJ4DpiIeDNZxu/npmlk3zKoQNv6nu9iLmmNfgbMKoze/2iNoTWjQkmGuhKkZbTPo
S/WPkVqhX0K4Rs/cf/wvJhcq/xxo5SC+nq/V3+HPnDECwZrVwZU4IUxHystDi+9+
mFOox5fWeGCwx3k6HjrDSV3xUniqjKKUCWMvWnWb9AdpoHFhT+LeqzFWGsWz/HLI
R5qyBGdh3R6l8JCKwu5Vmg3SCKZRP0AO05jltHUVJBz6I+9M0RgiMxdap5o6I2nW
wNBjY/EAqnqUiyp13WxyMaLz2a7E4zbeyrQEvqjY159Rnb13+DfJOe0ZTj6Wr5AK
noofAW3gByzBGhG92px0wHy4ksSGotzeVwolT3QK2WK569JVSrK4t+x581GKz9CQ
rXcSxCNEUZVqzq1xrXKvmrTDVJ0nBYGTKu04PEnHpkshRWzumC7y/ew7iH1JxwSu
2fTeUB+o7eMa41UCLR4fP4PF9/22lQg5yvE5hDdTD9Zb0dOqglDH+j/s26WZk4/1
wy81RIwIE8xLinIZzxuln5rBZp/9wRKsgi9Vt45AwmYr+Sg70JN5Rw3kbuzNfTDQ
ghgt+aLGOS8hlZsLG3WT6phfo4vhhJXamJHwBQ2mwFV457sH48/4XNtHyPwA3gol
BOwKfoRX1uF3P7YPhuiULmqW39vuZotTtCBOvDth4z1OPZB17qizgsZIlLdkxAPl
MZOAz2tg74qeuQeEwxYPBjnWKQTF6xb9bp5W8VWE5N3eiwPjnHze3uknCgEfPMNd
j99ULhnc5MakfirJNOoPm1qndjzrmXY0nFy09qwSX25zld69et6L3ryMdNUqS935
ViPwLvxX0X5sGd9gcgLuwfAL0pHxafv/2E/3ibKEtRYL7KUAKGMRyzibXo6UzLJO
LT62s4F/fuzKiTcwOpzxlFoGpinpshrowDrTaIY1NM1foAr+5qwxbi1vd5k3T8RR
4eBZW1bUE2fI4PSDp4Bph6nsXYeuI6WNndXrCpyrNUzxB/44uRXkkj0vJisA7Euf
xsbpzOKWoPhI+aJ6Ll1isoGEWP+yHmYnNxT539H0vsAcK8vVyTak75tdcB+OfexD
f3IXQAWsJZcaSSeiSGjGMfvR5PRRg812EZronAT5Of2jEbH9D8h+hsHgXxxP0ysX
0TrApkYnFyS6zDBgp1LlrzEcCNrV4xVz076cML8VMSUYWU1CutZROr2NGI0o34Mj
YL0/mBZLlenT3zsFWIhS7iC9MxQ5N//FT3xaYDAU9Jr8D3N9+kEYCTmzWIJ3/zcm
LCOvz7xiaPgRi1wajx0EQII9Q9QPaVzV7cFcIvwJGbl7Nw93vriAcoxBYastP518
KXOLl65+PfBXnZujfi/V6O0y9aktV3FufNPjPTE+eioO3dtiXUD3XUUZJm0q4eGd
NoE3Cc7BcaInj11iukntC2ukH4eVZEr0fCBgNtzxV4tilO8MEwVyh2uzrSefKhQk
37+R4s6v/dyrytpOktbZEJPZYs8z+iIZJMsVtuBRHhPg2chvAwIaxwTx7dLECjeM
aNYyE6TQdjTpTsBXgy0ll4R3vqeeHhyhB6mHtUw41PYSP/jUeEFG67jWZ7j13OKa
m0NnvieH2UgbKD7ZKpwLJwEfjngxSGEYN8OYT2FK9/iv/DE+xxUsVPZCDe4iCccC
RhOUkBJTlGX9FyjGpy4wtiyJb8OkEzufGhL7gqUPRHUHzHge/UVugYiOfL98cZK0
jq+pqDDfn7MMaXF+Yj4p6yq8rXXVUP3MNs3nHahofNL0AO+KbrNJ5tQ2HOUpCdhg
kT1jJRiABX/z9jjC4V91mtEf+kCoiTqci3hJRe9/mJ8mCKHRxBe1kYgMoYUEvF8g
EZ5IHysQlxEThYAfEdiPOBrG8CxZmMQw+myV4gMUzu0DAetYZnE5M4ivvsdPSTgd
btpupNzgUu3kL3yfYUzvnk6Op9efb92HaXm/xLk+QctUPyZAvc9qb1vLeebbyzWH
ADyVZkcSbXTypphEIkS/erFyJ3MSGEWrEtxup/khXN5hgDtznDoJYr5Jtp8j5lbN
cY4wR/9vH+I0HblEtAoThFevQJM8fHCYTrrI9TKMdN4WHNnlohHk4EPhwE30Yvog
jwBW2fTt3YxjGEBAUFlbQlHUwiGKuzBlJXHQEn50CXAf/UQkJFBnwVg4vTLt/s9E
uIzjASl5/IRf+2ob7MNV1XG7KTMmCgLBbebSRh6IaFRvnO4ZeGn6JG3Rc2m6VFRV
9xuuMke8ND1fJhzWj5o+E+/C3GF4eZpSBN8yjZPdPzJB7I8Km6iSgpcda7R8LgKf
oCcSFpEb2DOPfdHjk7LnEtWFgT7LM4eE30pX/f5uBWDVSAaK2htG1YPqGRAVj8NP
vGiWD/x/xOOeSocsGIJ4RnU+omtqmdWaNamBWQAoWlJxzWcKCoctVOpZ6w1n5tQX
RluXAo3Cw0paZmCpPbKlmYtH0s5PIoYl52xlKNzFFa0W7H3EkfGabeHN+ndxK0Mj
/K5hIYyGB7AW/Q11MqqYpOkAKvjY65JNjnYcyYLFk7My+GI70YGiml2o3y7kKqMz
hr9LzQLTJ3ZNX7mH+qs3kQGZGbduEjau2hBJhRWBv5pPHIjnI2qMuabmR4ud/sQD
5JqTJrtuFQQpvot0HIHEBT5o5AHFCkMqB1yON3aLF+j5sp1m46W03J9uaQifJETF
zGhkMgME8ELii/X5NP29aGvE6Z2yZZ+1WUk/WQ3d0YneE0jAu+KOmhuu7gFzOvEX
M11BgjolvCzo6xeYiSLeNsddGVGfMjcciT2fQcu3ui/tmKEAROL2uCkXfFdB530Y
4GDcUmxGEFZsWrUdRxFt4SK7e5bWDAFSJECknWj5TKhnsB/G6qgRF/EB5Q1UBJZr
w74nVEaReN9WgrTqDYwJjzhecZbyXtQO3aSJss7syfeKOuZqLExCRCOD1uvjZati
szCDNFUSurpj3RKvcruXC+AWjV53u5li48bmWt17nQrML0B/lnKTy3xBQ/eA1euF
rikTP7FPik7glMJPNvUYLgSQrH8CRxzGA1evwyU4KvHeLK0PczHz/m7i6na5DrQV
oqVFEf0sIbg5j7oGZtarwNm/SJJySBj5hu2BP8B6YoH6zCqHYrvB67keAOheNHpf
TK/B/Xj3DbS5+Cnol3BYY1RtUa6Ou9wHyolOX59v4ym09sBchLp4z8CZFSZaOFmu
q6idhcUm5r85cbSSkhN1d4N7o21fvgVPubj2UQAhHPz8pqZlTpQ5s4s8oH9cMPfD
T0cFOgFaHOcbkBiCJPvgB55G9IGXOMCHW5aT+JoXrg63Q7RLVcQu3HUkGL2g+o8u
lL+KCmaLc8AzOJ7sFIffrkFLYZo6oeSJeZU2m+etmoxCZNAi7QvfLb75i1cB/iFM
9zVH/smFMeM4zSpWJyWC8KD0LbIfiRj58z9aqjGIBSPZp0HQoNva9w2e26tFTsXt
WxO0i0PKCSWmGoS8HKIwAzZ+o52OeaKVCnV4Eif8dViN/AfXW/kklL8OCSOc7CSk
W0AHLZqcbgCgsCfoj4hd9lnYCXJBjUzK0ZAFJaM5OF+mBChHewcJu/kgR2VWoB+h
flo75BVmzUYmNrFC3IyRsyI8ojNu2HXjCRvSjEu160B1s9kcexV6sjIIXvI9VMBe
ncwX6zPqpZStv22Pch7YSnVgH0PK2F7DYmdWZKnQYwFUcMsHrS8mkilxeGVn2Tdg
S+fGLCyra95w2hNyPmPMsxZ/DJvF+oqZBhHxI0eFSd0FpSffuDshhHHuy6cRSDHh
PHh5mtv3lkIsUcvNDBUUzOfsP0avO4kkfogg1rv4Z3CvxYTjBoChgGKVZio7flJr
qJioRfZmgGOn1ij+HDpXKXDC/ZJzRj1oVW5Q9NuItEqf7uV85YqfyAVg3JjJr1Ix
frF1yU3oj+oWvs25sFKIF9902meXs+M1agItDgJ2keey/saEw+8dSlqm7OX0cxA8
gtEDDWVPdK8+65GV7YlCXoSvGKvcdix2R22oLZjK0UFI1QFtVdatn+a/Dx+6SkfD
+dwvkidCOHmAatM+YBcaFE9cSFap1mpxzeJOfIG7kt+karWsoIft6eXifBVPrc7F
7jV7U+kvQrRp06ewDYmRfM80sd7zhvIStHG3zNkJpHn5dOHNAeoX3w/YR9oOBRNW
fy/2RRcdGERTlrjphkZPahvukvJiEQa/0bLnU/1hLIf0pBeEVI88jzL25zznieQY
85BkEyowk9VynGbqBEgYptmjEiccIu8RhD3KZfSnfNmml6U6KV1sMmALgK8u7BFC
i1BNxPDxNsLM1t3iwvMyiyBEFCVt/Am6QaZ+/zb6FWe02YtxK01aAXIK5Cp3PC+k
KFoDnT6arwKPZ6vDsuSa3wbJxr4qOCtSwiv60sPUEBGB14x1Fd9G9zDGdtfruBwC
CbZEz34ylq3HHZ4MdpcBbCAX4IoAayScREjhhimsHGrS1E3KcEMwQYQmaE2ky1qX
Sych9m0LRmATGSneefgv1z/0Es0NS39GpRU1otHOOzUw3Eis7LktnXSpFRnJwMY4
YvnxNRYzBGhd0cTBiyh6Z0qcgxQD7tYlCMFXI6uIYOiCstpgH9MgLyT9LQUW3oDo
hA7PNiejf7QGiPMNK4kGhjQd9PS/VSPxMB9QWx4FE2qx4JE5xLmvBXeKEttmp81F
ivzWAF9wwTmyhBkbVFqp6II/2VPPyhwhwCuRZoSXVXxP9MZpUzGuaDY6THSPCJ3d
l22aQ8m8YXxxpLbTJrKRFDGNeRqzKhda/x7NLnYor4w4SzKljD1jMN6tKa0VMhft
udyHsFZA/2kKcWTTojBNJqhGPi08cDI99MPKO7iv0D7nXDxZlZEXgXDkmaBCIxKt
O75O6jWP3LJq29s7UcvnUjrX+mUJPYexMb4BIuGAbmA3by0Eo46umQD0nbOgdykG
PUTj23qSkYW5BSta4PGAPacUbJ90bigo/nynV+jJiU1vWi5ip5+7n0AWDnW43Sjx
QV96CTx915eF783/mfXgZVxW+NPJ4E83lIg9O3uJSQUQ538xuOxcUPP1wLQaaMKv
hXaUsJTm9uR6m8PtwaAR6RZb3/9j1/+bhndiYIiMLpC4KlGz2jAenlJkX05iNXSQ
tSKkoIZDB47WYnRdZtvuOREyJaKmD9EU9vv/JgKW/AgCa38InbfsgXzTvixf5/gf
tX/7r58hzbaw4Bs0cscvwB7Jjb+OCKV1HklPXYHel6I2athTUOVNF6TqW5F4gbJw
YS7ZcoqVEgfajf8nSVzI3giOoshJpwV8hFPR+09gDzjlajKusqADUTXmvv1+Fqt2
s41TMZ/jAFZ8s1IzIt8qCVmDmvRq1C+onGDU4BZ52Iuw3IBbQ1pmvWJe65zFKEeu
Y3tA60nj1Pk1PRuNWFJPWjyh3j66ntdAeQY/EAzmYO7iBc5YRwUt92Y8+YWifKO0
KvrYQnl1YrhkD0LttchCHMT5Lqz/2M8Ilh8UVTGaS+OF25ZujTHAVSYChHCFdEkR
HgYKMp4pAr6N231nG8mrQacjmxDkwC+/upjCK3AVHTjSQH0zcJCc1Snk1xhpNNCW
KNDpKxM6kgzLTPElARaJnMJOHDX2+pFasbejiMhKpg0Xk4B3tLlqPNuY5enn1RGX
N+edlJcUE5hlEWd2/o2AoQ4oriVOGvX+L1g6R3YQRcJj6A1GCKB/rizrFqu33rgA
ZPTic7bRkKbygGjt1XCXjau4o+PIaoIQyczbuxfPTPBf5dcd4ZU63uvIoJ9+bMsC
qqSuLX9yx9DmWGrK9OAE3I1/sRj/qRI7DAzPaFh3hqNNg+r5Qc191zNDxey4fb/M
jPczPmUldN4GmwMWWP2exJ4Js9P5D4Vw7MFS5y9Y4tJWk5dXlpHfHH2nn5iqPmae
uXcSyR8ittQTT9TWandMCfvjaCQc9WU7Adeq0QxnwOwyCWgigyANMPWsmo2F4tHE
1SB8CMUkxq8YeQT9PzLdcjOtd2tUIDViyRksUH1xYU7ZmxsfeRt1HdYSCVe4HYAD
Acatd4QBobMBx6XTFqSL0UztDMQsYVpTwVM9v+9PKFPwvNHT66l8XFpymbrsxhSO
M/0ZGSdBy7JpFZ7BH9ODLqMeONaUO+CdyEorgkx/rbbzbZetJEKO2vIh6x4jts5W
zooQnxJ2OSYZSbrAlMiHRdf2u+ujBN9uubfNyKeeHrF51aHV7p7I0Z/Ix0qhiv8Q
dWX0fNNzP4E9CfD/dw2gloHd1cupGktjISmS2PE3ewwYecVROt0zf5YZPBbqyzuf
xOfIYLi1ejLgiwTcGAab+pKQb/EwfFq6MdMgoJpOjxDtNhP/t9eRFzkGQQCU3k9k
R+UYsMgPk9boVw2msUhQ+tgyqlEEGUdYri39iahRxT+nc1E6OZadx7rUkEvb4at/
ENVaFifAXW1fViSw9vlENtGp1zDyQi+WtJ2nIu6JCBsQZ8O/jl6Cio277bIp3Vje
N3XdhvKM4kD/20fqquEiVSqzHgOuMw7iEIZm7B+UCWdyXB5PL0kx2RX1ZERf/ZiM
9QFgYUeJQtI3EXqlC8FzgJLSpYrwVIK3tuR2sriZNdjT0CysGLzqJCiPqToyFOk7
d9DwZvwKcm+tNaPJVR5rGSz4dkztmYnA89EzSmDAw4aLjPf6UZNvfFVJ+p0AVgNO
Ho1Gw5sc1rEf87e0aMe6vZPLUP5t474CgvfWtrGpRxI0Q96c7WaqIG9wWS9aDxR+
nm6Mfq+2Eg/oaW9msBLKAxN50/W7BGs6QPGcPzxtjsIhH+bdMTiIOi4Ilv1ZosjU
cmoM7Buad068gUUCUDWpD1BMcQPDe72P711zXp1U074nHFOfDZ0Y6hcA+yikE37s
Wm/ESgdJ8UMlYq9Y7w00De85MYJsgUgC8RGRJoJkuLspK0UUi90Lb2AcAzHZCZNR
onuM54Je2/ic3poNUslhTXiPpuoMlSkuedrJwnoAOHMl9GtqjMjQo7AV1aeeOcdy
pjKvaf5rYTDaCo2CwPdIXm3kvhitIvkSaUSJzOntll0zlTjHNJul5WaijlWCJhEF
fydWFwOqdRG89XrcKukC8CFkGNmIuQ0Nen9kH9vcPTWnC4kB+06IPRbxunZtId0q
QzxLGgX30Xz3mS0z8xNX9eGGowXgQsLcXuxBXSZnRPCTdccvL/N0DNUG75ann9hU
GO/ueBkS2tb5boK+uxjfcjkRjcrcnS9cH/4wImlkHg7h2kbrXN4M6EdNwSLgVAdh
C/Ozaz5f/e+F6IUVO9Z938N9aVjm/W6N6LgLGqrFbTMtWZ16NzFgCSgWv7PBaYVY
UYGm2LAAMKJp8R6v/EG2CVP9g8/25Wfv78i2sI9ehuJgEzYoQLG3hJS61XPPMbOH
HvreFixlKwbBfdL+eT36OPvfitccySH7CSwRgYlGm93SePMwMRdEng1uXHSSdaBS
LvCxgUpTWnnqMQQi3ReLVfkw3zDvwN9kiCCAROl0DPBS4MlTfuWtNcuQv5xs+kmw
js4eefUGoZ0qaJn5wV6ykRK9/BN0r7oV553Tym8gcBtZAoFCY19/qlBFu2hvlZkz
/5aUPH8Om6sYJtIOZPdNakSJeySBrTQH+AXfQetUzr1Z6BfN85/OQDqe0WTf2NE1
BIf7dBtvVcZ6Zsb3u8DzI4HMi3xJdQeAUBB7qBYEnsgk0DS2XyMLrgvgEWVjxGg2
it0dMxO1jl4Eg8jLRpDxWftPPr3sev8W6ZJaWblGfs0KlTKzXfC5T0Pw11kYwP2k
RDS4x0IAls2H1veWWpGUS9oXHnlQ9B39HKPG7yP8jqVp+HlJ7gr+nMgSu+W9FfRf
KK+oB4ILM0hRsUg4t/NXkG9ppdoBF07Y6BQH5jiJbi7sH6EKyxJoEhxOLshXntI/
U6GHjjdtQ9J6kBLmfoSe0K+amyXaHzoLovzFWNhRF7aaTZmJjdr0giKlfJ+XbzaJ
Af2doEETeZc/5OFU3OR8jRFewu2n2HCwdjMg+AI1MipJ+PnnRhBuGbrfBawbAsvv
niEWJ+BGh+WCxJrlXKoJJq8s5ZBWxMa8orQZqvOLvnNWJCiNBU9Z70wq5hI4ZQXn
qNM5I/h6f9ONFyI4qj41fLZhEjksesmODLBnCkJhpMDv+auRCzT2oaknRGnQP206
VP0o7+lr9u+HfyDkyKcxp7fhKxj1QH0M+dhKObbHoMzXD0B8pJh/SqKoPj9dK3yj
DKqRMRvbQjmTCUzYN5/r7mczXmQReny3KWa9gBnh2Hqmy10tO9Tk/ZUDCYy4Ri4l
Gl7/QP5r8EqbPIq1ZSoe6p4RpXkAQhmDyf1bTGf+dht2u1/WK6C65hpTj3tYM3rZ
h2HyJce6KJOzSUyZ+71Mj0g2apOmD1UdxzblHoBL3rL4tbqxnKqee0nEFKerdbXd
yrtIEVuXZIpEnm3nqYLHQwLvOeuFAFLsQihFqtwhkzZksB2UMpnNFT/WSTFdBs6C
jJSuSpt+qTyspewruNrrAM6+tPElQbrUv6qLR9EcTLcCSMyeisJzW4dkr9A8465X
4kOu7UzGz4RW+NftigLyy4ZKsVq5PscjZmu1fZ6+8veAOqQcraD3LsuFzBrFMhkg
Y0GUy2c0UA/aRNu/rQGao0O9eZxrJYugtyG1ITH9p62qiXIG1mKZny4/zAXpE3v4
a1aJOM5w3jV7SJQ2YrJ9cS5Pn7nks8mPIbG+RC1FqUhp68r2+FMrrpntZqthsCbR
T/xeeh80Cn+zQFH+QdFTRMNBKIE3+EhwCdKTE3Lhm+nXomamVbNqadfxcLvbMAxh
axJlg1Gv+9TGN7EcL3DCmiYpilgoSeArO5wh4IdG3giNC08ctOwK08sc8f7pISL0
DrKrUp2kLwpOKdYupMZBcdH7tMZJ8VrMHXICHJnsr+1Je6wV0XXbCftNi+2KLbQF
sLAr6wuVSB9G5lVU5Xd7hYXeP+i/K/VyVqYktkIVISrttrUlRqbSmE5AIQJZbUvL
VdWQyzEHsHP8879LGDbDMZDDyCsMO6jOQCsPTbJk73UxZ/bmipODxlsHabcJr4iP
JJtiqOHKuQrmWmhQBRHqT4AUysGYUtJz/zHw/tNv1UmahjcSQJOL0ck6/Xq53Y04
f/RiDRZ2BHB/wBo3IcVl0Ha2gJpvf5vzZtUN310W+Qpecl/yu4D5RF3a1WsXrIIa
0CbY1LKvcLQ945ufgqgO+KyAI2MscHG/jmb/F7uUicyHPxHTGwH2lpPLsei7T+0i
FYqTBjdCUf/HHqZTxf3Nx1eueovisg/q/DlQ/DjeGxSJ4dseu05ZJjCVF7iZvAtx
fUgX4HrS/8Thop6nbTbZeZj+2VMK3hsPbmxbuI2BQajYm8G1TXO7tlYR3c+RnMMY
hVtJov9TxOBAUlWDXUfDqB6BdsJveBIIqyX7A25l/gzglDpDAxMuRjq/0s7Xmj4p
h2C02fDPqrdoH9vKsA/QonicqClU/OVDUts91BSSYQNADRbhKvBazu9pgBLjggT+
mRmypiQyY4vhoDeJDOD4nokcUZM170tfpOcRczIb9wudDyo/GBz7VBHbQmNGAokZ
lWdrtAURON3KMiWhV/taE0iNCkzvhnM7xuha9PqwyuX2C7TERBwRvIkXlAjtc+Tt
mP+TAUq45Xmo+IkRdud+QRFrTTxQ5vr3jobTcVLM4iQBjnTbXcHnpSM4mHgw/uLR
PX/gDvWSgsWS/P0f6J0SCJkSgSS7eXytiYnPM+qSldzD6da6vw0rpaERddt6tiyP
IE3lnVI+t8EfQWJRQD724bPhbf27+nEGXOI0LXFziCxK4TMEThsF8EtnjxuoOf/x
INpDYCMTepFenOG8RkfI1TCjHyms+2sIWftC1emKfBvTA8s03QDYT7r7iXX+AUzM
300YBPkn8Rs5+YdprxJF4s9Ze/jEMvyb2x8oTUWV3msOhfh6kaBAYGzUM9eO8pOr
jwNXtODXmGL4cmuMivzzHtIHmWhNAgbdcskov4D7d5senfl2eO2RVD4AyApaBrZ8
uXsIXDQuVTG6kJQnCWZndtUWD8VZr25yfNdQufS6C/C7nwP0XsEzGc86pZtg4/sU
J2SDfUatvUH+YOhc1CoFrd9oR4u65pwkNeZoUXfX03ITQyGT3knwVvxCi12DHMLn
C9S//Ht7yuu5cP7z5/Os1Zm60AOkwbAtWQtINejeYZ9o3JCPf547lyxbWdR35LAZ
KUOnM18pMATtOdP0soyiBeYmo+zgv3x4byJwn4+TClMNddbNiA+gBPygoMkaRZ/M
3yQbD8/Ze/bPQkidHrER+b3zAM9I0o7dF0/8oUKupWlfOjzRtPM04GC9057v+E9H
lLBwsMRY5obPiI6OyN1RzcZvcPkjg3G714Y0Sn/pKmNXvGS2JGTplVYTh6JNUrPy
Xn6K2nO21jKkakTxIjs1myGuQPY7BwD5ByVWpku0ar4rE7evB9M6jCcZY+1lIJS/
b+jUndOWsvjR2Yv2lBHsfWTY+AP8YSYpS02bKZG2zm6yZIz3QOrVT+aTxpHbL7wh
gCset8pIvczzPIggpjK5KDUBApvsWyv9eylCuTUSADTEKpASd/Tyu3EexXh0Fg4O
bt2CT5JQECrUCCIAEm9lz9Hy+L/Se1mUbFWxcwF60dGXIj6zL1VruUWs1S8va1Gq
WQKnJD0w3xCQ3nS3ks6xFeBKuhSbtAO+moAIMGhnUyYzUAu2bEvpW4qA6AXgGJJg
OxlINvhQiHn7n/DsAoa6PuHcteDqURXu+Nm7Oop1doWD3S5O4gvHq+g+cQQB9/Wi
hSLAKcfAnis+TU5XNaEymx/6z+Gwgdfh7qtYQeH5J6/rlJOqIOm3t9b/oBupqrO4
oNkyb1Cq4euDu46rFoRSJkflDAiRyue4Epa+NBcn1OKNIgLN8TT9ric1OEjY1VIL
dIoQ6Dv3uzn1shId/KgvBjdfHfvmdx9AvhVlNqbMx7Zbc3ae+jeEi+BSp2OMHQyi
haaxoih4UvuAXfrsR8f3eJVlRRmUwIRFi0/P8GSNt2Pc/2vrpUdIAjGzOORBRLLA
9AXI8KSNW7NMY0LySMAEZnTM/euPCR1uTyFgHezcXHkgEENQIv2eEn/FgzR/Bbw+
E9tOvOBy+BCt9siPdKgIHUZaPfpn8lyd0XosfB6MiVnSSWdyGTjMAjn4iZT6bTb9
9inNJeJcI7YOt7X8crnWIZWcsrsunndknBAhgTSaRJuT1e262LE90F96eJQ9RG4E
1mU0RucDf+1+GdYS84ggUMOKbFaN3HEh47VZHmZ3x+CWsVpH1e9nKo6Zi1KkV/Ai
p4jTsNN1yv/gIzTrLCe5tAIx/+ox2CsHTdZYlMHbeh6hu3dFKBIounDgS0PA8jfF
ysyNX6Sn6J2C/S02CVjPPVayjd4+lf1mGXCAA1Yd2ZHdmQKHQCOD6Ri+dCykp8/n
/u3vw8J6D5SYVgepXW1VvUs1PkYYGwpRGTrmN75FGVgb/vJTasCQuevyKODgs7Vt
5xitryQ5iHoPclxREbchjRiRKAFiv6Hdg6kmL6nkeEFJx+gjtheDFuSu+iJnWkUa
UTVs5BTKNXFa1jXGeAPGo7rjabcbMiRygOsG2aV3bl6jOggNRr6/N08AOKNi3BeW
7bku13v2VzAbbF4MiSp1kgqGls0BHWfdsl1rHxQZ9wV7ZGAwRwute2OiyWiwFxW7
SACzEAXKaeeXr/h2KbU6BnzavVaymfs6hs7KMJTwZ82lXXq7eBZB3xzSMDY17vaK
A2dqL/kDgWHYvk2ZevFD/uaqk+1MHccRNO9Wo3CVZSU94zvwIxZWiaNWL34ftdQb
3uXvHH61hwP67a4yMWY/0ivj7uwl1rQSgDdP+psxizghpc+FEbiNrQutHD/NYGBP
N1P7H9e1EnsmVoQ3yGrug8ZrK9ZEFKJT5g1uAAA8iHbWgWv4tofrbeg4iCRmNPxr
8lmmcfgDR4pjUKsYXhbhbVS4Lxg8lrL65yNdYz7El+6NbIion9Y40aKwtF4J/b4/
cirjHlaGyBaEGtWM/AscEdGKRGHUEoTaKA8SErYNm0eFHQXaVCHomHFAnABT9yNv
ILXmIrGzfaC4HK0Zzoo8cg1R5jjmxVqYjoHmWm9qxU7RYHil2Bu+H3sf6SRe7d+i
e2NjDJmKnkNOXbloYnGXW8xKAvld4MjeEwgGO6eqFAp1Y6B3OFgu8JRpzBSFX41Y
Ky0BFlhVFjcOVfII0zvMvt53sWUmGHBXTgKCzdwADqb25V4UJRvNIk+xI5PNkCT2
eTBQpUOOB/7M97AyshET8qG+NLwCcuODz71BaNY2AGXNnJDt1/vKa9Y9werXIKn5
SmDuy6zoUYjlFa9d3PhyNQ3QFsK9nj6O1AZVeEa03EUJc4BYr0Sc02ykM4vS1pln
2+gGJLbVgjAoOQkLa9y+NmLikcKM9IzPGhV1PaFAu7nn1kYeBrSklvmd/sq2TJHZ
XK3d96+5SGO9ZtFPG4eEnOldXmQUy1tv5FPUaBrM2UrS71Kj3HKYEBrcJVaFXN+E
zuW1JijvCRt5f6cjGydGGOhQThrDJZpE962vs4hbdZCa725INZYBcXMKU1zp7yC8
xLZPhvfZgIjafIzkfdEuYigHoiI3Q2QDqbJHyyRnldVXNqgxx+WZtC+Bql2AMLAt
Z/Z4ergkAMQXY3P6h/P4TS/GaxfSmgDvL8JAYjFMBg69iH8/AHSUHcVu0cCRunWI
glL/uZvScR1iuXJfrgr7ljuj1UYct9eGtU48ozA3d/TbFXRFbV5WcsiaXDJ/hHFb
szjKkUhTGnc6WlKR5ZfsD7Q1rVKCwv6V9IWzRU/FDv1PAAXjBJejOjU7Up8hSlXP
bV1cFOmZsz22k3J3TtYOutZ82B66j0hbfMOnmPJKzxdUKetIfdWe48u7rQvR0wrO
YJiQCK3TuxRfwO99Cklu9iL6OHhSq6MIV08fUC0MvU1re4JD8zHi/Q9pN7qLP4tg
Ye83LqP2ATOCO7EaRNZi895k0qS0n7xiFQA/s3hBldMiziVI+tdbjanyRnEFGGTq
zl2dgzHKKOuY9V1O0DY6JdC2D1Rtxnm1g1O5ACq8TGrPcB5NXMxCe7KPltdJbOgi
8z50mn1HhnfJ3rNr2txZdS8Kq1Q+rnIcGEqmAAYhiPGhbMHBL0bSLGs+RldjYGvL
qbo7UEHtsrlOzujE/D/uB7waQRvG6U8Q2496fLmCGXlppD9Q7Yh1LoZukEEPsCqV
sSLUfdFEsN8JBjuZRAvqBviI4ooZ/gN4W94FixfcvP3P+0CenL8DhGbDDToCyR3X
/TLhN7XUanEQLTPF56UnFhSGkxZiqdVhwVrmfc7XeHDPR9vjMUgkl+p7ObP4MRV/
ExyG523hIhKOXY7XIjZg4OBJgaktsG4dP443srByzbWWnoSm//TPceo9yFQ4V6jk
Wo5MTEIU82mT6ZiOcVmDEn627D+uFLHlVPZKp3OQPzVT9BloPZbIlB83+4m1dib3
ZCqXmW9bK0h7blb9cN8Y2RnmYyCRc8WlbU6jIWqobdoV1Yuq15d0AcB+Z4fKZTly
/rK38m7foaBmSf+LraaDdgwAccT48nerABZzjp5bUr8qT8ALD4zwzANHiwQsMaXH
WX92EPPSHuqw71bQ3PTpObsCfEn58/UO5buqAC2dZ8YaAToSg1ehNPG0ZjC98R4a
+jtzewhNso6gax1326114fdvRHXszZkpL8zoWgQFcqE1Fm5av8vL6IictzjEshGC
t2brrgFn67agu26kjV1fBrxyra+DsRh3+T+g9l+I76U4gZ1TsU8tIrxHm/TY4KZB
6yEy8xxu4DsjmjIsxFJUCvNItQARO/Mfx0bXZyYdfrD4xYDB9OivVnja0G5pDEIU
yLoZZArr0nx1jHKCwuSmA9fnpmjA/T4ajt+nSLKVZkB6euKazKhsL+lLb53AVPI6
8kHaimLIklUn5LpXN9Pygazx9he9SWFKKLQYeURmHnLS/nvW7rjcyMX3WObkkj7d
DrjoVGm5fexVM5gQRZUSwm0svvvYS3oJH/FwylWpooPdiWQP0S47qRX4qfmvQFgD
guAXQXUzXi+QsoSPogJpQTG0EhjkTyrm7goqU3Vq9A50rDS39OkfafFTRAgJofFk
Bsd/yrS0u7/jrz83AmC4BSu0DM2XvaFjWl3URd3UwmuFztJb7TSw/hQ/O14Mt7hL
6T87rX1B2mb8Dh6WxP1JRzzVeB5iWeOVmVW2J79OOFDjTqRRJl2skurHlcvervcm
dtHG7sKCS0ZLPQsPMp8MMddYBxhJUJUOieOTiF7ybcby6cY/i1b90epqcHHx7yJv
RbprtrIgrDvc0WpeTVATRToO3RGEdVh3i0EK3WM5n8/lAkKaQSLAv0dHmCpXVyRz
9xzqUltn+aRiaP5GGPpn/iQJREORUpwFNJYYzMRcBNGppFpWW1ZyRC0BjQ5xF77s
oSMTgrbEKCuqEkdwFs/6aQH5RMvoWqbo3f6IVv747GYZCZuVj5Yd3bhwQjLu5m4d
lAFEVhpY3cZE0h43Dl1a8J6ye/u09L1FSrYhT6oYF0SDQyvDPpC1MZ0mECwwQmsy
7bxf20Pb/BVPNQPU2H7p/c2Pb8YTrc7Lhki0/+CXz4FTUA3Svgd5oH08hJzvjW5E
wor/+Wl6BgBBveS1NK43phjdhTcI52guP69z0KyZhcGf1uUhiCfFYOd18hLA69LI
x2jX95AbnGv40/hP5tIDXyeSgm2eGLTv/JlTmFJFKz0EvHR1XRLawg0wxh6cF4jm
cfQ2KgFyiD8IIATgwTE9kA1aL3qXi7UbVfAvOB5IOFijMFBbYPwCykYlfNiiBlDA
XbXbD1qPTvzdHnBUo++0iNZ/B3AsdHKCazqwv8L49vNyNHvik+TUZ+mrpPrRNjE/
5EI/n8u1h2vi9NsmDmMjh+UbGIWcos7nL8QVZkqS/C1nMmpxwa9oQ6hD4hNcHwu0
2WMbR+FgBmn7ylSVmAx8IYkX1dq8XI66UOHQw6EtvhX3hylXNAl+M8WFfCgv0LUf
ZQBMV4sv9qiNeoo3lUVzFAtzkY6JCTI2RlcgttfhN4J1LdMIs8FTtSkmdEEJhUoi
YKf70zuaf5j4TA6N5zULAGwaIYf6e9S8hzQN6V/I0cX23z66rt1er34abUFJQsuj
UooR1JmJTYD5YIOF430p9QoS5xgd9CTUGRiPPElkpOVQ7Q3smJaPwbnKScXQMNay
DDfiSq61u6oHW9Fc1YEJa/U67QrRYb7PYX/OGiiONUNy2L0nVceBiq0qIo7rqlk8
uB6H9fNKBY/+111kahReJ/QhUfo7zmbzQEuPuNKIN+NFFEXVK6o14yQYSCG5/OCR
2iy8hiwKZyx72y31kICqP0Mbq2nri0a0zi7lK2alKW2xukT5Kt4Suq95+4ba6LJK
MpkgIw444j/8MUVBWYchequH5J9UgXceNzkr+BS8u0zuUXuMxIed9FA6gOXBY1Dm
Ui1Ma2By7+5a3rNBzmWCNVMeNj4mDzAOYgNxcB+3hyiDB9lJGK8hON0vpMY5z//8
omhd1QzVBpp9hkjwfde8su/8ZGYW5XupAHK2IullKpLEIJBk4nXOY1eSdeB7Kd3C
4x0wLvUoO0KSTJq6NRFlmYXukFhvamxGahOlF8fJIDQgLzI4uzGT+fK5yvFiPRok
LpjRAuPWcpyWay8dyuKXCvyPAeKl0eYxF1bk0rRS4xI+o6ciduQ/mNsGrFocNffA
ylwGOfRZ4HfLaSB9XDQCFGWx7YXFm8tE30PBNlbMyfT1S+4HN1PakbNGkxAOPPdv
/cJjL9QPHImpgd/6qSVSZDcgkmuHld2PI/MFeo3nimY9+MsEzPzcKcaMCtW9/XhW
secwUWe52v43Wney9RFsGMINU51oAn50Wtej5nZwB4DDToBu2czXOJQ1FP73toAA
iE35CBRdME9xCbjWz8tU8DbijXDEL8e+2ubJyHqoG3bctU9fu/bpDgaRI8dPO2tp
lNXMfTojEGSBQsUFXjKfMIg4T5Ke84Qqh2ChFn6jIt9/cuefKGtWctI/9VAnDoGw
YVthwA+RrQNYKOIKGYFBfBKQnIgZYlSEMYbolzintoMawqHF+ORdYLfxOmFTudQS
c2zZfNNfBZUL/0Y4c70EduF5T8907WqIWKqodC69ot1YmWYjtaDgP/BMsszBuWBH
eOyZE92WDGDLXy4G6Vlm5cKj6ZsTuapRDbgRO6TvvD3d7Fn5j4vPQMdiVT0SF5/s
7aHWIX8g6eIsz+Hqn76c8XiRuvjbAi9hdXmP5XOxCZkN7y4yk24y1QXyHlI2ZsQ3
QQ81uiNCNh3LbC50RuZ9Q4wqDT3IPERVl5YqpFSmuj1fnOs+lYo6izGsNkuajCvO
DG9rez7vT32pm4v8W2cKkIBOPUoBzJI3LGR8xV8UxpkrOo8as/SrfhqhdOU3BFFq
TLO8fTYdYfPHYWw6+sDJmzEMVYOK3y/w8InQb5njEsENJ7YUxh45FW7N+DzLuXG8
ASL7ZyIKH91XCd2S7LKkqdLOlLuT+uMi10O96WyEg0BdbnORwZzwju20z/J1vtxf
WU8j30yDrACM9w0/WMSUI/JvCdDfRRfbFifRL9S2XOtj4URWmHDWAc67zXDMzPzF
wbWIB+qqCMI5UwONbTNP0Sx8/IV4DS7ygeqhiaHIpHsp+MMNno2c+Gg1UE7pnOvw
I6Pqmygy9ezl7Fur0X4OpknwYnysVYEjpAX08O/uvbyPnpK8+NNperPcrB21Nd+1
03eNSnr/v/kdkY41Nl3WOgeQZxDN7Bp1e2CB1Yus9FAPhVtWUD7wj5qgxs4sJEtJ
3Fn0fwwh0boir/o+NPNiGyRmu98RgT6zgG3ktITZI85LzPi81uGLIunrGQLDlBTm
pHNQgNOPfy9ngV/BqaVR7BYewto61PRy8nHjVYkYM9oDEp9NdAMd0ZF+yksjvshf
7f8sS6gOjVvBoLZ9pM2sLivsms6WzLAM+oKEyHFTLOSy3DKGnhNcmqSU1PLBKrgG
ONiNRK/OOPr2BrthhZl10pppAxzH7PrXOZNK10s0bbgK4KDMZr43vnPaxfRX1RtH
tdwuMK+tT57YpW6kmP6HvOv5UrMY6kky0H+EEUs6te7B8dkuhD3YFlkJhFichv+5
hCu6IgF0DxXVGSCtFbYlzYlRPF1HLQxAmkTW89fmQwMywmoBEsGOmkzw5N7Ot5bR
tyquT3e7qQOoeSDq+9jQBKE0qJamHlCiM6FPVrvjMrVAqt22IkOibHkYg0Bn6mDI
vbwUApd82dhK9n4dLSwsMEaUTj8tSSVWnzqBdw8M07q5SSW7T1mrJKHHgwZunMia
/oNjR2kyOUWeN9P1Ebz8rNhoADe6tjkeKPzzAnKoezTC7x9yHFTfabJ44qTyRvaw
0txKLKhVuidjdqFIQmL0Dc33u1eKBvmRYWGh3Z+b05ONFLu2E91zcDRaZIg7+2c3
QoffXPXl2tfamrERA0LAAejaswaiZZb7dkwBJ0jCrMd521cnTgGVAu7aFt6dHdqZ
SkSSeUC3b7HYY5f6LiL7SNN0zHlHi25DTc7MGqyPvKymJ4G67333CWzyvXhZaNYo
l2foyfSw1jLHFaW8DC2zzQXUJJX2bLOy+q+B8uBQpvgjYOEykc3UfPlxIRISngXT
3fjXT9G22QToGeJQli5zaO64o5RTriANCBhD3eVIddYShowcOOjI0++URY2RC2dh
M6ef3RPom8pOLaikjvSgkBAQj8xvG8ug+ysxa/QAbsuu02xL50pb1GbfI+fXfLaU
p71Nl9PPavPEUHs5upfuu8lb/jUfP+29CKMzJQiFScP9foAlpPDBZEd78z3RtSjW
DY1sKKmYVwgdHDfpai/MQjse6T+7RuPbtswoOvJNizJQY2CEd1RMfPPDxkUbhXkB
ow+LYkxNfRS5A++oWyaaliqNobmgv7gKDQkGG3njuCVk8pH1TPb39boQoIAfnw/6
JeqST7tEWjHu9Y3WAiPzEBFrSkIjcIwPviXBg7LaRDrLZ9WXhfheyg/dYTWr/QaV
AONOA2lsOUu1M+HWz5TlV1YB21PN6lhnEu/+9fISCqmEQZAZCrPCiA9sSxPf8XsE
hnLMAv7UtuXWw8ZQXiegvqsordIGqS7W9Ks+xUfiKo62pHsLyqfShwCaMnv/iHi5
9ZrsUwWteFK9aUf3HMQ+oK1Z9GFNuNL2oOCWOxPEPUf9ObayZLIDpCYv/LCxIFf2
fYhhrerVS/UBI4ars5Vi/kAirRwAtLQJyLuZrFrxdIqwjwFBz3AcIRkfgVKU2XFQ
ZnGlg2pO9Y9Evd1QpDSye3klMYlchFbEGIV1ZbxNyNa9muUJ1/vVe8qOgvG2iArh
k41VgfeUZ00AvujgtXlG9kfhATURQzD7qWbDvmrjAZmSLI9NVKXg4wcC94oAQT31
J/0EL2wcNZmJJ8OC3BQlopKvZgyeFIv0IKkDVFBLYP+00nejSQsG5+HEDCFuyHJC
wO4w0MQgm/PSr/gNeLdBX08TNYbrFnXt+f9GRHHKKDhgwSr5t7be+k0GRqjDaYfA
Rgbx2khkTmKrzBpxk52Q28xiT66Jj4/CpDVqAWVI/e8/6F0oVFaud/vyaAAM/iS0
WUby39QkkqaO0YKJf/VfU6xtCWivdRurQoymGL5ntZNIF0QEmUKKEt9xotcflJA5
6Dq4sasOAryfEQBq1lUW6VqmpPA9K4HC1anQ3mSuAwp0B2YiHB9z+s8eCExj1PWM
hmWz1P3bWq/VsZPS4vvwuQLsowk87kiK8ES8TD92ZGJeBKRd+yp1CC9IHxqTTz1S
6AXUOOEa5emr6FvU5J7FCNQf0vNDJJvT8BlY6BVnE/dxNhhMg9ha18Wluz5Q75L6
xN5LfinPcM6fOUFxMMbxhFiLAo3foKpLbUll0rRpT3DWE3KTxW/pI6Gn45mXPyO0
1LXfIg3B5Qnb0raq2IOCP41rh1pc32V6ZGnhEHo3GvI1AJViE5O3VmF+bM+s4jsw
YqJQSoPFw9IiY8GcyXQadTB64qx68UwVFjaBuEAdRJQO/oxF4hQaKrGqfb0xqK6Q
X/ntErYEXKKE34KQY1dPs8+42nJ14w/C/34LY5fiW+WwvYEsl20T8sFJw1O/HC/R
HoH5MhKeZ2mbT4Jx9sNv9zletc3EFkSSV0OML4W+4xkOzG3lDHpJizOLSRA0+cHQ
Ats+/qSS2W79m/5ukr+2E27pNRe+GO7io+uboc7zxbBF9HfGaSqYGz19GF4f03m8
KL6KK3xF7c7cLvZNBfbILmY7GozoRxuyQqJnbNraXbCwIxnzXr0Mf/w/SG3EzYbu
u2feiKov10B7bmsCRAj3RqlO6ZoutN4oZP8ggDSjq0H3szSvPd27n5pLNgTBN239
1S4J2ZI8Mpz/fUgYLzqlSxMDHTmYS4sBsyjYiLYe9l2gGsKVxwomHIi72k6eia3y
Fv8wql/2dowhJBt9pAzBQpJIbhAC4ga+ejrGS+LgKnX/oAWiu6gyu5W2jwMCo+Id
9/Wz2uZyiQkZj2SiOxm9+zMKMh9/Nk24iTt3oxGU72e8508kJtQBkEHBibozoNjj
szpS9jpqXgXuonsYQlRTnClaeCFvVnrXW3B1PWSfRXktiNP6AZrj1CCZZBCl+zk3
MpPTFChhkYpqj3mIEbANKc9KmJnj/6iPzzve8mPBzgXQQoZU8cJ10qvegiPVcnPz
LILP8blRhyHVG9u3yBOK9r27Ew5Dgwg1myLgKAsc2KnZREYKHHCR/T7B+vUxszGh
DCbNRNNw9lNeyIuya+3dqo1YfVIz8+fVgNW1iWzn2Sk5xDD7IJCpb9IVG5eROqUc
qAfxATmY21fvaDGb/LlxDri5+koeIOUVschN6oLIeU7wHDihPO7caL2KqXHPtOhA
aVEDGhkt5Ae7wCso/BKKcbrYjgW5LJ2iokzmPRwDaR9+FfXuHFnuEm7bp26ayXJL
svOXXky+761X1Cb4hUs3/iF7oi7phrlKsyNY5JXOkmV/zf1lpWuxHZkMFuzJW2uY
PU0yK0vDbsrm+wl3IqbjOVdx5Ia6PXtkqBa03ET4jJYp5XKLTJvSWEt79drCZKhp
P0jgTe5NaBHVrvabNvq1BWwT6T+cz6pII5b59+y14HlO+HDPwApq8ZqTn1YK+Rfb
cyibOVVW4QkjZh3WwCHsb7lDgUlRz5TEiMiKzHZ1ut3inVkUi3kpr01LkBUVe8Q2
WGP8QrmjhwWXjCI3afjt5k4pytvcrSNDw/p7nb9GYzvYsp+bhI0D9/nhyctzzAAu
Hs/M3gRC32ixodncf6iF+czN9kqfr5yzPS6oWE9mNQQBmhgJB50+Cmy/DL7OF04G
CgcSPPkro/GGR2U+2q28+/XDYM8touv9rYdH5qeCydLCdG7eJRsImS3fwAnepkMe
+18TgYbAl9688AKLtBz1E7fEfj0T4vr5ORfjeb7Z4nXrDN9YnGuNl8inWxLIDrZa
wY7brOCLzCUhvjTWNNlqiV/3CIcxpi8Rc2ov8ldz9xdu5Aw0xlmcxC9ubaAYiIB/
FofD+y7YdWns1rgtjt0EDBfOhYY7OtVzeYEmsmUkk2AFLK4/y8leczJwcuirNN04
aJeZzdiOYlhSDz4nGDmwEQP9xfnZIikwwsa3zD+UV2SCfLFmVSXMJPwlGo5ZTC5A
Q+tz5yz10js3ZDWkaXvlfxEwrptArg02LDMXg0LIOXthJEhY7WFZcX1fyg3vGufU
OcR6vv1GALbQH4ce8fNA1ghc/wAf1MNGyEDgUWncfH/wdbirmyexcOZ4njwaSLXv
fHc4yKpVIX6y1+dDJO2qk7qrzOkra+0ViJ4GevMerLln9l1zt3Iddpzpu6SfrlAN
k9LdtRu1eG+tfQzIApwlcSxWM1A3U06Z0fqipRuimJlbDYK8wQR3wO+Yqe8hLEwC
+7eSDDExKlSpscpzacELT8MEeu3AGZE3LSO48e4QsdtA+yLrHTX31SiWqCSbOdew
mk173RqkYCfFCPUZ6h2tadIxKA5fJ69m9nE/eSwAopUoe7rSueCTaZL1WPYz9p88
rYSI8RxnYqM5Do9UMEWQAx2FIntzK60PI/d0hz1jm88lkVwVN5ya2p+UC+Rygc5r
4GxxEqgzm4dHhH1EkuRVPP10dPHyoSIFs2eiwzafsyHy5CBBs19IXfdcQuplQRJw
iUepijReL2ZIgiNaG1Pj62ShhB2l5QbQq28/v2iqtoeccYiAtLwIZA/7sakX+N32
r8nlyo8zallMkXrpHPSgzcfExQ67JtJcL7dPDx+kZUexc8T5/iltkCkM/o6YktEe
8yaFTRs7cwFCiD+KpIiD2ZVqDunEfLqp/WneGmA0y1CC5ti9WRC807EyGDoisV/T
4v8WVyB38mjCbC+AnVPp+73mxilazbNPo5RY/oG5JkE1D2XTRem6L6hP/R+IKfQo
bW94Cxj3sSmGII2SwNs4xNMiD9BaAZhJCsyNq7tzceJjen/lgYwv+nJ7h7QAjyuP
8piK7HLRW/bYDYlY1aaVET4k9JECPKmzLFcpyd1wpfq4HTAqxAqY2W829iQMp99h
Ou/8qlsheaQDN3onDoBS8JyOAd2U+mbQD+X9T+xexc6x0fdckepNkbFCaD99EJb3
YuOKHoKDEYDtb3gXXYP7ojiqcJ/FwNtjAoCqK5L+81ecg9/DzHrkdYH8oYWR6JRA
/Soi+7NNvlbTlMCIwfHRybm1Lz0cX+86JfFN0yM3v4xYqPK2+vNRE2Ev/Bcp6HzR
TviUcJHcCK8cM+ELhJUfwVYJQO0TP1r5d/2bCIrKZkxudKol7ExC+MSuvU4P2i3x
SUFO0HvbfYdIwPh1LzrFIGQSq4NvSIP+ItHtY/AazxMQ6aLDMYt4otmODeiXgTNa
WtYb/0FOGX/nGB4J+LzKmGxXbPEN5e9y/KcWSRyYV3dMyBfFtz+jWX8Djt51hkBF
zAXdKmJnHorUwkqNppzv/Or6d2FDeVBWPvVA0oi5cnpChcl8NZhDrGSlogrXMD3R
uTxVroUaD+G9J34SzCEUsQJHRoBxUY+wXekOJIXr5VFwbIxPJlb4P5vxztVyfaV0
qM5Hxl4fczmL+q5tMu+8BVA9QIXNdJEktaEBc0RK9hwm1WCfzMMSc2QMd1h4Rab0
Bg1xMaY/pTE1GE72DmAzhEdoVuomLkfxCw/dDaV6dWp1BEjID67p2aTJbvLq8iif
OLm5Qd/qdcgTjhAXplgnmD3S8+9SVVMQWpm7CV0LCEnL0UkJd0vAXga8zzgzBpIt
mjiMhfNcjCarrS2hLC/72LuAf+2jeWgXkNkYeAVwgZwVo6euEuofLGyt+nNLRB5M
ShcEinSnj8/+mrEbPrRI131IdEqRYkQOcjCI+i7UWqYRhobZZIBv/M9v1pZUyOcv
YB5QboVymA+BrF956yLM+uCaj6Qi9jLzji2uP9d1uHDLRjG368jM3Zo2+qncvdZH
NbP42mArVxDCPF/km/XJalZ7rEQOAeGdSxlNSpJMBbbJ/u3A4hWnIwX2kT3KraK2
u1hxYfRtVwMzl2gtUS7LjfUOcKvMoSNskBNK0Tizl12vBYBqt/K+VmSHsvCtpdIN
LCVeP2QzIfLS3GLdYmrnjV8lFc2dp8UoyI0MoBkGZ9S277/bmADOaNdkD6vKG5sp
krjI4E9NvYPMkMRIECUpCEiYv/ViK7jJkk2VdT3vuqZXiYaHpc8E7iB7HXF7/t+m
WZmnk0cuzNc3kCpF1VkeCPzH0BD4KWamoXXXICBa3QxWlxei5JefijXvGoJzgO+G
nCkzqh+xEUXTYbxQDJ4r6XECdOCDStN9tZWkwDoF3sZkZRKB8EiZFrYiIGKFP7XI
VK/M1wezx9EDlwwpA2wv8z2DKbkobyTxwPd0YRj5fI90SrfVPDBjIZbK9korRhjh
k2cJw34txkROzH193cn7q/mRcB7lFXN9iLM2joWA/8F1Gb+m4yYKhiIvfvWhN9bm
MIQ6WbAp9lybnA4p8mtd60wxaMTXzNsL6e9Zqi5zz9TXdcdVlZTtwOtmwUYVC9ip
owv/Y8AEQoqDzT6gyT/rNfxvpx41s3NRk4CtLGN1tmcMV9WBMgCw6IETVgJcaAr5
gfZFhZRde9QtuD2FN2sHBiewBRWyGEdEJlMiEVRRvxvomyEGJnBwDZsLHA3+xfo+
MhMYO5SHe9leLtOL67FFf859FZp6wZO1C/8LYNZHu+PGSJQ493rpJVA+t4cagHZ6
S9NXmldefA2KMJeMPpK8BawePMnoLLegcf53t3TZt6+xopoSvju0fM8LG5e1X49N
fesLYluuqZJRC0J7Fu3DAFnx6BjgJ5zuQ8hYTIBb5lvReo0999syUE+Gf+pmRLM6
A/0Mhqck+OnzmLdfYRdrTU0k4c4zRwN7tdRoixSz16MSTRXVfsMspboTTJO7RMSm
67Oup0Lqa20+8suuZxY36Q==
`pragma protect end_protected
