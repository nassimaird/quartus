��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_I
y�����
��)�z���i���t�ky��Xzm�BG�+�+S�ص���%��\��\H�H����ԑZ	N�<��,hi���lr�2c����J����B-&>sD����jx{0<�l~�Eɖ��x;0�O���n Y���7�!4�Ʒ�(P��"0����h)�
&��߆R��@\����ͯ�ZF{֞Uk���?�R��+H[vx�8l���1�7!��Q�j�8���6��s��P�cU.�Z���5_��_]z'Mq%��,;-G��.��n&��"��kw�'F� �za�%&ƿ���/�(I��zº6v�H�)=.ڜG'7
�;C�Y����A��o��*��h�7W�,�wH���<4]�q��݋~�4�)��t���p����tZ\�r��f�|��ɨD��w^����y��b�7M���i׮�P<������V	���z+Z�E��+)����Ri�k�ң���'V) �K�oٝXwA�ffUu��4�|��+N�9����㐎v��c�{Ni}�S*��of��0��!��T�C����E7���U��ω���`�R�P`t"�P�5�WG�r��2�K��w�k�u��AL��]+E�ع�b�,�0bݏy�|�C仧D��"r����70f�o�K�L�8�)-��lӎ�h�n���ԳZ�EdO�Ĩ�7
��t*"5���S� ����-T���gI$�^f��[X5c�0��h�i�}��4����6.��s�M���@�X��N/'����[�
[�'��ֿ/��]�HUuX��ѯ6��w+��(�+��Ͳ�4��&n��-/ގx�����試��� LŬn�5<�����-B�A�.w,�j�Z��i���V��B��O��e�G�{L/L�n�7y� �y����!э?��m<���zJ�'��tJ0 j25/���cc٢Ϫ��_Dec;̍�����͝a�!�جݽ�X��l;?��ɹ��H��{z�o$᭷�����)Q�6J�)8�~��*�����RK:�02C�[�S�$}���v	iQ�㏀��k�{r�~�f���P0����Й�}�A��l�V���97��)���|y�1��T��"S����;C�_G�]�sޕ��8�A�"���β!_������Z&�kOl�����cտ��v�~N�Q~��A��l[�Vjw�2u�g�vk5L�S���u|��B�� |&>Q$�,��C��&������R���#�H�	�?�M�/�T���_���ˌ�,�2<��5�N%��n��M<�u)�֛�`��0���'�u�h����
�����Gc�)s��s=�GT�wzD�w0R����'ڇY�h�w3E�FfX�$C/%�cH#[����l'���� K�d~gz����M1�XH3��E>>�jD-�d��>浈`:�Z�m�)��|�'L3���IW�H�����4��7�~/J1I�K�����j��U������e���#F��V�@]����e�RBT�G�"eU����.b���K%-sX8��ZV�a}M���`�Ζ��Q�q��JڄV�_ѵ8k��U!�WX[�K��!�D{yŒN�T�D��U�z)�D:�����s>�/����[z�>��Չ�P��T��$}~��g`��x���U��*�Dͺ��}+z�J:9�/�H��1�*��5�x����a��S\AF�S�j<g�r��8��``��N�4"s���Xc��t�c�<�7`��������/��������|?��`�x�L���l�ٴv��I�p��$�d]��[L/�@<r�l8bP��l9�ny�v,y�JtJ�|T�0��1���p�$�TP�0
ا�m��BxȨ���F~-I�
$ע�2��� �Q:0���b-�a2c�f�7E�`���c�HhC�q�d�n���Nez<nc,��T6l��c��	�_ U�i��i!�jv&'I]�)Wq�A�A�He=��-�	��m���,��IM\8E�cZ��+�!�CV$Gˡ�>6
k{�+t��	���_f��a$��* +h��O���H��MJ>#�s�L����2T�(��~���\���H%���憙�\�;̓h�S� �H`�#���YvZ(+��r���+l����1���js���=�C��u��tY�*���w\9�T�k��^��94�a8���^d�-h�.�&P��K��X͞�� ��rɀpF���2�b6����Ȍ�*�S��EqK���O�NV����E�^Z�Α}���ٌ.���B��poI�����d·Ⱦ�[S�Ϊ����|�P0��(�qU�Mg���h$K����(n�hP�Tؐ�O�۷+��N��M�x}0�����V�r�-��⚧c_�h���E�h�w\)�B��	#�w�n����Ո�/P@9�AwB$e˅�l�`�D�&Q	QG�.|�t
�M�
�8��z\��cI�eS�� -UVDc���L��i#����}?�������� �Dj�5d4E`�t���,'c�o���2�h�f��7�h �)�����3��	�C���R�u�K��'�~����e�&K"L��%4嚫`@��y�����6��/T�8a��?RrUHnG�������H���Z{~E S�_�7��C�����R��=
5Z��v�W�������M4ܩ	Il�N&���1�-���,��d��ʶ�Hhpo�.��yˬ��@2����=.��y�u�b���I��\!��Q����]�(�Տ�x����� #��֊�P�23^��?]4���rn�zS�R1^�5��� =_Xj3��-2O�o���'���W�>|�L�E$�n���̺&��O�܀�4���"wi���j��g�����][{�<3r>��I�(J:m&R>|O"!
�ϓ	���w������M!s֍���[Ρo$x�tUx̡��q9�F��pO�Imf|�I0>=�en�5�@�V���]o:*�)�����Q��z�gׂP�Mib�s���R���
���{u���fB��k��<�O���Ӎ�����$\�y�h�t$�9�+�ݑ0�.����{����p{1"+�i!k��9���a��(_E_��B�E:�ҧD��=#ӭO�h@�����н%{؍�7x���G���A��6?�R�)�pЪ�.GM+�;�
�G^�OӠ>$d)�>�[���n��,:)!�챡��Bs�5Lx��a1�
���«��n��� @y���0�����S��H����2����fB'9�V�b��.�/��>-�"�U�{�8��o�zM����$J��H=��[pU�%q��,������_���+�Ǐ~ԛ�::|O�Be�k<�?��<�xp�_��Wc՗�#3V �T����.�rbK��>�/~��ʎۦ��E&�T�gy�ߔ<�yS��k�Z��8�������	&�ʦ�q]�m��f���ܖ���x��������'��@e8wFE�m%��k���/&�~d���j����g����"��v��۱x�_�.�z��C��J� ����;oU�R<�@�%�C��A1Ƽ]�@��է#�_�]T> oY���$؍�U�(ݝ��EkB�M��+�,�g�t�F|`�&y��V,J��Y�fl�X����J�b����Gh A����c���	�_IZu�s޹�,�lo�� _Ep��5B���%�Q@Wo�����@ܵR=�����Y�qG'�oz��F�jJ���~��9�� j�5�<��v�7G�V��m�k�b�x"������r2���u�7u9��m���H�b#z��D�S�-�6�� 0ayB<�i6H�c�
����hb�Y'C�oֵ���{��@.r�t���Eg���p�ʑ8c7�ރ�a�����f�(� G�D�84�7� <�N���Z\Z��D�]7&��C_�i�di�x��	�Vw��=�`�Y�F���Y�e���B�ɏ��hnR$�P`L�By�j5��ON���2VF��U;�6A	�\�nNs��R�WFI�е�)�z��>弱V�y��h�+����_��ݣ�F�?6TK��F�3u��J	HEt���6p�