��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�2�2�*��l��3�t��X�ڇF��j&�^��7d@pY2�H�!��a�k�Y��(�l�K;^S88�]��ʵ�т���;�lM�E�H���*2��}��� ��D�	qm�4%��tݷ`��������hz.����u���tH[qJ7��d�!6� �תM��;��܇�����*+//W
��v��<�z��vYݮ���p�Q|��l♙���E tҪ��ʌ)��oIP�}���~'\
I2/]fv�j����0�zi���&���d�-c;�xՕ7����F^��7��C��
kxk�,�b�Ӵ��)*k��9�=IV����K*6*sC�a��6��PXؽ�ϋ�7��p�F�/��ןR�,}�{��2	���@j�B��s�ыhĩFn��)�/���|��N7������Ω�o-d���6��Չ�B|�}naSĽ{lŎ}�P�g�����T"V��ԣ*88#�Ufj���!#Q5҇,��j�0�ZK�Pr
n,�"��+����s�GX����z�ӆ^��pϡ��8��цY�ۦ&��ȕw���D�=j�a>�@�����i��󯣔�7�AW��vˀb�-���͌�@����
 !|gu_e5+���y��;�KFIH�����r�BB`(P(��~'�(v�N���B[���u�����t�Oٱ���9�1�x���s�&g����
(�W�{���Jt���LN�7Q
��������}*H{2��@޻s��m��L��JA<2�Yz3��S�Q�@��]'S�=��,_'���_�EJ������jĺ����,&"�q5�'��&\p�b��IJN�ޒ;�˷!�jpg���5S}X 	�(j�^6^V[-+�0����֙�03��4m`m �����*� ���Q���4kI�autX���H!.��'�����Y��n�8G�ҭ���JHs!2z��3m/'lr��%&8�_�����Ǣ�t�O�Ǆ\P1�nd��?(':�1��6+g
�p[D3f�4n�-kk{W{^z-WP9Ut0c��3F����	�Ԭz-���qd��Ʀ[>����ד�u.%r�V&�\���Td��uEmie �h[S�!�5C�:��
�LBJ��.�p�e��pa��*��׊gWw�W¦���5M�R6��uӸ:]	��N*`J/1n�Z�BLǔі����P}[��sq*���^F ��|�F7G��U �"u����&�c��/��+%2��������2X1����$���]#�tD·�u�>h�Ly��j�� � �����ƏkDX�yf�t�3s.k;���P�o��`������)�,U�?��/��2�Ԥ��Q��0 �7���G�P^�󀳤X+��P�jxP���P�:�-ה��rl�BJ`+��ɋ�����n1M�*NXxی�t�:��x��������u��n�alv�T�`8�E�;Y�م�s�~ 2j����e�r�Ϯ�j����|Y8�Ӏ�a��Զ��=Uڏ6����߷�X�7cx��� gTNC�JްgIg$D��&�>4[n�ߘ�]^�ԦM�u�h�g����:r��4�JA�܇�0�]k�8��ݛ�/vDycS�Dl��M��O�l������r�PR+��rV��@���*	=8g�1XV�6����Ni������"��
�/��RCɟ݄�o���o�������寃����Hy/��N�������Ȁ�u�G�KU^�(������W( ���	R���
2E�% �I��]�kj@�3l2��������h�m���E`�O����zYGY�:ԧ���N>���_�Ë'�@�����s�B�ٙUKj�����v�3��V�FQ��Ҥr��f��&i��M�u�{���X�i�P�Z��/�q�.���&f�N�lpe߿]c�T���r�z��5��W�V�g�O���`4�Nz��`TBڒ]v|ވO9��:h�*��Q�\�u*�^��%mA�a�O�>zc���[�,I䲹����2���U8�Y�}x�RQ�'�/)�|ỄZ��李��uRɑŽy0<�����)~�>�қY���9 ��l�����W�6&G6�� 3���z���֌��_�c�{������D�Q(�C4r�+�3�3��o���/��-r�N2n�{n�����~��g߭�_K�ܾa|��K.��^����6�aX�ȢƨR":Q�j�S�6���9�q�$.�ɷ�O)Y#sd8���*w
M�u&��|���.txy���ѻ�A��B�=o-ڛ��@��d1c�8��w�N�q$4�{�7�M:�k�gB[L3�'� X���F���G2VM��E��X�/~'�,X_TFۜ��M��QH���	[�ui�E`� �+�;�;��\2%����2��WZ�lm!b�fo�7*y���:پR����*� @�y�� �tt`H����'I����bL�_�T4�D�^6ٖ�gq�~�;̀u��S���t!�#s,�Ǳ��4E���9�g����za���N!��+s���qů����K�k7a�iT��Yļ���� �E�]�vC!��p|��8�z�	�Q1QS`TS�Y�/Ʒ��^��=�.&�%5�lE!�2�$�0�7IxE�i���v0ϊ�I�CZT�3I�����H����R���&��[>׉Ɋ|r%�v��F
� 5A\ͧa�	.��$<�cʬ��5��޸홗�(�2ґu��P��
���-D�I����zm�E%��K�����%�6N��O-�>Qݽ&b�q�k���\���Sp�dUW�Z�چ��� >��ǅ�GD>ipz��]���*l����ډ깸T2�"��U�Ro䶄�PԳ~S�L�7�8����2y�v�K���\�3v]��h���I����Tⷀ~�tC`���w?az�ù�*�����^�b�g-Vq͇-�頺���;�k��0G�M�z0YԷ~JF���{���XV���Peoe����k���.�eQt�Hh�'b~�u�T�y��e��*���^�&2�7�	_�UFf��ǖy;=��j�ɕ"��P(�Zȇ���wh�D�da�1�E���O�D�!��m��V�7�F�$�ա��|(i\����M	ht&k(\��}l��Deu��)����+M
5G
���!�V&��T�Ţ,�f?Ȑ��k"&�X�D�<T��U�G+��T�����.=Q�m�&�؝��/Nn���}�?8�~B_�y���������on�F�ba����Nǯ�4I�7*4�6i��:,R�z���b����\�N�0eBP�S�ew��P�}omc�o8�[�V�������j�r凅d���� �:{y��� 9j�x����[��F�2�6��ב�	Jp%�}IS+
:R�c��0�Q�X3]B�늶V$�H�m�aw�H@&2I�L�����ib�4N�d� �����uI��G�/�sM�|�Z捑�����k PT@�u�֍Lq[�5�e®9P5%=�=�nN?��%)�A�N���*RT`K�Pv
��}i�]�Y��z�oA�,�>G��^� ֙��0�2�^�"-C�fR݆)}��3�0�sW�,�c�br�}����0��)�w�_u
�N�˟5����%��g���͞V��0��il�ʑh� ��b��ĐY,�c�ha��|��J��P����E`�ϫ+`#�qM[��F%_��N�`w�D�P�\\��_Y�g6�kg��e�^�*:(��e
{����O�@K]ǹ'X�Md}V�\Do{e��u�N=�*�,�6��TT9N`�����?���iI��k�꬞���u���I
���)�O0q�&��4�%��CG��Z.�T�rx-�v=���%�W�HOwec1�S2�Ne4�Y�ٳ�7�pb�����������U��˺y�t={��\;M5�vA����,�[̈�~|�`������&�|B&3�C�k��6���ѹ��$2<�U��e�ݶ��?A��l�׵��r�&m�G) ��1-�#��� ?���,�s�<�]��B�7J��m^��(�7�s^�.\U{-��4�XS��R2A�� �K��l��r@�����!;#������6�6�TO�:��|�9�*x�JgJ����#
���qk8����m��;M~z�ۚ���u�HI'�<YF���8����OA�����HET�|�|�9�K���F�B�b��c��$"��"Q��0]}��ǈ�҇ê�)"��K��>�`!ي|G�v��@�����M�RӅ@Ai;
FY����W��L����?��+Тh� ��f�Hm�}���A�)����"�y�숹{��-O�����35����u�Q���(Ԟn����@�-��%eB媮�#Ը@�C[�#q���G~º"���[py�����2�5E*���t:�˗���V��6��֬^�V��lF��(b�.�vo��
L�]��	��Ý0��_Ҕ�z�2��M	8z�T����V�z��]��B��h[[��"�Y��D�fȀQ�7�����Xo6G+z4d�[O��I1Y�Nar�P�>|16�����3�-����@���_k��usVSM3��*
^���Yf��?U��-(~^� �=�u�ő���!��o��9��n��Й ��8���u���L��jʫ/��xl�@�Q8����������ٛ��,z�ą
�B�z�'���!Sq��R�1�T�o
���<�2t��5F�'~o�|c�O��l� ��k'᭫#^��E��*仐L758U�o�J�6�}"���i�
���rz\�k<���::��p:�b����+�,&�_���Ԋ�^�|H������g\���-}/H.�̓@?CP[��5z�_s�+ゐ��Z���m�}�]l��%�-�gU���~�pOl�_�cܼ�wi���KQd��	����a����%UӲb� *z�!�w��9 <IS�^�����5!D��,��c�V���M]��^颺HY���Na���tO�z��x�����▧��g�`#���+��,򗵕�$���B���Ċ��n�N��=�Fha�l���)&~�P�vN�RFJ��2��V��z8�^6�|� v`�~I�q����q�����H�����+߭f�N~g�=-Y�h��<c�.:���+��o��/2��<z�� l-���AZ�����Vq��_�4W�'��^Ju�Ɯöu��z�GvMjp g��:�?���wE6�i�BR��h�%��b��y�^�|;��]��ɿk3ć��N���L�ݥ�}�� �ӗ�c�h%�B�O��U�:��a&uc�͟�'խL�ܼ �C�yO�(����K��v^�*c�̶��Q�t킎���Tگ(k�l�HiI0F e�^�����v���{v�	��F}KF�N���-8�m��;��!jg'��T�ӄ�n���uL�"�w�Cg���VJp0?��uN�#�]��Q�.�S\��2��+:�)���������>�*z�<�ql����+��?4��!�B�K�P�j�	Y��~ �m�@�Fl�AWh�r��G�;�'�`I=�q����"�ٕ ��q>N��d� ��e��?���Q�\BR*�C���������Д���r��3�GB/�����3�����$�m~Ho�7������=y��qa�����ƽT�}c����؊sl��0�ĸP'����3��ZoG�Y4�@����C��c�v�鱫Zo~y6�N�>Kn��� ��R}�a��6N�i�����u;M�a�F`*����x�c嗂��M7�v��c�#~���6�P�	�ϼ�ڗ��^��BѸ��h���P!����o|}���PR������A$��r��I���\�',N�$m�Ü��5DP��ؚ�Ο�n�����S�l�7��%�/��7p�������u�&��%�0dl����Цcx�mo�c`)�񙔧�V�q��䏹�Jf�>8}X �l,&��`f%C���6R*��a���ա���V��yBY˳��U���||��ل�3�bOY��C+��d�����g��Fy�=}�`���_�Zv�=��h��q:���������/�����$����Kȉ�4�������-_��ʆ�k�e%����WQmU�2��𢡼�
�t�ޤ'���eQ�Or�������Z5�z�ms=&;�B[�8��W^�m7�Cz�s��>�o�h�z��Z;n��p�K���>M��`'0��?�A�:#�^��? �����(���;���<���7���ë֜�mqn�r�o~B��\35�S �V�.���t����B�!�9.��:�s(!�41��K����B8	ec:�� ۛ@��܊is=���F�6�g�i�Kp)6���ܧ�XP�s��k��R�4c9-��C���R;�@��&�90�����S�J�?�I�Z�!���`~%`���ue�XHu�:e�$������m!	����|o�=������v���!�%3��L�W�%O�Y���^1"�{&��s��d����2�]O��>�h���2��n��
#+Q6�O�(�	����v�0�_=�(a*~���MVZx>�5z���ɅYo��D��&:t��C�������:捉��A����:0Or�ڤ�����ř̜�������nF	�w�W�%��=�I�`YE.T��r�"����p�9.�l�G*��H>�|��d��Ae�%�@d"���xV���
�VO�Tՠ��mm!Y��W��Z����R��|�>���.��"rz1^y�V�}hH$���j�:_C�TH(�K�꾮��g�&l�������c�ܼ�|җ�C������a�^�
�C���u�[���Z�;���[QH�O_'#E��<��G7jR��tZ�����7~��+�x�e�����y�
�������:pRK�����J怉�*D�g�SО2~��[����7��p�w�A�=6f�ZѬ��@�P1���A�8Sj��4��,��W���HG����`��01Y)+�췸nz~��w����I>��X�v9?����]0�2�L8��)�R�LM��[=	xҒ�XڥqV�����=)([D/jX~�X������Y�e��"d�T��8ʟ�Z��FX���し��A!���R���/���y��bGf39Yn�	Dj!`��K9QZIK����W��[�G߳/�'?`���2$��M�L�"#i�v��lT����m��js}���CS�F� Fo3�����ݹ"�yNi�'������՜�>؆� �OV����@I�$n��d����xcQ&j����0M]A1�>3\����Zn�z�V-0�A��������2d0�P���Z?��K�D`�K�q�@�w`��cے?�<�U��5ħ�ߘEÈ^�s�^�����$�cQ����DT����T;����W�ѫ�c�/G�.��͝T�Z!������c�Le�r�b6��1���*�q���I�:���T�}�h�g�2t�^�B>u0��\��Z������f�2n� ���25|m�뉤.&��=瀩��	-�v��; 7� ����b�|m6�$�+��0�s�Qe�e<\&�_�t�BY2�U)�f����	j��ާ���e�.�'7"��s�]�і~�:Ѕ#n��P9��أ�ɇ��S�c�2����4B*�T��u�lS���DD�?�ǘrG�ې����O�_��C�GZ�$�9��#|Ԑ��s
�zN��KՠE�T�����x���:�hodGd�P���1�/�Wl��B�r��&�P4{^���/��"� N��B�N�E���$\4�3.��1r�q�J'�.:�/����}G`�+x�� ��H�
8/�3YA�N���9t��*������k����g�%
X{L�S��X��6����W4Ll�ν�3[�5����H ����Ʃ��H	R��E�I߫�z,�' @�4S��4�1�2��ae7�AV>E�zx��M���\v��EY	�*���P}�m0��a����j?!2�!6���]��|x\u"�Y��ų��+*���@�q��m�`���X�\
�`�#���O*�y9asѢ�؁q[�����?���ﵘ7&I CC���>��g���g�֬F�M_�F��<��+�"����;������N�*��W�G�uM'FzB��bf���B�8��8���Qk[�6Mp�	9�MT�sC��%��j^�&�G���f�T(@������ρ�k���q���؂,b�h�a�fD�,��d��{!�uG��T���(�l��;����P$IJQ�q����.��V��(J��,��s� $�0s؇�Rj���	�{��E�����ч�H��K��6����;7pu,����bW��"Aئ��)���ϝT$���f�v�������.�r�J��JB�P���I�O��<̅�]0���:�^7S헿�����kXmC�JINw)ޮ�t�Ҿ��V3S�ڥ�3�F<D��M�1r�ق!ef���{uY���˨��9��H��;��<|�k��NZ@������3;Q鋣�5�ư-��I�8k|;H\s�$k�)�$���d����H����W��´��w�ݸ�O�y�H0�0�!S�I�="L�|���7���4Y����H?8q`��V��%��Z��Xc����O=2�*�%dJ�ݨ uS�>�zi,�"�� N��=��*݊���1L
h�٫`V�[=�<��0[��l�*���G�m��5�!T�-�=���w'P<����po�q��;#|��e[�'@�
�G�d��lkrR:�"�