��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG��_ �9FLC^��� ]��,�u�P۹��_=kB�8g�/�K)q0�0�T��rD���o�!m����-��
��'(��Y�ft��kƵwU�8�M6<B��3����mT�o|v���oO��>⽄����q�_h��P�T����$��u�&�� �_k3��\��;$�B��=�$�����	ƅ
 ���I� +�u���&�2+�k�k� bk��@d�_.�<�Jo�"��?b�H�I�u� ��F8@�ZvDSw����<�*k���̐,�xه���d�*��2��әt��%_�߃[��=~��^��}�ӣ .�L$����lcؙET����i�:�?u'O�v+D�V'��B:���X�K�i\��ޫ�iN��ѣ�oґ�%�V��+�uS|$xs��x�q�� Š;��X_�Vh-�͇@�y��l�_^�����ފOp2�I@��f��\��v�l��h�����7F�+���2��MP�8�n�oH��?L;ϧ��402�/k��}�M�d�Wƀ��3�FQQ4�?�a����]���h8xz�����]���`��f (�����^
��%I��t����s� ��yk��t���m�{3|4t���<D�
�� E��"�U�� �)�6yEA"6<'���dB���2�B�b�>�=��8���.�2	��lnI�D���[��yO�6G`��h��e��ɷ�2�z�4�F~	Iy%l`�Ӭ[�H��#�)L���A^Q~)_dܢ�-=�U�� v:�=��k���+XozG�sMz~~��̝�&�5y_�����y��z�ٖث_����H�<��s�EF����htp��f0q`��[u�#W4�b�A��m5��i¨j(Ymɟ�ȹ�B�$B���c�-y�KW�|JS܅s���;WS��6;b>{��
�H��#U�{:�ĝ+���㖯�rb[�D�B�ƕ��(A)����@�+���a�'H��m-%�%'��؄'<��<ʼ�yϻt�3��*��`�+��FaUpjshd�`�Uc>gC��A� �]�/򻵘/fJo�ո�G��m�D���nW���}0�e(�tK�o�T����?����������k��y���SQ���4b�ϛֿ@?�#p�Qb�wѻt��ep��ӜI}�Z��t#�^2OI�Mx�LB�8˰��\l��Y��,�:�`pe�<u`rH��xh��|qg�=:�p`՞��Y��"�iّ���sN�Sb�����B[��S��j ���]�LKōo,�wK��ck�e�aZ�_BJ������� �ɀ�w��S����	��ۣ��������{��f����+n>�7Z�O�T-�W?p��=KR�w��,<M�P�Û��K5
�ź���c��/�T��>�7�S6��>������-��z��ʋ&�"'�
��h��tC�`��ɸ\�譗�'o���dC�+O���?��u�Y������*�x�5���#��]g��caS�I��o@�y�J�40E䉒/Nk@l���`��4v�qt񱸤����ڌ<qj@������*RH�Z�+�E �=d ���m�O�}S�+�F/�;�\��)�'�G�	 ��D����*I��	0-.�,B��U�Rٍ�	vi	H��̀�L�7O�܀wlos<����T�o�<�
��㜨�Z���*��O�[f/\^/;z�H�<�ek���t��k�s$�e�teW�2K���=᣾�tJ����7xz��c�#�k��(� R���T����1ڻc*�������mj'Aկ��R� ]�>q�8,h�r�
Ţ��x{9��[޺>��c��Kl��W��_d32lZ�i���hz�����k��	�Ǝ�|�`>�Ү],)�;�+:�mo<R���`�s�Nq�c�j��}#F��H�A_�"1�y݇�cͤp]���tMnI�k��# �b�7͇%nv\��, 72���B��,K�R�z�O�!oE�-���V5g���+�ԑ�/,�����m����6��WML�``�Tj�r�g�Uf~��SI��y3��>u��Zm�f?�ٞ�/���20V��@�eP�p��Q�ѸY�'��%juV^bO)��d��S�|�u�
-Z�1�[�!'[H�?F����4�)���%�7����x_����f��:?�햻`L��@��M;�M�}~P��"UrV�J�l%������0M��O���@�n�(+���rS3O(B�I��{d�_v#8�!%ˁ:d,ܚ�cŹ����&h�d����)hQ��'�P�f�ϖ�J@P�ӓ��(�2e��U��%���L�Ow;���{��S:"S{��S�.���(og*�I��g�#����h��HO���Ou	���`ϯ�K$A0=x���42�$��=�IMc��ԩ}�܀!�4��ժ�U�q�qz��2da� ���y��A��ĥ���}��9�x��)��W��>h��%��?�GpJ�9�6Ç�3��G���X�tx�7�:=D�#��A�K�@#ˑ7�P�f7I�k��U7�lf�Wyr���Ի����<�ª�d3�@��vL���_�_�A�$��qy4DLH�%R��SZ�]A�'��x� �Q�S�id�=�n؜�,2����q1�9<����߿���ߌ.�d�)�����~.��8�\g6(k�q;\�-H|g��=�#l?�>�xaBܑj�As�>��h� �(;M�cZ�U����Z�6�f��FΗD�� �s3f��jؗg�q%K�-u*Y�80}E.�h<Dd��.�K6�\�a���pa����)�躱��j�ȰPm7������tSq5�^�֞T>ic��0 ��
�f�1�i��Λ6��l�x��ָ`��Z{>��^d ��)D�ɧIpS,��q7;��j��9�9����Ѥ��7%�Ҙԏ�^܄쥖�-�4���n�?��-pAQ	y��b6����iOx�
���&t�C4߀E"ʘp/'t����L�¿/3�C�g���^��P�1^r<PĄ&���`׏4��i/��ą6��T�|����˗.�L5}�	-�-|���ݺ�V
l�g �H�6�������j0ɨ>d�����!�^����kV�]oCu��2�r�p�B?8 �O8�ӻ0�$�O�7�FZwLw(�zح�4hJ 'W�]3'�iU�F�*H��D6�؇ �̤�!�yR�Vg�g=�?�~��K�=�<榠
J��j�J��p(V�<w�|��_N���vt�:.�Y&�[��hш�:2���a�ۓXr� �R�̊���$�/k���KPT�n��
0R^������Se�U�0ǌ� ����s �b�KN��ZGF-$y-��'qX٬�I��Ղ��,G%Ր����ɩ*��B}"��ꘓ�����G}>���܂�IQ茣9��$7愲�7j�W2S�񾘿l��/e�q�b�R���?�1|0s�� }�L������*Dk�y��)�RㄟU1�����@���ҵ��Be���$�L	ЛT�I�e8��ɞ=���q.V�rƍ]���ʧ������.��@�]��{�9�,�Z�g�g½ndl��j!�=)��iZ�2��=�/��M�7�/A�X�\�\���;�mp�ᾥ_J5�|�_
p�bgwFaNNƓ$x�ck�LM� �0����g= ���A ��a�%S4&�{�� `B��`ļ*���Yl��T�p�#^T4���V`�+��n�C��P�ͩ�%�`*�� QQG[���9\�C)���{R�4�%F\�_uQ��?�:�DAv���
Y���t=g�"����v�Ϡ��G������s)��+[�N4�ʫX��`�v�1v7m|�"�N�,��B]�����u���yo�/��0����W驏�'�gxȡl��ik@^N�g�Bm(�ܿ�k�K��ƀ�k�ŋ?��C�k�4���Ta]�bBk#���/��I~H�����Cn��y��1̝���M}ׁМ�����q�T|C��H�f�8��h=���8���܆%�l.�����(M��7�c����"(ڵ�������R��j�cPՉ��>QX��>W��҆���(��;�ѝQ��:����b}QHS�_�<�y�ӕ�A�	�~c��	^l��ry�#�-{`Y<��G����Ζ�O�����RT����Q�g�f����3T��Շ`\l8�l���O��(�@~���8����3g���y��w� #u0��%e��
1�X:��)Z_����|hz�p/��(�Eb!NI�sԶGT��q���^�̏���a6�B�_i�+遵t�/���D�J���ق�L�j��s8�d;��N��rDA\��V����O���d# Ati\� ������5�G��Jp�,a6ڍ~�֗cŢ.ȷ��媔�}EN�uAhg�6L��2�2Ύa_�	*Q>�~6�XqȨX�[a�Zh�3�c&§�Q�Oel�VੋuO`	X�ue��hF�����Դ<��hj��B�L�f���i����<B�Xք��X��R3�xA��d�B=(�v�ۦ e-��vԑ	Ddx}#��=G2;S�N�g����H��Y�~  �Y;���-9���4�v�K��]kµ��p��פ���c�#yصt:.M���{�J@6g�L{"ߣ�l����"����*.�9���!=��RE�lKP�U(�c'�Ж�^,�����m�%2�>��{�B&+��y_Ĩ�#�s|q`H�W|'@�,�3�v�-/H��jxpѯi��7��>D�8�@�̮Ec���(�ayW����UĪ��.=7���/�?��G��:�8�8����X-��iY]|r ��5�8�����
Qhڴ�O|B'�\�.�jYݸgg�=���l�#�a2l?������8�{nE��Y�Q�*�K*�A��7���D!7M�EwG\O�z����k��� ������]��,�g�h���y-g���c&Q��؈,�b�aףL0��}�Zi�_�W}a�z�9���փW�[#���C�2<�t鍄��>�|LB��݃x�j?N��8|⵹/4�TnR�}w�9
��>=�F]��-��K�E�iS��4�-'$q�G�y
:+��ؤ̳���}N��1�5��z_�;�����&ci��6L��8?T�6�n����E|x�A��)� ����r;�v���f��l�l��}7��-��V�sd �s�VR��$f�)xs_�H&�a�X=�W�\D.@����ܵ`v�s�s��g��1�e��C	��~��D�������/�Ģ�,�M)�v�Y���A���8
ۆ� 	Cc&D}W�yj�!�gx,�M�:�
hfE1n�`X㴬�](}5,���/��y#B��Z���6Ǿ�,H� <Ȳ��0 |B�3�*i�S�͚%��3��g)������ٓ���� ����}lE,}s�DRq�%��_~{R=l��R�/c��G�?\Ų�d�%�c�S���B�Ǵ1�g
�(r���8n0z${]�~��cm�ҶH�ԯ��O�(�����N�~9�˿��c��ї����s؂�>W'w�u��G��ƌ�/��ӶJ� &�sZ�7v���ȏ��'@'mO.�cj	6��'�9&.�,��D"�,�4���%+\E�i��ՖR �@�W��/�v��_� U$����-2e��t`������q8-�//ws�W�I�%d��ߵ5"!�ı�a��c�p��iB����bU�'�����"�񮫑j���V��5^�v�nUa��|"����2$�������v&9��B�l��l������x��a�5�9*{�mm-v	}��9�dިm�7&�d'���MMh%���+9�uy��T�GB^�����)��>�77��[���5ˡ���L�;u�n��A�0����S�0G��.��2jF]H{���C[�U�ޏ��=�����q*�F���p�UM1|�����$-a��Wp��^ a{�_@��_��