`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c5Oc3Zzv2HWBtYarAwLq797W6/rcZcL6z6WIiKir9xICWbOvB47Tbegu5DNhVaKC
Ol1CwB2D/ion0hd/LVT//0sKhYUDEykdMKMsDUfbkRhSQLknUV2LQtG9hEz9mZKu
kfTEbCLa9f6etkMbkFYsElVa1PRoZ36Kz77PfHZczjU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35344)
1bKVlpTMGULSVE4x3Q1OfqxBS6m6HuHBmxWsTbFwv5Y7aE7kSW7cJmKCKQbj3bqg
anXvVARMNpuZ71FRLTcrOXWp3pe6yNT9jEtqO+YbfskED2+DWQM3EoS/1MDMXaDN
EfSDqykIY5dQZMH4SgCM9zwtQx9hghR1lX3eiZjfMZlCZrK2TE41HbtAks5+lyqP
THrnDKd2tyyrLPDCMuTaAZQw966n5/H8nwvZJSoCo9gbXhZxHcnC9eblyVOuBBc/
GwexlOyXQxklvyzFKaGBpPSf18fq332cGELxG3IZECRPD2o97jMNQv25kSKNAJ2o
yDyJiEIajZgBTsIuIttTH5rMgbKWkNMH0gKqlkyW/Ho6YGbNIiiTKZzLt7LumiIB
pQy7jpyPt+uS7GNBqxJjPocPyzbAZ7TyuEl9y9t9AETSuEyMphjs+j20VvMxa9la
TgxDyNpfDy6cJ9FecY7tPZZwntA2GVAQi46BFQpXl8Gq0Kk0HlKdJA1MnY4yYJ8o
Ej7nppX48LHLlBrUW9F87XOk2HORmvZukQDI8Lwszown9vWDlx2HyB8TjYBxMecR
VbOp/4WyoNANK3Zc97dON3W9f9lqYALaBJz+4HtLKveHhnw4vcu3Y/otYe1SNRrk
p3ITn02GhhFJF56Jur5HMbtH1Zz56ZZI1E63nTE7ZGgWI/AHLxT85h2ElfMmaH5b
4qBiiwo5PgFzot7htwVl0B98syNzQU1nnZQSFlTXY3s5r2Zt/YRUQoIBNoCi4ji5
R2OnSRPRXrF3AD7+2kwr3QednFbAeO3svzrFiWJgSFoiN8YfGKC+F9lS/YL34wwf
BtUgShUJgqYP3tmkU23Sn3+s0476nLypKon/jLbu35kabAFJC+lUMXRC5d52C36P
VlZp//RC3RjCaBCiToiGxmg7wkBNamFRiGUoTcz9mEuFIsIqVxmqjO+5dGLKDHsc
SWmpaBsobiHH/MRgojPDJKGG3y8sl4u/Ve4EIBlxd8aoZYkqfR1sg4PRMcDwGmyU
d+ScyQqiqcVM47h02rQrPlFAYLZAkA98PMxBNfGKIbAwd+k07SaQ+gQ0M9jg4Ypf
jUX0jHXxTZ/hGSBKZ4Pmp3/RI0h2zwGFM2w1WKR+aQQQIt+lSVtWbPlt5rhSnabe
5Qy3l8CPsccZP8ZQ47Jd7lpUUmkJR4KtoKLrsCLBsWuJqNM0ojPw3dOpNqLVGyfo
GIwMUtuy6qmlAo6mZr/2dQvaZZESgP0I3Ij+J85ekJYLrRumctXbJkVNMYQSkqGS
OSKXOpuYjHDIiyuHqRhB50dPT5WJIMs6uaGkG6Zi8CB5L8gEhvi8WbqhoQk24+F5
opk9lf/fbVAvvkvlVpw9WIcARSoCByq6oaHhwHKP7Dv++BbgPyAqYazMnWlEFMvz
K9qBfu/mpDxNICRzolPjXTUzwqJRHgOpxNy4VOOqThW2S96wr0WM38IyY2z8VdMh
fM5LK9QTv6EkVERGsNakyWkC9Dq3xDnB8aWy54LuLobwyIkCISj2FG4/SDWHFBIs
ygVD24STxg9pSv33Emrtwtoea0WgxVpiGZURjo34qnBKoTxHDJktgQL+FxzgezJ3
VaRK0y9t8yWGly2QlmBFWJnrQGhIS4idrm353fRDehjpVDjg4KeBmYvsH6XqSM0F
WLsUi3iKymUdXnwvaNP2zwwtMqpLo9xqZzrXKthJUUnOjrUGjy95MgNIbd+SHQvs
TFY/RNBUolh8c6pGcVyG203mIxHCDMAL9jEFUoGoZYbsT/0E7LNKvdcRgN5id0BM
+8E2Bl1tPrry+7vqeNTAll0vIX3unjRyPhQRjkreYP8h2JxNy1HTZEelhrDobAeN
DXejQQMOrxSwM4vAQDyNvRLhGTojYVDT8tFVz+zuGIrczS4le/PdbIlySgAnFMBv
fiFv+8mh/2VXSyF5Ew5cajM2yF22GKTejDzgAlFMt63ktdNf1UtC5k4duDaIz6Z/
F0FHstI17OPe42GpEEqr8SQ11vCpySDCTC2f638RcLLuvV2XaGCh9hkz6F64rVf6
4+sFTdCuqV4JvqJkApyaL7c5sx4sy7GwLGcsv+oF61+mc+PpABL+LGeKeGEL3Uq8
MtQJ1XJCoTC+Ycs3Viehdqu4mKNLH3TumUGDJJ2Vpblnoek9MMCFKXuWAYMwFzOn
3b9kd1llyDGAZkABGi4+TCjPV35kIChcMwxBdcPdvkbZbyPBpOiym62+JZp/D1yt
hLtpZOP2pfAz3KLft2OtmhWs92Y50EMNspgz1UhMdaHPud/0VLNZVlrZfBDLnF2z
UEzqHsHyRsHJy4ts6fJTTd4tZEA9m5Tr5N6RTVKE5MHLr8B85n4oCba48LLHkhiI
WS1i9LDDJ1r9UbQo+XR8y1Np9zOh2HDyQouOP5HSfB2fXmYFqZiT1hLxltAdHo7r
f3khb+vabo57jebZ0lRP39p9UHcUI3uW/fwiy3enDI6wZwNpzA6ycVIS6lvMnABa
TWd5FAm6C3LLD7dNU22458tvJ18ADq79O2t6t1/82hG9gLkXPkO9aQhGXcElfX8L
lutbVGz5h9y/IjXde5/Oojsft7Kd5poFD/lZncMxVzuLEpehqfN5M/Gewx2RT+Dj
Ee2ndtRUloMBmQcnFEvXgt6DG+BaFPCR8FK9iChkm4a40fgqzoTMfazpk3itO0mg
rWCHQMFH5tgFpGJQZNLt37BCgS6VsCihzS5cSZ4/ubUt+/rcvFCrWPsTZEK7VCmN
zi3lQ28s0Lf++iaucwhAaTzeZm3KotvgianmQRPBFlpv+dDrX34lpB/F5jxowPT0
aoBZFgq/u4RA7qSuJznW+3H2ATNIAesXDT19nCy12o0PHZWWCrSl2GzHVB+usm0X
mOolAJubBT9D8G+tIqabZDwRZr7JFKyEIlhu36EmALB3O935sHgtoene1WNt9tYy
0FVmXt6Av9VziZDbtNUL7D8Cqo2zzMMtjHGaxzu6pq0VJjemUu3tyuAc1AbTNV8D
/I5cjlBpAXTMOy4ctLf2NRP/l1/ICDnKg8wZwux8lRt0Q3oEKdr2kzt2DvDZJXUa
LQ8YNu0WBag9ya8UFqqnbCa7vrrmhCyTWfCM/qmEt9tT+rh02kPfrofc4ZWgxWEX
ZhlbCwChTUx66gghm8umhBx6s8bPB0rVB85X/NTQ0oA1OpAME535yYVC7SmCmR3u
7Clp9te72ajWZhx7E7opK9PD1X+YSo0J6PbODzpNqweWIZgnu9+vsI+ThWfqVzPr
3nsLHxmYAR0DCbAvz5ReiSBF9S8Z3kdRUhzY7Qpw7831W74QlNVnE2aihoMHlMGx
i8Ut07mgfwInKUPoXttkWk6h1t/bI6TaRz9vyTWIbzsE668nIrMpJaVmZ0Y5NfMY
Hxq3b97Up4Crjkw9ssgLeZoEJStHHATmT3gpxbb5QSqjKIbPplI0ng7pmXf1H0xe
DT0rnqtFm+E7aTGtHv01kSPo4P8GbO6WJ3WDEpUeq3eI83ZBqIKw1iUHfEApEH05
zhOgzqFd2xD218T1k8t5zXg/lbVDMM9TJTptJLo/zEttQU+M6qydvThjtQri/oyV
H3j3rcuV8Ic6fa6sVyGIlvl4fcXc6gzJA5WtkYbkQahUWqBeRJUnp2dr/hElQ6kJ
r1dGiWw4/XHxPNN6pL7cjx62CldKjYJVJ4T9CuKvD6rGQz74vO18h+bcJkp6rLA+
BRhCa7Yb8ilJFtv6DPMmA6RP7Fp7AFBQmmHEiq0t9vfctDpMbngier4DQaw+rxxv
2sphsUIueOIy4BZSDREmg5RrtnDvA2UrSxT5WnWc8FAVF4Sw+YgQpe5iOw9hKZ5H
Fm595pBxLT/85cRZNexcZCxuDH8D8Te83q2RV1ZO6wiA6i07EbKobcE1IhUj0SSM
wqLidNBX4EJmVvsAzqaofWfbi6cP/WZ4pNEpdNUNUMZWHJFHuo4MEsg+8zTy82Ci
k9tJSOCE0YJ+PkYGD3F8EPvmBneKaPQWZQEXSQ1kOe5pBn+EjJrbFS7Qniq1u8Y5
mm/eAbfUsVfjI9U2yVx4OLAvrWkdoeR7OhDP6KJE/BCA0D/GkqNux5PR31dH9tnQ
nLRhCIBv4Iek2puOIjkBtNk6RbRkn7UXblBcMsoqAR5WZkEBfL0Cj3stynKMii6O
EqTGFS2f+7XZODvulgu3vgFRwEHEm+hHQDV03WSDjGjInISGldjs1/eCkLS37xtR
ygly0JAmJCcWuXSU8+xMLqXpv33AUktNKYt40FgxmFuNzkUnxssRsfq3aOD8LBu3
LJfW0bCluVEBMnLXwUIZxgHZswSC7e2P673CdYwVxxfWDYdjnIToJ62jloWA/21x
lBQRQ1xODo9VUbxwdI9styWSGDeb+WNVetD818erXgu23uXEEXYBrASY2nChVRt7
ixGnRgNny9LWnvVqKG4cJULWg8pbbD/uqU2ym5LN1jCCXCzalOoZfre4uB4YjeYy
yuRuk46+BsXHpVjwiKUO0HqsiO7gwEiqKYlIaOy4jpOFhJ934PfLCEJJHAWk3O+7
mXnIyl4d2VvwjVZvm3MSk84jzZNd0WsGib3Q+K0RV5IbCFeQUnpWNHh6wX3Ohaqq
ivVUk6RJpiDf+bFb0/Iz7Iaz9TdqUJCrTKnoCB1oOA7WsmqdvNmBXBYoQ//G8zkz
B9kHEjpKrbbUeo11qr9smFrsqKDaoGov9vx26IaqyZU5/L/So4joKbMovtoWnu5W
6pBNuiq7WQDtYIabRgmZohUPF24CJksnuFneVOjtiI3trjOAyPJDlfp63GJI63h2
iE08zaf6m+Npe6ltWWgetjo9F2NirOXOzjJ/wzLu6A/EqZmHJ+6wPFJxwM2L5GJ8
shAXnqKenMAhWstq/ED5vgusdgU/sSmRBf8tVKaLz5xT2cWvie2dutaLUPW0XRTM
ibL8hXauuTobQLf3iXYOcfuKZCbK2ZJkCvOf3BvzOiwbe/k7vQShuEskgYZM+NPA
wRQVybZkzCCU/r10Rrg1xC3SMRQ0WaJmQspGd+5nDg7WNVsj4kNxonU9jKbRp0kM
hQN/yOVZpG0MeJ/kgbki9UW+4z2RuVbarXiRZxRacZqq3wBrFOaDZq2QaO0I//vx
9zSV93yZmJmXI2UfpHOnNcQP+6XNZ4mxEnN+CepBYeA/N7Ni2CO0Ob/lCADJsNS8
qV+WomRjDJwgWJSbhNKx7QzU1RtFJgiDZkNAAmcp/adINK9G8ViEGLpvxsODPScq
09VRx9UXJ0vsnlSk/ClFJpu4OM7LoWUklBZpOq0KwnVE9Q8mp3K8WjuA7VA4Jnuq
2olvNyuLfPGfuLw3trBVXvYngB35ji0g2N56FpaVhZUPlYZRoWXQydg7yII8P/Jw
7KjCGejVSU7u2BmxiARJJSEnNk/n7a3a4OBo1PgQ55s4wDjd4hjHme4gLFdzMsHU
Skmask+/iJSKla+QA0whE5CCabFz8d0RKGBQaYr4gwQ5m+bwxM9+2R/c4la+o2oI
6/lIUM++9UnMvlz928FpF8MPjhiiV6pXSUi6laZHqro6YMsQ40lCxWA8sNNUdOB6
J83eRv5UilrWqGiEwRGAhCdBbp1ECtZ+y8cBB/ZnN/h52gcvw6LT0S/U2kxMBXyx
AJ/ox80oS9HfqSomNl76Gn1i4Si5F+q2B6hjC3Fno9F+pDB+A4TlrvQyPN1EderI
Rn1+ISdXh4qSm1rnvMGbmKX3zW52AZmip9WtXhj4UM/vjEWGDanWNtgHAk6vUuYz
AGjRRM7duiBur+Dx2Or7kVEhdJXYtBlNyjHTfOSEkzhcovD9LZWC58DPK/Shvt2X
PCVQhwmbnZTVqsm3MuH57GyqYgyDthVDWfk0oW5YqbY0dGkKXkRUJ8ayDrPk+VjG
0waPw9ZQ9mQhNFrty4nMwFwzkQftyf8Wno+0eimiMQT6s+dC9t4IFMiOC7E/RQAJ
s55m9TIyT0dXlECbSwwtmhBJskllgXFGi8QJRhQEbIZtgMgnICJF+vhjXNH4L/UE
C/4UyaO0tRsPXHoRbEaTN40/8gyZOJS2RqcA/p4AxRn8c7v2g2jJEqd1auO1Gkbh
GHdYzfVQNNF9sErLdDzmVMB48Iz4uLhhBY0fGMY9G5IAt2WbNVNA2AkIZ9t200hO
FZC617ZpWDWzFMmQQBxIjTUn9ULOttvqgNXENaPpLVTzR/K/BWVXXDDa7rsxFKxH
dLgoy1yB4NipKdSVDc67BIspWjLY4LMd+o6e/I4cExypJs37v5RjbwEikXBjvwLS
lbfgyVYg4nmOlScSQrfJIGDPmXBRzV9rUI+XpHlUaS469fRNUZZUyDbmhGpsBz5/
7737WtLA2lrM4smhfHl35o7FwsqM9nHWHLQ2mPy+edS4zAifPOjRqEecEaoOTZnh
kjkeICPilqVY7V5BnYl9nCKSxNi2JzgRprp2Q8nLqbzUNrRggPj1dlb9mLUqT2MI
5bWImUHvs4D5O7M+RQ6ci/IOqEzALU7+KRhU8hyf5bpgSnvF2CP0Uf9aXJutxrDq
14l3SYpO6A1J6+/sjkDb8NLOx8y+ikdjqS4fqD2RX5Bkppmz8EhgQEGhEXQSB274
9n3qdA91O3WlPvNDXRiah9M7RLmEgMoBmows98SAOwsHGd186UVq3lrJYt8QntMh
DOPDpM30vxkenzDgecg2zPDLWMeDGlZVAQQIAdOToDKB+qGJOAjh9ODbA6BunJPt
grBGn8dUAB7k/65gOYL4FOsmpojtOnjUvnVcRRwDt0eT4mYQlB1bi2mNu33VsTiD
QadmlpbnnW/ezj94k2bSa+GT0EBXRlBnEUUXOcCaKeeUBN9D9YtTuxb8o6fJVo2n
pTnb6UB0KGOA6h3RO14k+QcOqyFLDvDQzUP37vBVw1J1cJOoIpg2UfKcBLTugSSt
P0cQyntQCwnSltd3isuzUAleYJxHvLwjumejSTCy4POqs0RjOKP3728XBeipE5yM
yTN297vl6VpCwqZq9OjwPSKu9S8A/HkG+v28cqRDXKih4JELmC0131sJ7U1OtfQn
N9X74bzh+OrZjnVnRxNi/ihIrUeWpDPVN74uwS+ZXYwkrpQjRRzMD+g4zxpEsAWJ
nlb1xR2VoRwFUqwyBmb/l8s8J0s4HvgrRYigtm16uRmt2+oZTtMzJqfVIm4Uijl0
CL080Sk7rR8ZdbnrUtzKSpAy0jnQ6SuMrTkgXBlCjqGeuMa+jiT+ZKEtmqHS6Wat
NpYi+23LNglGhMj5J4CjJctbK7GmVieE/9X4i/UCvtOpFXQrcXtS184v3H3HFSbh
gCmHstDH1+ww2FkTPGco0UPJ6wcdiiFaEAwB815SRcPA0Yhk7ba87pscx8FgJhI3
AY2DMd4XuJ4Xr7do22U+8JOBzsG1uRYJE6CfOF/c3jvsAVrqHeeZztK91Dku6Gw8
rzzuaD5KdMxVNQVI3n1zRQcOEvBxZ7uiYgiBg7ZClW7+YljoQ6+/r0JhrTpbN3To
ApYW8ZjHGHMnO6uMwWtePElPKqXqIQI+XDr/V0wKnfKMtZFwMhXSDEA/rTfhQiwZ
7wSue6un4HIbL88vWtV6NdKgcCfaVsCv66Ih5M7K4lN/6AR8Qy61S4816HtPObwE
BYDlPtg4Zt9wxOIUmNnbtZ7dFe52fTnzLnUUR5Dxwr0qTvatT7oQhKbIEtZaHAAa
4FhNy8z9DQl6GhHsde3nLB4cZz5AXs2Kx4NZHPG73eH6HQdVknmk38m8GcDBqh3/
NGC+mBXZOjW7U7p0uuCzUEPDj4MdA10RqeSG7bDTkLJepTLM7r39SQR3COXm8Nq1
UmOBXX3mhZL1ZuisID5BrKjYslNbekFyPY84VweCQT3JHPsB8OSwP9I2RJNGU3qX
jR3kqeXvIpH/DGd2r2NweqeaQuW488KJCIlA0+r6LF/q1fqFdZ99NseqVnmiHDLF
JPo5CQUjxgPi+p9bVZ4vdLJ/OTuyEqMDBFibVs9XF9xMBv9YOt0hxnjsmi+czTpI
w9ArSn04mXkqSgZV8snRne19MZG3tm2NWlVHlQYR2e+EkjA0zIA0qZO1yJUHUUid
j4Ce7PQhtUpCw7NAlgEbtBh8hUyAxYuITbXSwyI8dFoQJ6u5OU5znv0926gd+4g3
Ju+p+eXTrWUDekhchGnZ8M70iHC4b/VjvJZ/JjXxcNaDeairTvde5dR+CNHW0KAM
uo06wnklLFG9pILFPyPk7+iDvYdhlHTLjHV2EeEwi5105+kdl2cZ9bAjWH8DecB3
x45mQMWzMTsdQEkb/6uy0JwNnmpp4iwq9TK0O/rZbsRvZZFMRnVDHaIg/ZI6QLa7
4BAawbdsSgMbWBbL+xX/6dwjecpoE5ZqfdqGSRNKJb/8nkktcSAft+1eG+QtMudU
jCUDtLY1E8gOif5paZNFsICjhCTKfpi4Uo8+6DZBtlI/LSebrnj7tNo1CLtw27iI
Q9u+js7rdJyBJ/igVm+pp2hblriVSRQM97R4T/6RQZLuXQdKvSvdJLnW3P9yKjZO
k+A8Cql2ZD/Fm7fnLibSdjgUvrBoVk1phW4tI02+niPp+A7cRYCy2Foe+kO5K4rM
P8ZMi6rO8j2wurcmOwzGWBQmRyhSXZTaM01LHDiSWXXBCLvvvQW/RkMLyUSP1law
jLI+G+sT+Mg0YRC7AxRPvydwH5trjYkTOO7VXfURwggVIfxlzWKE/mJ+NyfhiIDo
7Cv8mbhVKGgZa/qsAKJQfMrHQb8JR5BLiuhy6qfD4P3/vPaIufWYTPsf0bFjHaom
woALjejtE3L12TOC3gdgNZp6FO8xeqVFPWofFizafUwinxjO/btgg1jCEtBp/DTu
3hEERjk25ZTFYqt5ABG9FG/CgF04Os4eCj0HkpQgfJd0gJ1aQ3nseZHQZr1qozhe
gmoaa0waB20dQKCRN5YIVcEpiTqF4x2anynlqm8mPBcuV8UUKMOGnQ0mX/dkUhfo
jPsAZrq4w7qUZyyMVLWPdR/8VRGqtD9y7v5KnDENV/ga87H4p97bR0vlNyEVEZHO
NrtHR8WrjUzSd1gygQL8skRb0FEYVl5FAVtcvfIgFI86O77DSFSRm7kbVPAMEbsD
nUi9tMtTbl+o/Rk7v318COA4xBQlh0wNZ2cJHR4d7spTMFdScUvHdHUuz0frLcKx
yTsD+n9ktphT8AQoVu2pkl2whUCzfl2AjsnaA+rM/xaYngUqDn9CI+py1UbIgFiC
AafnPdi/ZLLgflK97bNRqum7An/9peOa5z08ajVoNzaNjt8tQLZq4zv9t8VITW1d
ylC8TidgTRuEOucemxE08oT6f6dYU9MVYTS9vTkyf2aAvIdh7ct/V504QnhWSztq
L0M6E9qlBXhOjrOwRerQxI/3IuNbY/U3EJrImJFeILmPZrEuYpZabFS6XBcVIMcC
zHUSP525shrgfy+0IZ4A2i87YkdxGHTY7EGy/tLNpV0e0me+3Nnva9+XoenhgReg
hxDDZIl2v+mcL3z7JnV/iR9kKqwHcmYlRDkBOVG1Xb1friugn9IbWApqWfgLoiP+
RUaAzd8Oj5ZMETzpx6gfPZQ8N6CGtki5uHyQqfMGzK6W2Vmp8pIIvSQ9Uekv85IQ
t8Z/bhlWttzZuEl/m5+niHDUG4DlkNJGdOT8S76sZO81MIthfTm82/FW+XY2iH7H
0moR1VOssgxzjK0Q01bs65iTBEUrpXYgEKiEh92bymzo+WMTH0t0u2S4/1yDywPS
RyBTO86bge2a2OdS2rnM7YR60Hyx3o3myc2bUOjeoZYMw0yrwaAharq/C6t0FWt/
OKVnrMgmQDgYt5Iiwvv6/xIEXtPYCrOjANld8JHQeHkWv6T2fCs6X3mpUjrn9/QQ
BwlDHncvF1XfGKFXMi685IGtBwhJwFSoNkjMWFBMp33m/RRVfCZVFFJz0n17trEh
AZ9ZAEFSsGZfjLLp1aNTVm4dml/8/ot+6X5jRVH/1WwhbN2rkB8zBNbT8y4Y436x
9Rbf46hxrrdbhcKTD+seNOTnHM44RiQ74sC41ffkG0SFUWFkH87lVG44Rqn3Bymz
2xIH6FuToywQQa+4VvrAk5qYBe+UJzmxwyM5TKQciPkyn/Pbpl11f/AbZV23tgE9
4r2ZO2UKRwzjvdjg9xP+eX5aO9WiwTHKKmBY4A/b4Vef7nGybg75awo/CeBdhhz2
YVsyLiZbZUHQlk4pGeGDqCMdV8RlkE8ZzCp3KRtUNyxcZvnNA8vAaZr3zDhUD0X5
cPyYvzHYnBYn8Kq6eJHjdH7faoYTvuPnhVvtU+m5fL9ZYWftqHaEkwUYsDpnxZJn
+cuWlx4dfn82vgvbeO71stDHlCNXa1BnTxobHRp0Sz2uhfFJRKPSk+VNA3R8qLOk
roqOdmef40mdeWVwqA4W64EwcEUC1xRU1/44rB7s3SLof+CAfeeR1ywrSXwjAmPC
NxQXJqgNy3kh7tPmach/OJbmVhPvXbD1golf5XZMtlgFWg4S8vx8Rgkv4zXaCzJG
vOslMwlixmOtyLj1pF3EUrjMPEGqZnktMdSqjmEHj2PhKDOWTxWtLvwkHH/CVwvb
zAv8rVKoJ7e8wa4gRZ7Jmvucnqk1n9j//xgWMeRlwuBIlZlNfEmcvVKmjCqiK/nE
4GmhwbUMPYtphvcJ1gpLEdQwdqs8s1qba1gLjPB2TAD75lIlJpncbMg4ptj1kFIX
jODpumbCNOCKQpSRDb1dlPXCQ3HKRmNuRwZUTlqeQ3baZ+OojOsmRfhpgugnyor7
VjT9XmAn/aDwv1+LJSgFf+FBNjAlTuTZzzb6pZ3VyWDsTTQwxHqG5DtFPwS4dawq
XYUXaBpjcGGeCPWEjt+vp4r/i+BsNRjbzBhRIAu1IRTo2CF1YE6LPkgOzO81g4cX
KlwGlrj+IsY5Wu6NHr93FfTiHNkeJsAbRMsuSFn+bq1Rbp+sRhfHCJ1sQ5SkowvO
/T2awj0EtVux1ezTIdlQaodcGHdxrRFJWk7hbKY2carqtvHbpEHvM0WCng7Sbgbw
rAhqQhPVt07CVMbQOzuSPyw7t1Or2ZiiZSWATF1J5cX5rHQbaaCOs7MISKCku1Jz
WFIA48P2tfrz9fyGvvF3ddxx9mXU+CHhEgRP7LuUt8ujwADw1VhNZ80tO7ykAg7S
uwpGL7JmoWwbdB2DSxek7KmM8EgxKq7fqzZFdF7YKgo2d44Tyvky4EhWi68W/132
qKmzlgdDw8rXNgekP5Eo5cqWz8F1LJH+wz71wgnG+UW+WPbUccNoQu7+iRVf9Asa
nB9zCHEgFiwroKMnTXhYRHQME95i8izQ85hZgGUS9qiqwpq3oM5D/t6iPdJ3y8rw
N5vRL8JQylwHA84Ev62Ncg3wZ7eILS7q79UbpPYOi+NcjvtT2Zqvp9F1jkWidzSJ
ujwdAq6Ly9ckaDXFMF4cqFDACwMKCMPVF9jb+LZONBCYcYAD+tswNBxME0O4Ebz7
Mg0HlQ9Ko6ExKGfShw6VZ3bJ/iyP7smEs7E8lek/b0notRahaaPviKL8tcn0QVcE
FUCisv8okwH0wrvEFWjIRJYKVRBHltRhnNVL0m2SvUe4jnMUUC+sb8z7ljzrER/1
VhR/oEXv1grz2w5I5Oddh534W09OqxEC5LFIv7v7fXs3t9mCLk+BB4rCLgbZWFAD
xzH3EXnv4r2sOw8Qx9pVJjxnXvfPFjsnKW8Awn7TqbBF/0vmj+tuOFL+C/sH9ahW
oO4wMrK/VrfVQ2obsCGJ/b+e2SPDUi81sScb8E/WJknrHkg3bnTmGCPTwHU/Z/HJ
QeFXf/LC78U3egp7sP+4UsdFfjRknk+R2VAVURHnPGU4UzHMGX8f06+QHepVq7JD
vKs/Q0CgyppRNM+YNtgspKpTB/OCs5svzQ3hOVQQQHoUQQeETtFvAD/yEGgYlCaQ
veByp9rlpnryNFQ6c6YzFWWfAEiKf6jo6I+4AM6kLUaKM/vfzm5hcE8W6442q5ch
uQTZ9SvyuKqLW3fmzdYGDWkQ27SohNl5A/9x3QqM3IQ3/LrgBgInytpCVgD6PJhu
dItyCUGOFC6H6kLz9UkoiekqxAz5uE+LC3AfusyJ5lM/Xc4Ra2A+QXPIrVRCxRtj
p2VP9647HYDgzSrhroC/AmAS5FB7eAFGW6BRm3aM057ByuoJ612qDDzXdQ7kdGYV
pQ+uJRpjy20vx8v0h6EHST0BkHSaS34nzoCjVF4G9u5XN6SOtD8IWh49yjoTTu+u
AHbxANWQN1I4xA4KpP2qKcxZEPSIBpqKpNA5QBOHVTR6ooRTPsc//FXzdkPt9Cxl
Dfmrq4ATfZeoQoayxlSUhLAomrKIH9z92xFFx+g+bfz6+cOzw4PzoJIW7PI/Rpsg
v8DE30mDuUR1xLDkM5dcPhUNpwxJ2AW7P83LvSkf27Yq4sOZmXAMxVAtctjH8PA9
aVyBrbxyuHMedtzpgYh9HHU3M98A9aucV56uh8SsDcPkEKF/2FKRiPYTFqj2kl1m
zprNKV3ulleVevwMiGLYtz+DwzANrU0aXBm4brAu89e6s2q4OWRDVEnOoZxtlRME
sogQtXqIV7k6eZWtz6yW5gO5xxsUwvUCCb4UppnbC1KO0i75qb074JNM3eQfmRQb
RdnQxzy/DRBRPTHJOW9olcOYSqTF2bnK7VON3mL6vo3TNIyduHeRKJrqH6JmPHLi
+NtFZI7FwhExn3x7+NTxIvv/KiNWbnd31TsSQEzGqUqjbDb773V7DKnC28ZogSKz
GVhcfeRhO0c746r2py0tojXkA4HxtqnF02/k81H8Rzo65QMunDbtZxAwT+IBZSlY
yFFVmjHCNkwNtcU45lyr4tsPzFR9C78vU95BeQjorLrbyGB8Ep07c4oep8IqYMJh
7AnlgdqHUBMhDTe2td7kBPWu/Kk6Rm/DyU/Pv5KHcGxZNI5e07vLd1bnJcgBY9Fz
Ubahlwxei4/KxPctkcX6GfnxQd1qJNDNlI9QZC5A96slZbu+dWGklu4e1wJeRqoZ
0BW2GtWyi0mMzYLGhzXCbY7rFlTmEITXSN2lZn/RVzkHlDVK6dE1MXg9cQDPAV3G
6qDDKwKosvC5BfNuEPYRR/bqRKeUo2IS9rpnzZ66kHSEwjixX0kLAwRFzbSYFVqE
sudMnzjCJYUZCwXxKXXBL4jRnUMiYLDln2E2YjseOVONNuvIM6V5TzHadXms0y8Z
x96iVCF7RtxR/z0qfLZ1+Xn+rbvGyQTmdoqHjogp/MTN3y4c8jJ4peyajBjGoQoy
5pMVBjbFk2uw+RZMs/o2+jaLu/pBCzoKxMzAh8wWiE1zz96fM7rNGld7HgGR4ed+
/97BASe6VDLc5uFbbMSq2zqpS4Dfk9oK5/cY866nUjOcDiaMbPIwLllwaJ5Mo+ml
IHOu7ckfn8DdpNEfkG2Q3y8r45TBYkGqJINLdu8eiOrPMsYbNb1q8N0hhGrKrGua
+XG706KYjHfDAn1BR+MKklc5igcntdqgTKc7qNHapC1dLSjyIq4lHzbfoAbwu/A3
v++1NihMlvV2x8Ik2Fz85ZVDTEWRP8sOD/pyX+c78ouxldeABOGiKAo07BILjP4N
i2aetGwhLkMBvd2RPyTX/Qkv0DlXN1WTOXO/SXke5hUTjKW1EuWjrDUQyYn3Mhzz
acrqcMReD0SQ8wn6zjzPivdWas6rfFkTnehFLXbdMHcUfxaCFS4iVPcVxzK/pPPX
AF6x15jx6ZrpkFDSex09lW9H46kphBxFDE0hb5sf/nU8S4qdacWo+F25ZzAQAoJr
Oo7MGQuD0mOW4ZWTah3CkJi326ZMrjzK3kZuP6ScC6J3tUycWGDqYuXX/Ng6DoBq
Iafz1lTTlA0ootHgWs59IDSblQSFXCLL0ulhEMnvBwXPZ0buc0+0tksFfjoM5Zsw
eap6NcF8LMQCPhTQ0u1iQen3iviRya7nYvPyAlyxyGd+KBioXrF8VWXJvoFIxEKE
SaFwRffxO9HAePoO38f17/gVahj8woizCDvY/eUhXNs77ns5GLyM+QJjmHLlZkNL
4MLUE6hlRcRsl5lEJAPB+l7U3sjQUrzRfd4oS2sRT7b2F1cNJXyXjkRPBotR5EQn
/tB15c612nAozzZlmUTBcWK56TizRupr12rOyCboNdzJtBVG3CU71JAlB+hNKOLa
LB9agJICmUgFc/M1my/9has+pq3ZaftCVkeTA4QZuXwlSkIW+ZWd6ICz2hI5x/nV
dvygXPA5INZhYGogLur2YivmxUBW1nKh0NXm8P7t/kCFhSpzSK85gmBNK2weCP9E
llHB/ZG8RLwIZsPrRMnR+ELw/I9JkAt4zcN+2koWYorhSeiIsDukIKFDMjFbCvwB
8BNbdx1HO8a/egJ1Kkpk9jnKIJISa7x6cxMBmymfFRYILqfiAsIzmjX7WDOTfcxn
L9SUqFUfnv9mrlPEasx3yAFhLBZrbIjEykZaR4izMgXbx6qk9SGnOL627yudakPI
XRRUZ7vw57sZy4ju+hApYHX8Xfw/U+42/G0NKx+N3epp5hc32P66APfz8U2YHhrM
pCnBEMxDiPUCfNSVAT6/WLFwjzAG52oA4wfcEivEsVKRRmU9NOSc4aMehlFWKB1p
5sCJbmIrUqZ4FxR03naxoed7bVW19n1ndKZ6BNoDqp0ZpPCrBdA5rErNec9OIQIh
HYMTI2qSrEqYafE08E4l59tJXNHxbOgzl5AS/IEj3+ZIr/+/6einam7y18bXBVDc
mQMElnR2iwa3sq1QbUQ92tPjym60pqJHgYoG8HgTickN1Gd4AUCVyYQ+I98bi4Xk
EdOmaLV5NseZm5nx4Sdbg2xK1Ztg/fAmU4VuIrD8YusQf0LHF4ppr+Y7hWSdVt03
W3DqflXOEMycggfh88w9NX7oGr4wPSsp9sjjgHZ4Dx0cStk4YHYWsAPlIG+cRm0V
Ngn+aoIs2oHlWMXq5f7eEcRhYfzqeTZFyIfPJhljxpeE2N8t4i+xbuwFk3gRvAsU
PX0tqGcU7vwXhHUDwh24n50FSoi2xTB5ghK4ypApT93Wytos1oVCRMQZ4ezYEGdY
sytuT3g6dMvU2DmF7n19H0Eu7yC27cmef+TsHtCurFT6v2Efbx1TauGitr3xRTMl
luwdFyd23XIJKFPflQ6gKPKcSIZHtfuL2XpXOPllbVbheJyFPGgQ1D6gybufQ23Z
gFynbt+sbqjB37t3E1mZav7rcWD9mUxYpTiIylsWJbS+zQMOMGZMp7K1NxDeyyJ0
Z2OYS79NmCtd1A+mVng0uOuQDY5M38IVMmnSC0O+uBhajCLC7AnkGfub/XiTV7FY
K4JaVmIOGItKHjhtFcpZ0fbsZ6qaSeqsh9Slc1w43YtANW8iPYyYlKn6Inat63CZ
p2DoGAcDzkBjTVqtapFU/XCjdVsafG1BkNL1uKcWIG5fP4pGmOBrH08Jnd7Tvzx0
lFgSMbLps3589qVFGkNQZ49JJdmMNWXGUsrR/nb9BycpPsiMUQu5bRD7B5aKTv8Z
bc3yA9c07Kn6jCQxrb0CYmPHxJ1O3oZWGgAW2Baa2m/rYvS4JoV/hWezyfmEcAxX
DO2n7m7k23ChllEpILWbD1Sxyl3BVrcWrKODRAXDxMOTz+t/sf/Uk3lehaF9YjkQ
Uw7HJNHKXQfC3fT1BUE+DFnGuHhAvfeD5zgc0NVGO8gH7nXfrTFQ1gJJvlvh0scq
c6zTlEuAt8vLgC9atKJcItnNjWvt/rVYc6bA21vbQPhGrVhvGypvXIusDIL4OxiL
5OGxM1etu1ndTNgCFyFVTSJlHwis9IyFSrBlZZEif0vCNQPj4KGQxCrM+iFIKkWI
RgqcVTOwHPdBZcDFCMlPrHnHCAjmjEcS8tcVJmx5IrL2HdSfEFp4BD0MtqNpQXVg
iiU3pb9MHRXgr8xW9oXQkMVOJwQx00Eam3JTbwBnhe9CTTPJr19LTdFChmHzifOH
XAsP1b+dFeNzSIRknHyk99coRkeYql8DPZipUXeSGq6suwapthrCZDY3ekVSLjCl
4p4PwEY7ZWobv3FNrDfyO85C7ZpmF6CyYjgBIM82L8ita2tphb4Vsfm5j7HWdJ4f
vOkWxaEzlKNmAB8YN1p5y0IiHpmxE7IVfkZdT8bUYBijYpEZZmoN5E9izXtbU8vD
2+auLbVrcoAlv13mF2AHoe3t/xEygLtyv6/RCgxZw4vaAkyqb95VTBt010BpSDzr
Z8UOBsSuldxR6RRjEQD/dMbwzcZ7VXNlmBC42s4uKXXTG35V9K46/rVHrH06+TKb
8B1UTAJOzDZhjR2UZADk8FUw23/o8/+bIA7RO57FNH5uszaZ2PBYMcGUM9fvnwb1
F/ZHyj5SndFMcxel7nklTFhR7OaYZg0gUWVj4N3IsGis2vkcZc4dzNO/7Dl0ZeA4
nWsR/uJmnieROnUK0TXGX9A9yuHry/toA/ZFiYOa4E8I8fOS11aKux7Wp0+W7h+Q
GJrXbFF5Xto/CSzL8eyq3LRFL8eXJvMDq090GKIjvd61ywDdZssz8x65BGUaWP0x
PHVYoHUTxzuNILSlzy6g50LCa299YBNjAkSJyVjGasQwaDkzQqYV9kGlDW4Sg1MF
CHCEgvaANQ5bmOCYHsA9cOrII7/hzZ/GtceJs+tdCxPE2KWlpTn0gdibo8FDvYii
uRqGrNQ+bC87iTXHg/xbCbhl9XDxReAQZfNwFLgTVQmY+IIMZrb9aPtzixfWCxSh
810LPEfCyaK+ZEV3Dai+4gfHzRtJwH6ytqrj/7e8RDON3LkpNL77ZZ9RnBWAahaa
8buI2mG0KyJam21yqNdeNggyXN9kmzBxBa1x19+PjT9/6IAjpT3fx3nVMLwAqQix
yt9XZauKfUe1NOTiZzedkR2ERCe5LQgEpgJqNEve1disOA8VC9nBPoha+cPHU1Dv
ihgQEbbjVWeKP7zpCrcL1YpHK4YkhlWiBkbt1+WSVeWmG+w4jg4lTvOiJqYlKYcL
P8G9+giYr/ip+V8U9K9ZEzAaVDF/UZFaeKBkJSqty0jGLPDI+HEHVFXwfawJN1SN
tfaSfOxUX1flccdkrsWm91A9vHj2CJq7B7UTN6PYXJwvnDx6UwCbr5yxPYKl18Df
0rTLQjPyvRS0D0mKcRxZzuNi90SrUsx7drhe6HdVffIXwYF3hs9V7tc4j1SRUvjd
UzOsp6MR47uVWzEEGH29Aq3lWjAXqV4qTYglAZZOkIJq3y8/uU1DdxJ4C6zhvWee
ogfm13gb6W4PsQNVFtmfKtwA/u00CL0e5pn4IPFkvU2nHEawzB2cmTVTMIPDARrW
yozAzgvrNDONdFnWypiUDKA1TnhqNdw4p4hc0UIX9WYZ2H/j2orQ6Lu7wT7WAPdQ
+1j6vyxuepleE07ICYdWjPWKXLewuIGLFQJsftfPaqArn44N1AvWGTreL3BxkKrZ
jGW1R71t/vkkyFKU+NiuvmdncUr5mArejGwdQyfoOibjVbesyySoqG/KRBKricgA
J73z66cj8ILtKH9fDXgSJCW8tBVVvaujgsNWBrRq0Rka4z4pSV9sm4qQ4mGma7yD
Aik1kZCWOMHqS7sgaVM42DamrggfTmEKZggzrR1K/4Cab362/Pw6q0Q7jnZ+tZmp
0EIH6rsSAS5lQeB6cqE7cRNaXHP5w1aomloiiveFM9KQFzNzwILlORxr9Z6QcHDk
BVhfdWcwiGbO8eUU3yIHi7WLwMl1sEh6CVapun9sBVK5EtlKoi/Ln/nyvKEToB1W
aIXHzxEs49loszUo93a4TbW/MVjAFBt8beR0vqfOwcn7DpVA9rrqBxWeoMk4trfR
awMmMy3ctjFOLqF/gUpfxbBsrtznOCjl2jRcrvv0hnGLv7jb3cbJBGluRHlnAA5x
zkMT1zKwDdGFRYHk/SgRL8HEZirLlhvNvizVyF1JHi7j3Owsu0jSGHEmWb93HdTW
omlicf4j7BXNQnfNYtrs57qosHpitmWId/exByNL4VmMY7smdf6wvkHwD3HFHoHt
9rbeDAVeelJBg7ibBaR/8xjm6IcH0LqQ85TBeu26PCNeJd17Jg+Gzcs5OKhJcYCW
8MSIo68GpTKWf1rVC/9Y7i2cnUQn44PO++UmPCsS+NagrYk36Vy6D6zTEawiRqmq
B4V0CUJNADXHM6PWHPEkUjUSqAyDUntVhCMwwZtPEkOVhgUb817eo8zYFrpzOyZ1
6SJrQ8ZzIXwmRnGtbZGa6QN59n3LWttQenB/feE8hK3VqhK7YWTBOCvqn94yUcMB
DfFMy/r4/oBv7XGyGf5D55DteJnulppU0N3A+vGTYL3z2OIsQYXGT+G+5HoPerLV
ObkB85jklkp/6HPi/XgLtC2/qRFjdjawvjlhhxRqg0/Gkc8DlMTjQm8ANSA9utXI
IL10nbnFxBarDKMP8+D2kJa/QoVdXbo0eTNM4zRxFRn/5CajnENeIoDkv5CTDvAJ
Qw2vS1b10tuJZP/3LTYvlZLd7RWzIx/SvF7DNBflt3vzYI3dESCpy5RGePW360Hw
dGqFZmpRM0Fj2ZNFfVOBxovDYNtyXrYddVzz9C8DH7Xbm2zgTdNSFNvYyEbEpoxa
Qv1hOvk6oFvF/ckrLcwXHMxw+ISVbQxf5jP7nq+ZYhqKF0jhvyV3NAivn+6Df0ak
CiTk8e0OcVySaddPAYIXc2mm4WVO6982eRcpyuQwjOcijv+6zlooW//GocJUCeAr
SXFWegdk/3GGWWmvSzVrAROE1jhlDbe8oSeV+DdORmMOYa6nw0SHbEVnyfVNylcd
RVgzUaj8kieBEAwkdP4mKcEFeqG4/Qz7qHkOv/zYCC1sUOelNN6wlARLGv6cAN4g
buj/Y4Tg3im6f/rds3bq1r1GgQLF5ukonYyjeE0SvnlmDM2qhUMTuk4QU57+E4/5
G0iFlOvLdJKleSPOHi8dKA4nbQolmQaXD1xTacH6NW/ADAI5h7IC+YpVikq4IQlq
WnAimoy2x4/uxVo1BjfXNXv04eQbQ6B5hxLb3rQjAcfa3HPYOFkQ5pgKmAuDT7H+
3Y4ifvDNtTWTzHJJBvVFoB9lfEjQ9y0UcuRs32HoSn3pT/ZCwPxTZZvJ3NCKS7hw
cQlkK68s6ryWvjOSSyFUx+zMXNRo5h/oU9OFqz+uGzOTo2uWvskT9uwwUzN3hFhY
kJTYjpNEMzy3RADlh9LAWNPZnAArwh2340NHreGop2rMIAp/RG5RsdVtm1ip7wqQ
4WuRyUnXEE7kupJ1cDQA3vVBxa7B+Sfl4gF6ZPUUh9SR8idSX73PBIjLSggNhZy2
cMDAfwWDC5EGHSabmxSTDPkEiO7OH9FbYmysIoeAc896vLOMqOQqvxoquN9QAseS
8N42q1b7XJuvjE8Os18Rac+mXHO5TXemHrXP3obFrgEDUX0Od8C9pHgFtNj9VReN
XC8JcAjtxhZ0D1r1HYOJLTwy6UcwWMEQs/JYmTG7dAFfV4qmVlMaj2Sku8CX+htS
4b8omJIImcc2D2rkO5MSt3OjH4PUwYqXVNFjeLoOeBPKzGssItXH74d2eAXuevDI
4TsSJDH/ftUDSe8HZGitjzZCsNgXB0BydYPRybu5HHOYALSSadc8HwZHwqkNJXgQ
fxrckJOBAdfFgo0G+hFvBdQZglXeqMkWmmvtTU4PjmexDcQ79sN8DOnxqodOCIt3
BvcpAVmsSKXGxVmz8t7i8uvEgZMg2zF8sZsp0V5Eun4WEb4hJ0rO7a6KdjTJlTVM
6YtZPM5IAHR12KJd5m8/gm4gLYEYi2br4VNsQD3WtncNSK/qdgUbhBPwi8nVdZTk
y2fNxwSAylhX1Lm962l9DF+P0Wgo1OkPi6XYyz0y2aJES1xUXFZV5lqICMsV5Q9c
WeJ5FT3uj2uyjsQYeZuAZap/hT7zKm4jc8CM2DnY4sqA65F8Ru5S58mtVb54gpwB
9ApiGggslbcoJb24Ho2nm/dUzf7GYKSOBB11f3xX4gkCJ1FLHSXAHJrki3xeXMMm
oBUdQkJ+kYlhloApAlqlgppXsJK7sq7hLIC8XLLUjDSooqt/C3TYOAxA0ZbVkkr5
E094xLSR70ddbMUhQ2geP1kgCCQnFemzA20WaTKoUA9o13DanxA4p9+0lrnlBIvq
xh352g8RmqNbzin4vRn41LhWrUXhaVymM63Ckioll7t0d8K59rjEVnbwfAlwlVd7
Cq3z4bs4ILoBWjmIQaAXv5wT5VFKqqkAjxCx3AMHdTuz2YntfmBi6nOSSDDCrcWk
seu77hdSASronFKSQh1qWn+b770BhY+bHAkag8SsCHT1MdKdKl9qZvRl4joYTKjA
256xOZpaszjD18l6pcHgdBpGDq2x8uTcas72TROy5nM88XY2llKdptawNGJMeyHZ
4YoOWcaiZlsLRLY5wTAJJNZ+ybz13CDy+VAiM0F1Caqx2+9FZeQxoIhCpYOVdweP
GN4QcMvx8QPvncJe1MEPaYdAIZDK/IOAfdTJE35d8zD/oSfgmu3iT8NjP8pQ8NkQ
do4R/HMnICVRDGEv8x/q2D62K6kxkBPVmYA+f6pHM9Vi/dG+JfY57sRqnkxGKvtH
jTDLdfDRiwRxFLYJK4Nhlz8TTRSQpiXZ2whddP0JYA31F4Ce7OCgew/fd6mrGJpW
J3/iIY0UA0YQgdGPSZMNmtPSDG4veJKqd31wMrTDzehOtv+fw+jjD3Oap5pR/0UF
ly3lWlIOB7Som2fABSQ1RdDP7gOMN1lMdsZleIs8yTt1V8rV240iduRJKwlJlDDk
bvG3WVZS8yxQEZkzN35fh89zKXrTL0rMiR7JeZeDR4UNB4bL2NyMhbD7j+86dl2k
Nky4MoIdTp2p05Ag360ZyZOnXs4kd9EuE7hYiFPf4QtqtIvjXcGAhr4drItB8NHM
ZCK1G0wUQhdVxmtaUfYrkrEeMkWoaqu3o9NGp37/ak5gtsxrnU6AW63IZ76RYpc7
s896CFz40QQ0CgLu2NLyzit0KbUeQXuCSj3N92d7J69j2ezp7kxwRSLw0Q2DoAYF
OJ+F1gyMCqnuNNYJHX9JrWm6FnzG3Ls34OKOq72J6Lhd+JjDaWUnfAJUNPDAHO4G
hEuVCSqn6PAzZp05pS+G1xI7EykzTruh9cWpmoCf/H/p15jtEltakPsM9M3PJ39E
8ttn4esMX5WylP7VYUJy9+vTqIQWNRnfDghX7+GmSExzBBxG6qcHRTw762eyiprj
6uZvF+cBpvbzrpmlDA19Q2eFxyiEpOoSP37ocxm77+O6RCUlLb/pIqwmYD7cJR3u
YOYyI/A6wBwvGRMs0lBRUBLHt5nDqX9iih8dHHhUAGaVMwkXKFSxOzT8euQFc5qv
r5d9p/ldma87Dbg6usDx1PajZAbPwPaaDS0Eq80MqAaylV15BcqBx+93O4YBLSbu
B7BdWYbpm60Bbn+pviGAFDrbaP+IegYLJ7d0kULu5162VSOukuyU1nhQFbuOzDCf
bt5Fw/raBEWu4uDFtzei7nuXedSZAupjJ8qjRM9NumZGMfZqhaUFRwT/04GQ0vfE
rUpQi9+JqSdEU6GsOGShnWOzprWCvJ1k7cnB7kl7y8X7muzv8py5xFlS6jt6d4pv
Rp7W2ap48VYZxm0+LH5zHBSc1OM8cF+/H3MObM2npEvp6ypfe5qaYuCwBsgy5qGc
xyHMxTvEEL0ChYORBpuKy+7vOOh/ZhXrVXx5OyZlXpNWEMAiCd41szJQsTNcEKUs
0VDLZvrzE/zRDtL0yCIqms4c6bLNWg3X9TetTSBbaBlGoSJ3xJybHEgkF9340im5
VkGE09t8D8YrPE7nLUarxB/pC8rLtdKcUdklRzLHyeM39EhOHtfs8OWPAxGJ56UB
q3KYY1i4uCAxhEDNPR0fxzOgYI0VP8gHP/kbLtC+GZ3GRQns7/r7EVwLy8xR5E9m
l89XzvPxf5QiJwMCX0NorMqQNZ+x8C7+U61S7gZo5jrqcPWOoeK8h4uxH5H42q4v
OBodsg+bq44RWkpeczJXXsfprkPjpnQUabegEMmWRw/Pg7FiH9K3VYBzy+2EdAeb
VmR/1ZsI+Pj/VaLhYb9QbLk5TiY29gIGFAbL5kE76N/kigTFUjxXE+DT0ttZH7Bq
wBrq7WvhXPFopQfNRAx5K5SCefJIv8MkdnXLCGOL5qXiYGPc4fy2cjjKaPDf4l9l
0Z4g74BPGCRxTqdsCJd51/QLVOJvTpt60rcnCiPwv5JTZHs6u9KAQ1LwHYZqxnx1
iYvQKfUfZw/pIsmdmJ2s3sXiI8ABb5xbQpNkf0mBkB+tnALh5O3B+D5FxDTlwK+I
xP33/zUkAl8p+xNX4Gnp1oEv+p240rq2uPUTkyk6UYTG1dbH6RYSPup2pI1TS8TW
PYGcl3I5eBaf7ANIeYzVnwHZlFRCK+E+ZSFNNc7+QK/LIF+DO+N3L6nJUF+4fvog
8MQ73VX++vAK+zKQI99JCFRiZsG2dqN9Z5xanvVtg10j0AzsAi4QhecRAOww5AUe
d7fbWhZyK4K3pSZdMRtENH7Ne+k4XTj8Ql4ZwpHE9QZBrmO+VQbET40QoWS0iiu+
3PEY9vN+0kewGPeHWph+fC8Ld5FMskRT/i9AomGPUxEH63EQzPuaET5IdNGNqA+a
hmUah+leUfXBlvVpoV5gHu2GIJbLKTGZWhQkecPNkGKDD4zeAEC/6dMxpx8X/dE8
hDPixbDW7mHEBGE+fLN8QHh5+x1p0UIg5lTTiQ//iRW/u7yvfPnkip1VQn/EJSuP
8bnYQP8mvHjOXsy5RlLZtOX+cUaWv4qOfHb6uPmxyfG83sKvXKWcw6iIuJOJ/klt
wP643PJjA1VXa6mRPns27JfgWm6MmQ6FTiDQ3waF2mD4K6eSjwuaJTdIlhioN+vq
EEjkOo8xrPE427u3QqOmHHi8Yq15bY98/tBH05uDng/fDu7URbHoXNc/fzZ9eVmo
e3Y1bT2N/xHGOCfLhiyX9R5tTqomSh0+awRhSigY2xt9n9YPkLZ0UXJWCL1IwJgP
D7kkBZD3j8pmSEZ34CUfTNHm1OwrxSnSyEXPCN5Tcjlny+X5RBZiyuLfZSN7Hhg4
0+ZJDCUx176oqsWpoK0qKLevsa5fjAiAtjySXhconoT+qpH4zll/aXQYYUslgFP3
iWWF67aqI0po84RDgxEk9lcDkw5EB+tCt7cS7diwJuaDVljlnvvUz812KRSmaqzS
U0auV6j6JeNl6dIT3Q7MUqzlwFyqscUks53g6KKPwPEWIy4Gx4B3nnqXFfNY+l+e
7TrwEDMREqWWGVF3J/Nemk4JQLEzizVTFXCIjJXg1TZOVqugAHPpBxEmz8zp7e5f
074NTBiAoIeax/2qghZreOZJAB75r37U8EXrtZTHNuI4x650afrfOqsHXjOTXN6b
bD99XF9zwVD+bLHWs919gMLj/ZZoSgit7tRLxMlq0OAXDcEUV8nQQ8HwFSHRN4BA
QgzAj95LmBiaQsfEVPUTtMfxswE3297+5NjAmnhaI1UHH+YaBrdNT1xFJruqX5cW
IJc9Fvaxi06+fe0eY/TynFKZcUjLqOTYgBJ3rPicTrmc+V0dspDVsBkIFExyMgmv
lsdh6nQlRIzpdMZKV1Pb/5466u7PbY/hM/lOGp7DgOmMd48V3dgluuI2IwrESjNl
Pk0xmXayVlvEB7/GUUOHYd0cI6QdaeNrm/JwjWPsKBXOpc3v6J7FxomiEPXON+zp
Du4ZDX6Vw5XL5UHp/gh9B1gzeTohsyVivoVuCCoPmjUQRY1DbHYjCTHpuJXsv/Cx
wNjz0ELKT8TT+GT6nru0s+JNrxzLRe8YX+u11XpOHr/1rdR4W32CxShKMoh+iUwG
x2oesUUTD0Gwf23ZLXNL5DpNG+QR+ZVGBUpNUEbYGYyRBwNe/e7bC/i9b8Q302FJ
030OLZwjbekadFEHFE37po3t5MpymEA5cV9TMPckBPhfLJJtJvFOWRIrPrAzx5PO
4BWgNCTf/54FgvzE3XTgWNlpJALGFs0sM1bCggoezRWQgFP5C7Avb2KdduiCPIB+
ra6iL5EQozruv3ASYsYMsQRxq4jhs2nVynu8h5ABHpCK+JFTdFDpbSYXwpKYLddS
UJzU601FwnxW3Gx/DkAaF+dGcDxJir87ka5FXiKb1tXjfWrY58AO5r/xZ56X8qiM
t2HDzw6utHkBmT6gx50cfPf5MDk+LcZN2o4uEqNTLXcZbgc21pZdaxRQGGTOtEZy
uIBKzeY9cugFhQHHRAL/6G8+Nm6qQ3DfwSeF+fu1VtN6CDMOHCO9aBvs8r5S1eCV
NksNpyYz8jMkFKaWrz5EpaHlg3Uy2JntaLcMO88gSJl00d88wDQ/7mA/KhMaNEJ6
vIRpKz6II2fyqw5xd5433w25HC/Fh3WBLG8pA7ZBcrbzePrjiSqExbDQzJ+yIfdk
SQXDFeaasjP+mMnjS+CLNGt7S9B+6wD/8nSHtyDnenaXSFlRRYEDaH7jmKfXsiPL
Ixb2gJt2ExKUEjtZtjbotlscfMZ3KWdSKKQXNxUSgC6DnibYyXzqtXN8WW4eo6W8
JYQ0yfk8OynQXN3FkxOiUVJ2WPSrHigoAs7F1Nx94vR4wgdPUHrCyoZN/5Kcv2FI
zt3EI+aEhcsDcZtxePurO66Pir699L0+dzYvqSNyzCGxt6DuPBCJq+djQI6t4y1m
QeObQGr7+9GISjpsr+aS1+yF0ApfPYr3UVl8iqDfTOSjZvrpoH9YUMKgKd5LYj/d
NtFpAYcwwf/LCinU2YN4/dVnHyhnsIAIz4FSwuQd54+9/C36+n4kvK7ttNU/G5YR
sBic6XuHt7x90GzRJv1i14wkWToD1QExN1ojWmxvwYOPN85I8aFJVTn+0DF99tzW
8xzCJowZhSG0VkhbxKwOtJMO+odMyRjLJOSFugsLZHSa2wI/W52/0ePL2I1IznwB
rKghCak6sPpKFoPQj9u4VD0Q3fSzayeiH5yZOKssRB7G4UHjXIgH9e2UyD4qMdQL
F6SPlFhoD0u1FVieyAErXufbATFPTA9Fd19d4yww+0Yts213k81Zy0T5Dc/LM8CZ
329/YqDgCzYoNUSLb1hHacg8zmKElQuVGl2KFL48/iDWLg9MOFFYUoU1v+xQ5AWB
qD97s0fuNIo6aGf2x2Xghijj/z7ZE/L2fYRzTJa8Nnun4je2M/cj4khGwV0EadSX
KRGvHn7kHoQwU9AO/tl5DSXlclWKKcNcLRZRRYwfM8bNIotTxMMB+yy4n8Qg/6Kx
rWSSYus0Qm1Ie55H7wXVzKo9LKeLQjRNTguvkiWdVNPjjuCLQmrmCF+6nGtNIQyF
DvCcfuy+cyUGnrYmPz7TiqIRh+tORX2OymwxB5QKib6u22r7GulQoj/+O2YzFoV8
8HY+9NgbkknZfBLRUMV/QsmBOa8lM2tHP+J1ZZyPej690EihQm+FQvM108d/79v9
Pnff8t7Z8Hd532bBYZxuNATTayDnebnYibnHnb3tKxWmCl7NmRIijbh3fl/mdohX
tjKcy/3IsNL5ZF7b8ytlFAYnd+p/raTGgZfxnLHBVVRgMIMSGS+dlQS566nSnSKi
Ld7BRVJmMWvZMMi+UrXo453Ket8yN1u3E/euqWHbyrWk/0leJ82NRRPi/w+Nq5m/
wBxBrLIcCgP2Cac8szLZ3yjXFH08I5vRwOEoBoob4tg2Wwmaj5A3/wqAug/5piuC
K579SlU0th9LmdIytYxSo0bc6DVo+VYsYmXxeBgP2+ofLzDokNlLKILQ/8p7RmoS
tFTB/5tGlOriIMRovgTJQ1svB0JR7SBB9Lt+i4cOf1ErZLXukN2go3MicTUKY0iu
ZtSkvowGawNpmep5iEWiI3WzoMHUoVk7CN3wvwm3cqVTk/AhmEsqWXhLOTMMmgQj
YWqcmha8T6dH4KUPwGLdbjo4pPcpwsYr3+LkqHjNyXNiMfCvErd7gxvC9YfLQgwy
9GFaSiFqOCYUn3ndp4aMkPeTwf0SzZMmmsohm8g/xkoICvoP0Bl93weWr7645Z5V
B/0JOdZuwnE/MRxwOV/C9qGjnWY9AS8nL27w2h+7pog2K/DifqMrocTUCLkFga6e
HiPFfoNUZZzOExZtUfeoROPcEQ83doFZfjUWVYQX4JujDWpOgou74BemGhG80cti
mjeibIlwGIMVfVOVCupOtapThjSAdHIeBLelQzG6MBUioth3g09Yh4YH3NxtWGE2
uOtHz4PDGvQJbl6jrYeO7EmV7jikVDhuO0f0jCmYI5wG15/6NXVDIEMgBhHT59Ar
gAnimirOZjjqmG/SkGxd/Q56QZfjXV92rscP4X9E4+NwjE6F4HQv7GKsTS/0vhAW
yrUwLkKe3Jf5TRnuZRgSTHikugIhC88OAXlQNGYIu+hAhw+79BHnh0gPgMv+Kp2z
TqosR938iK4yk+QswoWmdtsS8YTjoRLgCXobrs7NVCTK0BDVcuF5NXDlqlfGidmK
NhJqveXOGANmiZcCjv4UdbqLeoJ1EEC633mlm3pFexSIAwQnPLYnhIP063XennUu
7HkJCOSwCSQCS5K6vr7fDpyaN7k3jf5HZ3AydnTmRTVZPJ7RszbCE20A+wte4uKx
TbQHf6mq0XspN/ccCzgpChrAOsykme+lj+ftVcO3aAhmbNIwDewpRajz/hezwW7X
bur/76yuUBLILELHwBuDrbXLIfe2KVN1j/3d6M2NTmwkc3q5+pk/rHz/i5JpCOP2
433ZYMC5Q/0kP/C/beOwWHuWj2RE6JJU3v9N9Wa5A6thqvtsoAg8KjlHUPfzyCdZ
G7bdTW7Hbd8GhBD5ZUvJq70u9WLxV9t9yGCE5bVMjKYgLqn4/mxpPny63GnuqFjD
sKjYZdbWD2WIuitsy7YxyciCYFyN/hmrgrpjtdf3KryWOkW0bN0uZ2ZJggPQt0LQ
fPuLfPvBpVENRmFm5e3PDpigNJt6osRUo0eovOucf727MhvA+rNfWSCN2RJeVHNI
LB6906b4c9cSwrkOxIkadvFk4cyx/vC0FzKblpSKts95EcPHzTFWUakeGHp7zhZb
Lx7h3G7RaKmK96MGM+PfsLDyTMzyLcol3zdNkXwWAc32WZVabRIzsogLmE7iBeSM
u4gRcYX3u28SqYU5HGZPFweItp20FB6D38NHcBrLNni8qrDMudA3x/7MW46Bgo41
909gqUsHjvqpp64GMMlVI4U4XGgLJjqt2u0dXGHs4MbSCGiWY9rP6gCRglvHr2xY
VGn25c2xYFhvEtF6ff6unykFfoUG0RbWA38+FsumIfQBj2Jdc8HY+mI5UtANYWSO
ZJBehSznGi7Upre65RJfHYF4U+lBa3159kcwMfFrNWFGuN9Eg30jjn/Vla7FqKYv
MmDe1dU1EiG47tW2LqKWIIIBK1deQNXMmFTkgYEQyTSepQDJTwZIrVwo83c6eofH
IbZsWTLAJa3Zd6TN/OqdEQLZE51a2jgfhXxpKUNdoTsCxOZpLESH5Dxo3p1g5XXz
3J7W+oOk2kTgu5tj/tg3iXZNJu4XCDTBA+Ic1JQgxDGsHz1PFhSk4YLxZ15KofoS
vst5Ln9Bl3KmVZbER7QeXNllLEk1G9yv5DNpJeBtUhz34ZPLo1bs3ljaL1Vxm9AF
Zd23P/FogzHcaWqz17UQt3kB9s6vu6hO2u4Qq691AE8qii4xUYAHHQojQGZllF9s
Z2uCbMJA6utKBK/r1N8U9bRpnPJjhhsK8Hry6rluHqiBdDEUpKq8E0B7bJVjlz9J
aeDffaoAFKpzkqGr8hbVQrxpF/YBgvmAF3fQDcxPRhR00MsmMxYD8jInGYYuDS+W
t73MLLpspyRL1mZNc/l+kGLaPE8xFHcAfgOdXr8PqAuOBgjPqWW8XRXmGM2Y8+F3
9pZJJAcA5QpJ+KfO5JV+5jrZmEp35uBSTiDZwWD/KToQglJHKnalzZerZI8UKILa
fnvd+kogn3l2cEjpd5hLtfW5bG+lRGPjcxuIa2NHvs936TOeLyTEcXR/qUdhcTS0
yrLTawtwmLM2Ky6UB0diWPm3+h4JmY8a/UD3C75o9941cm0SmickNQGFhNGHOg0K
ZrIIBowu0uUgyf+FR7s2SWIf8elNLayJQ7oeSH662p3eZvuh/sL34slNsemXckTk
t0tDYIrgQRHAcrQvWG7NiiwjkCrKiZ5B26XFBN1n9bZL51yFCjesQsJLlFIsV5GM
SJx8XSq5SNOQYl/GDPb/dATY9HOKAH2SkkNOMgt90n732L1VKVYJlRqaAGEFX1tM
jO44GZkAzvc3y8Q1ACpEhlk+zBvuvNQxkgV1qdyLnsVPuUDyANgj05V1Y7MnMy/j
X8TEngafBQRFtr0LRU17LpC2oRwDK/oLAEB6HEkvsFT15wTyL56A2X7uI8jJ+Qaj
D8PXeL40lYHyX53LtNOLoqPmyQcCI5EOydn99WpFNl1J9Q4PStm1xofxwHHeS7Im
xN7Z/sWLhxKBi9Gu+3UIDRlNE9RG+mu/U2Tf0bsT3jXvYk8/vC5PzMgpLTHQfKVA
FOLFC3KWmXB66t6U//UQGe6pZcFQJ9aB7C4TGvIcVGcPGxEKYMBiK7gRY0pPqoLu
E+CGopwA+vGpquLhBsqiNF8gzDqgt16zzx0BNSNdRLKZdQx3kCLvQwtxzwpJWpbh
IZsxT/xYcA2OrMDeQpZFOKbS6hKxCGzhmSsUCcGb2CIppK+gIT4LcDrIn0Z2zNJs
YpXVQO/NcMkmknYAnw2gXd08jvYLvq/3sfq7soofd0JGQdwAba+XuA2fSn6VR62h
xX3AtA9IxR5xUU6XcDoE5aV5LKl9YheJg7zBmFKH1GzvBmROC7FyVgfa2eec6qS+
+K9Fzy8tGsXxhvqUmzLdtbvtnqHuLVqaJltLhxeAWrNdi/L4/LpakfduVKPDS/tm
BOeKy7Jov8ZLiokoJvCwEy4ZTqRmh2ofrV16xKuut9rYSRcdiVs03kR32Lj7Dq6t
5nFtkfg5Nix8Pv22xF7o9iKkY1TCWYV56iMDvE4wYUZxLH4B7IijAA3jTzEjtr8N
6u1CsULti8yWZULJhlNTSIt9AaBfol7PX9t9rivnXfhrF2Zf6o/CgoZhkBtod8vO
x4u0zWIK0b1SStPOqfMZ4HHJLH196z2w7TmagUfFjLLvoCfJmXa9GLSdbLZSvgA5
fJkUOotEennua5BndE9O756XkesRf+6lBI9JFM74JnXMtePvYcfqTgqmTe0/V/T6
ROJVYRKXmvjX44SWSauhDEI1aT2AhOqAwzlH0358QS3ErsFrXYBwov6GflEQU8OA
KmhwdGiqHFL4T5bP1dIWurAQJkVHGwxZhVtLgaRvLlOh0ZWKyA9EgEJkn2Np4WkF
Y2msBQt0pLxAxqfJVz6CM9Uf2x+hSHis1EsoH9Ogswt5/K6Zue+v2FqHNTnZNAh2
enop7+QeMh6C0dI6b1pQNIF6Oczi1Nyabo0lid8tfJFvue7U4zjtivPZAw2VPBzM
ballAQ4NNBnBu4bbRfqkSFR05lJ5/4P7Xfu2XLEwGSubjkQK9mAnYaUSttrojAjC
s8wQuEvTonF2yfb7jzYMOTLiCD3x98O/1fbJHNKWmNFyd1vzE9A55fmBfonFXIcF
i3ufLdP47yL88TzmA4FKESwkjBGKAQRop1Oh0C6EBlMndTcQUGFEgIjih9pr/F3G
j0h9HZUcCZTbLrht3XijC2wBkR/c2r2C7mzHJ5W/c7HR6YaWU0vTgEVe73A4d5iF
IZ5fEMznIBfzJP2laMAvbs6gcZXrdzrq/QscPN7+6c78ZxFFKDuD8ug5/No69y31
Ve2WouvNhD1ZJtfh0An/h81lTQgKqo85eqt144Rk95df7koPd43JaW3bZVZd1YJH
YuxmCjRdh5KoGx+VRplfkCCY3QtZMMWLEzHgztKVoaHffaGxuK82xDhXzaQ38j9P
tfFN1qp2FYjeVT2syexFBDsy599AR2vq+rCxZ4SOCVbGkm/xLhjgkivXXSXE8S/I
Y0vk99+uKlqruDNB+BBcBir2RN0i5WzGfcbD8lE1a3epKP1Vg6MTnWzK3NoVpSAw
32W5cUZG5yJ2sZ0U/xcROk0Ej3UU1OZsEqOwzXw7JS2fGYW918ocW3a6ctSjVLoe
TyQMT+ksRzQ4qEuRtB38iD+i2v+W4fEBTTm05JsNQBrl2POrQ7uiNmplOyvMv5xg
GKyCZLHo3jnI4tYmNp7Ty2B+yyiFCnunF2D2nJjnxrZVZW4PuKHpPvyRGFVZ27gZ
zlMNH8LRs6jf/iq7Fal6e1Lw0UZ3gSWTpKyHcTmxP66S+U/avp+zFE8yoMlYxlwz
0dnP2cNd+Kut1M/LybQM3ALhU7hLkA0onLCTzYvdPQSmH+lHigGaXnMT+2ra7hey
1GT74zzAJ4f7ufhTZ+RPntfWS/ZraAFHN2a1/rYv0sShXtRn/vNrekAX61h4Ae7V
H1YupXQE3EspJzufR/x1qN5rv3NGktl5jFb872hCmUBp6m9eHOuCYMB8ZylSDrGs
Y9l0644to4QGRmfr79Vz3Sc8CiGpsytNqqdqeSnkkw4rQFU6G5XQPvBzeBB+I5JO
8y9rYvDzfp//Gob3GURBfVgOTrKtF2x7J2Gzw0tumOO5F71+LgA5qtI/kEH/oViK
OqdZaiQlfKv3+bfDVH2qUNfxe1e6rZvH1utwCn2wsaGFrNFXx9WDjQAyaHq90OnO
wqyivH6qsuQXKQFdAZa2Eg4tUK0Pvyb5NBUrhrJAIhVA5R0hLLB3Ry2ItdxbhoiR
3JmnJx8M7OtD1FuWOmlWzl9fU0TbU7znQImsPOWN8r/mixAchGeBy2A+WAR5JP54
g1+CcnG0bKa7VEG1CrxN9cQlUADsajQGfwSb9T6EeYU2dCwuI8dJHCpFOCnHybR/
KAigZuQQJ0BQjJ0v0JjGOnHtdD5pCneQ7lrgm+6/UrFXA+jierHdALw6ygvmGeHc
5tQeekhrvUWkS/thlqlCVvzHlyKidLLWWGk3Q/fjyJvIg2WyRzYWR4JnLp98kBMk
pztHJhAZqCPyUfE/+1EZok7dEfMn6de+TKE24OloW7gBSEItf70izhg+DfQreV5Y
BGKCx9UBOD8qjKoUos8ByAuC4ekEmlOxWqigmLKCUBs02gmyewf6Pa1Fv4RQ6llh
071nFhbVc/Mmp8DU2hjnKrOfBBuKGyftQ4MmeQYJjDfp7IEG8snzUo2/6wuyvQ0C
JpYrkR5/igGQowOpkCxA8+qRCftoqG+iVfZ7B54uJ6FzjD3rY8WCifX803/3d5mP
K1ROuaVMXmCGzUAtv++p7w57+5cu5vlgJ+q42yWtXQ0AT4oqOjUI6XpNhNObLnBt
Ry3HutO9Br2BGDobVoB/j2LUtCLiRVaTCKtmbo9+5TVonSosYmEspCM308HJy+10
tVqdeEJfea2fYG22fFIFQENi92pS3Z1q8AdNwIM4Mq8EgMK//uVmAJj5p7VPNnG0
UG38CCXPnZhpeALcnS8mDKtD9zfusMjkAWtY9pny+e4ETBbK7oi6eCAHMrCWs7/H
LjcoI4tveILpKGaW8GpOh8k4QBz4EhZtv3tqxir7IQtJcScM9u6Zb7Y9GaBA6WiM
xahXi/Ilyw3bFLaN2sADdAUMV9J85/gvIND6Tp6T01oXvtZuZlNItWSiLOQli7tB
9oT5KeGXzhNHBHmZLs73ofYjpS2kP8qiJd8TdPm+OHn9JA2iHhN4A6pDQ2Oq/gdr
kRjOyQhe2Qgz+72h/J75gB4DC10TDwwQZXj53DdV9d0Ty/u5nO2M3vcmwPKYWAec
/mc+haBdVJRhO4Cs4eFuXkytI5L1kTnJvFuG7ozjujvtP7Yuiz4+Bun5zrUpGdWc
flX65DLFn/5AuQGMkkwCgHc7TIfp1/yVYeJbAlQlkynEG9E136y4OEruvK94bp+4
k2UP1trlGT/kTqbLvBbV6+D2IvtBZKDowPahl6dHFOdooTBjKcOXw6BxvrUnVhhy
pMY5KLZwmV5Fxi8zCrl5Cmu+JpBA0nPgYAZyqx8CtM2qBnr31gCL7qS28jOSoIVw
whVuBrBE6rHy9zHMqCY2/IRtt8f1hWl2PJEkUQ0ntFDaWKabQEPjQbmzm2/Py5QM
EeWpQBCovOphHLa2K7wAjDdt7KglMFqA7jwd83Jzb86nF8XQ6E8W9T8tGzBttXjy
9USHIlzaLKoUz/DA1F6ZVN9CeZWPc+fgFHtFMfDUG8g7jjrPOW+HOqFH7PPHcOO1
C2xRT2/gWJTOv8lDlldxjGXYX3VgzOs4ULdYSf1qwyckjEgchWJBZO7NMd6Rc71h
d/s2YU2qNO6R9n4Tcv1kaT3EX2s9jxlDL6HfPcvW+AGaTrdchU4cDv5SlRM4oAqM
35x+l0sh/Z8EIh8IaQgj9Kvt2nov5MUrvuE2L0gSSwfF9a6j7OVcWPMv9YkQsvAS
53HhmBhzP1WWqYidXvurzgyhMOOXK2E4difaad9k6lw0IoBj8mK1cq1/N2j9CsUy
+krIefsWneN6JspB5LPdc0wjPYwpm9iJepJY/XAePh9XZJJCc5a45ggbkbIg45JO
cksfQ4Qvge5/dWrAG5HokGjUyvkyjLUj+87bewjJ5ScydbVHGBmy4nslNKV1+rXu
+rmfRS2YlPAF/WY0hJDPpfe5LIcdYbCNI6QQb4W5B3BTqvWmllwcLw+KY2wlNeFq
BVtyhY1qhmYvJUSdH1nagLtw6Q+3SOalrLAVxOg5cAcLFYoOhZ21J5rkoyhFfo4p
JLg9yRBWW85jOqZp9NpJJ/kLfwdWgw/wx1Jk+z66n9+r/u2UlRzwkNtkpLcTPEpg
vTXXjMoKPDZbfYEJA8zh3YWLohH0vHC4RjNZThUQu0WDCebYggn1JENmvER8SHRM
ZQnCR/Adp3JG5C9MxZxFtCTVYcpg+Azf1ug5lo6F9sO4QpEf7IfeP4DuWwL+5Csj
kOA12iDPK7cs/jI0HjYm8Oj6RReXdKOARc0HmsisjJbEA43zHfRCJ5zz+S6liyle
JSb+God1gMaIudjy4vQBApqVcphVVQFNMG9j7rSe7/Xxskd5JHLQoUrV6ZdUmAoB
waYTxMjiQBEI+qLo8uzKXxFoTxxkL72eH7CiTdpPfwnvSXx+lsRs0lDlF/rxLNT3
0oilPwodckEcYAebysSHWncwW1hENujKNZR8YGpq/Mj3FBUsBea6mNBg2tEOCOAR
wgS5jDoiVGIYCk54EIadaM+aq3/eHDd3SlfSp89qDOnmRAPn6O/fEkoYanug5lvu
RCpeKbh9QGfUzsgU/QBQFi6OHMK4GIpXcU4io3hQmFapAC0GpiGEJbpBA3kjTC+6
5SIopV9Xw/8yY4GMqK/50dF1npxNAwyWHjkEBR+3hytGVO0WsqZRl4vCeUn7dJM9
wUKNZOo+dSCSzJ5TygK4ZZMNYiTnqA425oZrVMvDooy+xIGO5rpGXxcrlCTTNG2M
TLVKBFnz+g9ZOCLRmmLyPaSSjsC7OqulIf0ASbMzD7jyFiC1mwQheUsBLMPflKRn
svsIlMdHGN75w6mUgOB37bzstHy5R0/IJnZXu/HXRI1EIYc6a2OlaNMJ7akuw9G/
KQV4QC9pYPSpj0CkwrKWPpppKVoxmb4wKMXxReUe0pyvZzBz0HvDNVicLGxpc13r
7pBzSCWaXKMyB0Fh0JTfwqljJdXykYRtQOtjU2FJWm5BOFFTLcbEAurNcZGT+9D/
th+sDTXwYLv32+UuYwTAmBS6fOSdAAS83jmh/1z418V4R/KdyVHHJ6XRTTeiz9FI
ANI/D2unQJMc8kOFpCfzhPyxJ3FL1zpGN8IHUrmOO3PHD+hIjKUKeDY3oaJmSBiB
bYV0aNEuyorITOZxEw2TlPHcN6gNNO0oEtM8oLHDCZb8/OcRpAKSu2iEcIcCyiBM
mqvk790O7KWlNT7oh4kGBb2w7owVWTcxnMlcnQ6zpruZtCyrqiccTqinPbqPcwYv
cZiv3ensxXR1ErMYPNcrlW/omnHsu+64RS705M8D1JHOGaF8U89VDgGtrE1r+VAC
RBeFp+dti4DpSGJx1PVP5I+z1hQ78GCkDg71SAnuEccDKERta8VfwhkjzqdK+nzs
skQTszEzeAmjf9rouKy5EvPfVkTlhsopzCpfJ5wQnXi+N7MJgUaoswKjx01eSYNI
sxWwgYCURNpYPvrSYT0rghQ5cVtFgF93y/h/kw9Tj4kI7TjbZaRBhutJurpf7i2F
wxGw4k5eG1iA+tx7sMdpNbHIkrDBGPVVhjMP5jgXlCV+ZgYugm9Ddg+Pn1HSZP0z
iCwymuu2AVL22EKa5L0BWQ0WRAjfWEiv1VZN3pMYALIWSrj4DdDY5xHNpIAFuQDN
l4Ph40OcWeQ84FrNhf/lT3NANTItPvXE8ckPMQ5SGLNESJtIKSCo+CH3IkuKUJ8t
yWT42LDbNjceqBFtZlPy4JEW735jNJhwKjn4/qhN+PK4XKF9FlPOfSdcncljQc2j
9vceKk/Z1kwOR8z6ZmQNCMN4UDTrtp+DC35Tif/mvaNd7p+JzDMG1trON2iwuCsB
i4AtthbemYukm4fLFN7zlY2+zxprDV/YgoOSdz/vr/0WgjWcDHC/TgkysmgBTVrD
+v6NZhAyPizNQxypoRCAK/f0oN2b19Xr3tT8y1OQNPXTcYcKbKYF36y0ReWu12LN
Cu491uOn6kYXgKp9yQtS3miUWvNmPpPKRO30PYemltxCJMhA6jUBCXOrSdpf1ZXM
RZ3QYznN43cZJEy4LxSPVLTX+tNOP4oa6dtaw05tIPIS5QJ2PDA7FoeVD/rIe+m7
9oJCVAs1OonmfWHKrNUAN6um8tmAOt6bqXI5096lScrr/1STaaC4D1X27vEIfTIj
U8047WywjhLTV5Zw9KGFPZ92BG1ANRIFKPbFo4o+Eqms6/B/kKBcem353zdGv5lJ
C8vqZeMQqAr8zqb88SXpbjLUtNi5imbAIfwQQotjFSN3tDSsvkYTtL8HPPmqJZJo
RJDuaJuKfvuLF8ILQIbK4OPrOIvwwHD1QjieRQwgir6lGZnJUN23AA+JV4L8r10S
0CcaX687DXUPYPeC40fAnmxBv31Hr954IciyHEYqZtBXMADOOrBwGRGgnuyhOY62
CmEEQiV2S4u4vt/pwvEp9zdmPEylDnGymyCmscWANo2vYze3aNqvfE+Pc7jhWZlx
aRQ4yVOYyj83xWiWH9Y70n8M73fJRWBidNu6nuvmUN0zQXttbmTglRcRMJg/ya2n
BX+f2EfuUHI+1SANIzBrZXtZFvvGn7ZuJqJIGxc0/vCYAY4RIQsbsX+uS/i7nTWS
tiUvgor9sCh/8+wH39K2ROAwdUacdBix6+KMUg8+vMMkkpOJMg7Zn180qxqzh1Bo
SEJ6xo1BfXNqgXPw6sUKx4qcxkILwblw17NX+GagfgUNmirpH4rK53fh8fFpN01J
kj+2VSjiUlXilT+WIuK34TAe5/DEhn97JZCIxsod78l5plnJtnWCvHsLzCVk/Shj
wB1RLBZkFGr5n5s29IbOG2GthxHMQ0z8V9mRJsx/HtIHR6E+RLjShMEEL256Ob5B
YND5WnvfG0ljXpC+ZL2Bdni5L1cxygOn1XYCgVEZTDcz00OLN3Ux2fxLXTq5g6U/
YeEKIOtvVUJDsBHtEj84gJ3wbm1XILrbOki4F1kY5VhWP2qGtcB42MqK4iBmoM++
LKGVVIsajoTatXORHVOCGveKNTO9jjCVbtaJ4DNL//fweltf1oEJNrB5uqvOoc2m
BBKe5w7uCMAgjxsnijBQ+vAuJoYaW6+N3wy9ViyiP8MmxQScqq9rOKcHEICFXWvT
3fvCT1/iqlXKS7BD9iYftXuIH3uP6NjcrT92kUcZjOa/IDp6hO2HKyIiaS2QHkyR
9ljY8E2gpIBGXTKm9QpB14Qzn72kBVNk6uVk36oHsAYVQtv43RP/oTWPhfhfJcVn
lXRWa9f7v6gZuovj/F6AndNs7lJvID8QdP70qw1M76kqdQ3JBZhGwJu3NBzFvBpn
wyIGLGvD7utmgQS8O3DjZcC05GZpjpSXTutraIrR6jTCB4/aatHqg5oix8vi1tLZ
3HHnelGcfeXTynl5JKJv2LAzDsrjmcipkY85znkJozS8HzQLSbn7VZ1ZNKZXhm6h
/bIPDbV5Tz9+EEu04L/r3T535DRGTpzFPj87B1wgZE4KV1DfvmUerXWZWTvCn7gD
ucTOrHwqTTshA2PwLnDL4VcE4HYyWvV2WmEw0MXtwasnMmsiD0yGn4XgtlKBXn3o
A27vypTIkrMcJqnXZNK2x1knIC88QnHvnMXXFZKFYV9lEVFUVGITee9x+A7gm5C2
yqs8EfYUePSvAo8E7QWO8n7NvWWo5atm6Z6uUVnR0dErT6flSWhACj8zJi41Cbvn
xj4HicMzJ7ipnFuxlDg+F1KKMQgSM2AF6O4v7NYGV0qpluN8y6R4B9uDwvFHcNJe
Yt/NAKotDlC1+UEZeQa5dBRLwL3aH4LREt21Cjj6WkakSVQobS8ajiqs2vsHozj5
0oPOvdpWfcGss/Wsdpg7PrpGVegD8kct4n4JzHfrIelf8fkLpwCRo2dhS07c6AE5
MbXGPSgeoLIDJ2ebIbZJiW3uNDfquRMuBThOWS3MtUqULFBsXEQ/9RmtjyMREa8N
6kbsKoFBkVwYgvge1+4VWxzFpsaV4Q2KdUSqsKtuXIQ+DsQKwTbQTALuohk0xTY0
8qTo/6NCukGtkx1ALgtv4Lw3vJqJEIhK9WiOgUUnwCKeQOCQfw64VCt7IqYN3olx
jDuvZD7qrQVIWkZWo8WUq1qbyAM3HwkXzShYWufOHOyMAAoxR67SqEDYTOHidifi
/hRNMZRiV/+SMyeqjt/aX8rAxhYeS9T7Zh8ObJk+uDPJyj8lJO+iQKVofJBUJZOY
02WyZsYtVBZBQiXmHc0kpdk8og0cSnbryhDqzIA/oSdvN9mU2j32XP3NVRkdofA0
l/++64CpqFGbIZE4RRSNHqde+iHHLlfqXDpLyCJw5Rvm+aPLZ/D5TI7VJhSE781a
XhwoEikvah6pjdv1nTUrbobI90Y6mZVFaJkxYLfjbjpnjKqwgRL3QYgoJ73uOB0K
9qAL4QQWXoZy0IKdjnZ+hefN6LVveaqujbohOxT0YKH2xuBMNWWnrQMWwX/f6ceC
2XFhDMKiGOkHssmsmoSSSnnouz0NwJas+NuiAMORZahUuY2s/UMxTv7FvpLFY/Uj
Hjhc9nRV8iCZEme8jeTIDm/nDZ9LboKc5wLTxq8GBCEOCk+Oe4AjZSjby9d7mYN/
dk/1zZnOczFuP7etC4uMZeZp2H+P/BfPA8mLaBQ9DXwQmd/UxC+JjBu2WdlKSUK4
8tGjKcAgDE9N/1iw+mQSTHnqekylydWv0FiA5b8ub4Qg0gZxWqsHM15bgCkQuv3c
nwF9uIcb+oMcTBhOCm0vvUPGEiva3vE6N7ZCMQ7pDBzCuxy3INUR7XwBLfmC2G/R
tIf1PHrp5HlTyFLgXzy0VEMTpqn6KWXoLS7m5db34TzTskk4iuae8vIv6so7qX8R
BXNX+Xj2hEV+VFnSW5L1FOjZvUOXQRapLJ2jBm5YtE0HABHN4kFy/l5m4vud0wQP
1roe3HFAhU2xwwBUnPhBm8IHwDLV2+t3Hk0kiQLlD3HioAnt1ZNajf4aH7xWBWdi
6HBsDq3FNk9XPiTugEdpTiQCzKB1v6+CTVG+p+vsYNQs67+p3XD1zxEzQTdqreFN
r+97KZpk0VF0BpW0yHOx6gVKmd7dHSTelbyyHqInwbFxRj2ipgYWAe9HhNPU53Hv
9B3RcKnD6gZM3U4DH5vaRLB8JDTEdKzLJ8RzQxja15DZVoVdMUlIBMZs550u4y3F
tAbD1Z9hjPE5jMqDpMcG6pLapu2UcDc/H9EPFGv92SJT4zNL4f0YgprVTAVLGjD+
iRXJ7KXnweSAxBT0sU5rEs8Gu6qAyBEYc2VdHVGUOjOPml0ZIgVIO9vx+fOXX5CD
7DPK1SlYmdMxzun3TxFcY95vf977QthV2JhQJZjgL2MPBcZliUmU/sfzwrGx+thJ
SrAGF5NOgFQdjCRcZKKVVFspLCruruFJbFjcWZLp7/WKoX2NOka4ltScq9pgmv7A
FOmWBUiKj97h6xCUn9rcVMR1Dqoh5ekqTisdklEEnzxZ30Pnv9bijzk3rdlY669S
TXHGMQ/o4n01OBMsyiD8OCQhrvIQXpVX9okd4u0yY6hpoYBlH0oZ3gtndqxX7j1E
mmttQfDhEPv9bU13aMSQ+dmGFLiP7CEwqrRdSSBP8nXcXAnp6nTzHVgYmpoJdPFs
bdPqhWahuXeNjrN66e1lcx7L2YhIJcTbs7/jX0zTOJvTdbbsRWgQ1/db/MNzCo35
fKEqTBUecrDQ8a4hRYSWcQ4YrmpmLcsIaEzZtU4LtTVZgZ3xda2jwfZf6Byg2Ucx
NIJ67AL2oacWV0jhi7d79CVQx2ZUdsslzvixTH29SQaQ3hA4E+AQh0sr534fxhQH
MBFEuhP+ne0/ACUG1S8r5V7qEdsC0P/jA9xSqNDJLau/P9ETuF9LGREmgaKWdzL4
nvdo4jqQ38cUSQQVd3DAGJ7khNnpByNO0KV8Z3+MSqfuRZIAmY0ZVlon2eN/pkNf
9NKCbay+SX2lnWMR0kV2Q8jjOT/aoWMJCL/7n4bGwm8yGol8uLNt5eY4ic5y0POV
bqMLRENqmnI2zSHywWlTbKeRnmsj6h3wfCGZOeNH9q4fb9FGgkPObc3hsje1ovaA
w+TAb0taph6XOGbCEsw3Unkw2T7ezaIx/aUt1JzEcuIgwYVOoYdlVifO4WoGWNqD
gbxWxuk3Cuqw7HB9a3954+t+DrEoxy+BBK7uMQXRKDgSO5WD+ur+QIougYHu69/r
6jLIpvjuq+3GCBlJAwZxERofi8ShMTEqTFAJI/Eb5qeNJ6JysMo/d4RPQjx3r+9p
zrAIZSziofGAGgFzJ5w8gJztINLMp6Gugmdb6t8JnMunHf0R8TJdFo75GDW6vQZh
p7h7tytCDnnl996TSSmbGjKrbJpY7MZcUKyXxmGNZghsYrFes4g+zHMzXTWyu43j
2cyCXSz0vidUGKzYQv7vsobwm2BuYx4+iHpplBJ1FPkHSECGNnb2B5j4dUao4Ksf
k4xJgC6T1LQucR1vVUo/VU2dqGkyDD79cXNoPr13xYz6lGPyD7XeyhJ4N5nCOdP2
rVll3egRv2EWmdPQiWVNlquV1WLQgU3U0l5/po6gFdmyNZSmyhLoWKEkkZ1RX3+o
RFNjoUWiU7Rmz/5lu9qYBhorz7Jgcr3eyjyEi0P8Y3ejrH24dzZzNKRk78T0H6O5
GXLXyXIu2D4W4XqZ3xPnF3ZJL4M06gmaXth2+8w2us7IP7WRkBCboGxjYTI4UPL4
075AbhaEzvYelak19dJmn1kotdmH5D/cEyj0eWbEiQ64MBFwsa2FIaiTdWuW3mcE
1c7K586hpelt4WLswEPm2RZhyf5v0Ev5YdzPr82riCS3YiNwchEG/KsT1VgRkBwn
8Y6OqAXmLgDz34kEiPK82GjzFQtWHgWJQVM9OmFYK3EvvUeGRj3BMa1nzMysYwGI
8RQqLGv+oTRuZYuI3CJlyn20Z1GzxZfFL0cks1hEY0hsy3rhPmfuFjFT6UfrxUEU
t2olt/26ozwvMr4pH5eFVjySO2h5bRiuFa483ivUTfh9zkbis/G8sgUjmQBkKozz
SkIMdOKCY76u/HJSUSyMI0z0rio7FFgvdfvsTX8EFl4hDx1OfBKj5iYR3Kl4m0t6
ToHjeGDM4n9LtD42d87ZQ8D+IR4Wz+0NuYOmY0wUFwRGm4RT/aQP6xYGyN6yITYK
jVd35KMvRH/9qpfvJ6umdoJ32oqoBWQavlYSxA8dsbUqhELGzsPn+F/2TdVT5h9N
JN+FuyVuQ14X0MQNPqqJ66pn8M6FB71f4opRCTk0DLsTP9IOy+k+hYadfEdlvhLn
GF5CLoI2uAgHV7GqOpqVSTcWyjLT6Rdvt13qiBbbdSuFkWzLCsgd9L8g4VSiKttw
YJQXjkqkIvCI41VL9TTxrKDAw3Q9iwBwaKMPLwSiPKZQ87jLIOeUF+T9OIHdxfbS
ZRzGTXVHZSbnSqyiJpxtr2CMdYAZXwVe84NNBNj3s5u2o7F+XnN1rrhL+IkUBPIE
OZiBr4/ZYOc1k77gp5AmQuhhEPLiK/HEIc147WKimtSDKNz2Pdayr/uG76hFvL0t
ecQB/57WcRzREGXLvx1nAhZIeXxqrxPPvnw69XhwEKMdPlhu77f6mfRM68zb3FYx
kKN6EIl9Oxw2WkuqhH5wttRppwA0/EpF0CBNUnVDhM/HQEkP/dYZziTbluhnS2jG
Sg+iG3g2PvzzT48QHnw26kSHvmzUbOGd2c87fThz8JjshgjxjGN2Zd9/fYIr/Vc0
VjqGhvHuvHWexmFdURsdNcUgY9+kA5Zzm/tSDnwFLRxm/IkuUTXzSa7RkqGqZG6f
GuCdroTmXzn3UBCxpopDUrHC6sZCztnAHMqik4yET0CZaUDVmR0CJ5D5AssO82Y7
2P9PHzT2deBmklVrnwuplq0NthJ+KUsLPnRboQsfVNCQzscfQi8s/O0DJv9TVgWA
022860J4N1khEz/NnGkkkRLBhTgUl1q9BjFYBb6pC72vMbWGLX1PPzTcQvtLpgdq
lNmEeQYtBZJyfVRkiNT0DgPQhyKwO3CHvLJSB3Adu34MA6tQZDnS2igXr9cEKZ10
WP2dDegjMmmtEyITB5GY/9Us4liOFDCKWNVmDhhutB+sDPcYPuN3PrUofPzy1Agq
GVUp703mCIudpBcFNDuwa6PWRpY1I7pczNamyYn+rOOxZzqiEN1jKotZ0bnWJ+Br
51wN3yeDgDAFzJmYE1lIjwQt4sBh0Hynug1useYETRP0clqEs/A5YcwZsesikeLr
dSsLikWsBAHTi0IJRm0yT8y8D+TV72m+crJP5WtMs7euFfdI5ITYRds0SnkVAn2G
tWNAWlZhIdvZeZDOmZ60w+1FGuw1GQLZHCjppyo3bXxXleoY713iXujJK7K/OgUW
YPiUuYWuquHO9EHitapos6rEPjeEg8fMd5jdFzaiLY3UP152DgPj9uz9Z2MANZXS
keXW0I1WzZPrttWks1x4+9wI497amy2mvk3uX5ddhMvmR8RZzoVGvJNtkk38GaoX
LRmoajsmGWIAlmAF87wcCiNaeN9pEm4gtPXBy1NVlFb3sLD2374/aIAZh3wXsBDE
Jl6Sk0KZEM175xsr1BSXrZwknsTU72WNoltWYjNDsQjiUb6cOof9N9zTlFPM9luV
6pGRUxFmzntbsDt/VjAO0xND+x8hAXCIMBEZ5xVnal9OD3M6igK+U/PVJ8yJT+cp
+RYmVgjSLREsBbcBtmJIuFKoRxiu/C+oZonjlqGsDDaNDEZwTE3PKsQrMEw1690r
NaIxVPRy2MPd4sCuQJx9+4BNfOXSr0FSn9AaU+2QxpDdsWh6yRk4jM9hluWyfwtt
r1Ox1XSl2kA3lB0SBaLWTg0YEWJuzzIvETeBTojp1nNh0Sy7eTgMdrnNHJor60uT
aHeOOhRxOnDlK7an8fWMIvxg3+3sD68pFez0rhjnEHu9coClsEwoxnVK9VyfqLYu
dknA3E38pxCWy2W7obghBRhlr9QRz1LEbA9ppSEHSgb4w8EtPQRI8gyqUC0mD16Y
f6V84csde2RCQIuwtWS2JzVPtWEUDDdwon/BMJuS3iOFM1Ck7fioJrWc7wCcqQZK
vpODH9lujZbw+6GHdt2ucjGyQM+fouvzFZLURvNlv31UlmRb0A8iG2ItIgQNztX0
abpgzkjbWyRoqpY53GHKJxr/h1IUNe6hxZsXQCSWfjKfjpRJeSqvQcEXy7gUQndU
DW8+V/CD+HRR5lF9DC5BU9aH4s3zStwEqQoyQnAYsY2ugQR7v26f98HBQTFEu6Sj
Q6l/tfSoD7jiWphGm3kZROyl5ttpBZMaO1um4Sjx63KEOqpzsBlKyHiiq81bCrng
is1vEXQRsiuy3AMbxHdDJ8xEUld8BSjZxZl5nTJBmFv4en/UD0B7davckW19MnRm
lI6nWusQTIyJhCNe52d8VaNhaINEmZI/heQ+COtAsbAC10vD0jH5kSmrucxOw6Xq
MZAtmGJ7ofiPjFCISl1vRybD2HifDB2BFPsP5CciyXy2j+I6omXETpfm5yPXDpQ0
hOUjR76BfZDH2mQjn5ldeIkB3X22cnJs3gj+kIHq1SDrYtE8rY/B4BcclogSbpWk
uAjJOCuzy1AmVKmA6jRR4wAfX3kx5/LnHOhDIAx0M4a0ZLkso3Sm2jA5Bf0NS8Ko
Zgw0+uYZhRIVRIme9SXh6bkKdZis20xPYOoQbUK1GQmus0/P8qDf6rDe3uj4pkn8
WACZlNCsTNB8oatbENc+UQ1xfW4j63oR4Pnu/260T/4q2XdyerV1sL1d5p5RQvmp
yJNqHOzmbmJ053m3WKh5wcYGQtpXToU7IKV6IGvJAk+BgZ3zD07TaELcwRemj45m
ElTOsUtZrKJV05DQ1W0grVtIsGVUezO9Q4ZrX90FAZRPFZYG57UM6d9dlmguqb1Q
ocfhoSaqGEYIxxb1whHMCrureqZ39wW7p5aMBWXG1gQJ1cQn6hG6xgi40rEj8fKy
u5pqdlJW4OGjRZiUywyFC2qX69VsDgcnrzYt5P9jdG5if64r6S7ciUWL4NwCZ6z3
pevLJmmDr6KtmZLjVzUI3zZJdCevdyPL77pvlHR8ZUYkyRr0njWkihcb9yoCWr6R
9W6PsdlNM+qDh1+NLEoKEtUkaIHikYvpZUF7PcZ9KXzO/6Rffqw9GUAmkJA23Zu/
ovqcmKQ6GO10e3hfEavtBHstdEXu8KndfIoMzob3iXL7yvskENAsRXBpYhh0O4kz
QSPlP6c6QaV9Wa6Hj0yd5Jydyy/0p84e5gx9GUyodbALe6ZO3rt/7fnfUBzcSbh1
KnqzxipfDRl3rJ5YLfFfWdvv2ulW38bmwgOL9XxrXi9uNYjq3WpB1L6OZUU170XD
xH7Ezt1s6njdCZXiVzFS87CEwef0qH0ixgGQrPKUEXxHCuoUXl0y2eu/VH6hm1HG
eaNXbZ1KzLsXKqkEKO2PqefXJElwJLkgImKcYFsqinpZPJJ5Ie6upDKxSa/Zzn5s
fgzew93nI/jZe8WdExA8MNUDbfpt/SRy/nbpxx/zBAi65NKFfM3O2k4REazwW+di
rZCpNGW15t5TtCjX710RL8O2VXD1+bxjweqFfM5iS0stxFP6DgzGRPOwu+tFaP93
CfyOVxt6GDWL3xILJwAh0QowNS3HD21HAMay1398NncjzJd17pFp2NGEFxNWpBNv
EVC46weOkVQx24Ex9OagMXseFyT5z+701/KZW93NicTRsmp1S8uLrpkHH4V6g9EN
/XZmVRePevFaPWxi+c4CvQUOAzc1IhtxoMBCwm24A6NYkZSSZKmtAUEbbwv24VIr
YIauF6FHVrQxQR2qagPYA21pqpY8t5E5JOxqUZqLzs96fzj/QpScwfKbfcKO1Qxt
2LcTu5/lHLknZ+luDNYIHZnbCDzCLyOolv7q8/h/HZCtPh7KwgnCElFqAtarntLE
8Iid7vkXp+GRkJfgSkGJaOV0rhIWcCv3a/Mjn8QmIJ9/Sxv8/IuXfttLtjr9uad3
w2WxNzJUq9fuOGY8SgyA+K/yZD0TF5XeRZ09yD40JY8RVP8yradLv7n6AxATasQt
KcNF0exCe+73ZItsGlifdRwKdJjFbPoszO3776YodC4nJGPzo4Cf4TWtpdwrCwZ7
y8HmnW9UbQAZ6rTa8hDcNYlGjSgKpuV6AfxBJJ+v5/072dSHQM/YG1cJZOzRt6tR
htRjJRUuUAF1b7mCOVp+ZxjEp5hQzFH2AK49ZvJJzKsAhxX6O0flq09rfYwY6PqD
Hu3yIo9bw4st7q3huJMTPLUYEGAhVNQ1TgaEwMg4Yblb2FwtV7wGZydTWoWnsETp
o3NipwR0qCMohOrFqyxikAjSCO5OofXN7FHFXyqTqMv1A6wNIsV/9ImpNcQ+W4I8
0UP/4nshfEwlPyRDNS9XGO8A2b2vPZdhy4+kUs1oQdWtfoXABG8FUHCoJNlyAs/5
ip54CrOgMV5m+S/ifEeTB0M+j2tKsBnwKakN0RPIpe0sq0trMZSCchZqIyR9FftK
7LOUGA7iGYssNuKWXTBwkNmV/3hdZGQ8PcfeqZmx+Pex/Y07YWJSUbaFjwzETfTI
cfcaOqYnQPLs+hvGTXJhU6AEKF0qh0TfO7WfrLJDlFMgKRkmdxFXGyfDns4uSotn
69qkGJvRrhyqwNcrAkdNEd+2iRZnziLqsLdY2jlElkty73MDliZO1iWu9jNX0Fzs
ABH9y8gZ5p3A38I86qEuR0NFVTiUOvZCN0jHMCA6YsqVY2fUIefqSxnUX+S8Lv0w
JtyCbHsE1S/WlFpPQb/8WQ0IqcejZujZPNYVLxVLphLYik45UlQvUzKSVelMBkYo
Hqx8tN6d13s1Ktt1I8hzMWdJcoAtA4XhWymLhTd3PRy8ez5+IqChb27OY5InMvfq
/knQHFpLSjoThKYEZMYAI+icWE40/sPn4HakcBD7vp3lwzGHp4SCSRc3qZsSUFHA
9kFEYixh74D6O6Haku4Jn3FtrKk2iPDXgJYHpxKNFs3JC5ZnnF2kPqfCvLxlD1cq
uCXfsp9VGh2bh4t1bli8fYxpnShmTFteVzyXenU1keV58vyjs01N1Bltoy0sG+xD
iHorYSy67o+c1rJR+f18wImr2HKF68qBWA/iiAxU3fB3LoAym3swdXT5t4Hu8OUX
+jwKEXBAnmIw0tYzi3RSrATYCPR3EMayA5Ag4NS9+/LWQVwjV08brND42LoQFrn1
D8l36HmJPedQ13tbLCLGPZ52dt+bPPLgAj1c93OMcHypyxhnPL6zPSFJ22Jvy0/P
tAm9/6ZNV/nIyRyQrJlj+bocdpWEW1qv+Mwt/5mo9U+0ezlZOr3enX9OeFU6Zk41
2CErgfiqToiyUksD2tK4WQGnYzmR+IZbtpHTlx8oFCwVy9KFrMtUN26yBvjSjElo
lSf7RAgrcoh4gvbqll9R9ZbaRt2Zx+db92ofhuSRQ1O01gQRu0yVaqXpcAaXLR6o
z3v3NMqvPBfDQ8pyrA9dx2L9SQsb6SSXrLrNAJVyYVIYL1VtMtsA2giPwr+RgefQ
0pa3g6g9dYB7EcJjbSwFu1Xpu6CrmMmWnspCoR5dtAd5r9gcdxXZFreaz0f4kCxS
qrrb6ejbRPpPVArlGHL/GRlxK3g48oswmBGdSVHjLI/rEYJQUb5L9H+IFhhRImQE
RPDNdZOced6b2hQREEOhgzZQmgXomtIMAgq1tUHFLsbOsM+hLwhVJt57U0SGWCAc
J6MqDluEmEWeaaBh38jnTebImYrciFq4mmyMAoggGhUBJ9yzV6Gi871nuwKP1/ZX
uwu94C59sTg9uR9Jgivcc/nZv6KQgP7Nzc2O4F3yc6az8DGY5usEgHgShL1kRkzk
EeuePY6LHYOpm8UI6ugYeqldGnKubv6po8XpXpaBpivffls/UYPd/mA9UYMcz8V0
d4JO/J902Ds8lznG3D41LEQ7h6klsQrVe9w2uHyUsMvFVjyPwtf3+ex8YvyoamQK
ugkmws4aFfyebH37Divrsa4KjVu9//fjhp0tra3EHmdXqq0a87gH9mKTfQxKckOJ
s2LdMB1Kb2890TGsPJFyF8jcos8cBz2+Xfk0BbkpVKRlc3Vtb5jXSqYK34RBSbg2
GM3aXmjYO73Pt4zRz67xmAGDpKkXcDk0KcRCrK6nRkrEMvdnWnJ7RcfF/5YtV2AR
pIKqc083Mzq6Ybn2N1od1dfPymJRbDcQteQMuTIYBB9hc8xcinHPfP6WOxDyO+0R
2NoP9dm3cgZbawVmljwxwqdEHtVdNiUDtrIjkIgKBgA8S/lidDD26WrxwuyoSVao
r/0hoJxQ+wEPtJI5bOoQrxUP7FHcY2Ed10h3F0RSxMejiYzqTh9M2jYVEtsddvJa
DGS0cASTNkTBihCYKm3i8o/pnCJra9rWQtRnWIA01ZJnTMXgObtJJyHS6zoBlhOt
NyBT2pc3GtmG9U+tBvyXLn1KmD4uRv4GdYTT+3gFFdN3BJCVEZ/Q6lEp7yOEjBtf
uJG/WWg+nHd15DDWdS14ly5RzeVWEAp+ALJV2dZ1BdTIbF51JozN3gKJaB0vajPH
KoZCMS5ZfTFjGdXVbEQDkD6pMr/MF+VfONvNYuzPGvXLdpPLluA/E0GvKApTsBaI
VcbiC1zpTyzuFp8J6bLQLYuAjKT9olRCWvzX3t/KPS6pwiO6av5aBFzhAjiM62ap
4bvKMFvFPpwHcnoic7aCv8V/Zkmt3aAMg8Nwuaoo34Ux4uHkKEqhy3TXp6rjMVB+
5E4iNPbIeZPIbejGUzTJzdAZ7m0SPZFM4J7Ts40JZ3Neu5qQMeN4S36mIjpJt8ND
z59gGyhY6rRDmD1n+aXmMuYzPnTNiG9Htz53o/8PPAsLuDIaJIuEqISBl99clkR0
+nqLdedBn3o3CZotMe8HI1hxSnO95kEPUswHmh+/N9/RYakZ7DZDVZQnbao2dTMd
Gs5gPz3nVT7cGnXRJts9JCh07V6WsoNdYQrRIQBIdIRMjX4YpvVJOpkqEq8GdZpO
lWqGjH3dLiA8pr3Zks2UVXJVs3YAHG0sjDG+97QLW1WBR3Up8sGi3RMQJhVaLJPv
vLbD/VByQm7O4hNDXYTvrY5xtNb/1yePNBlfi2mp6zVSeHmmnAYJzXrkFdjmOcb0
2uhTVlxtgrPtZEoJJkjzPIM2k6eaFUqxJcwekBy3JshrIzvqKdx0Cr37eKNJSVte
jAOi3D9oBT8nBA4wn9kSJ18VM9DYvO6ZSuhRvPoExVffz+z0lBO88K1f5KguhY+V
dDzh3gVWlHSSP8QJICNv/k/vHXPKBw1U8ZWrKxh0YS9PQRj+InJtb2hD77W029Ug
VDYyu29BQmVCnyO94PZY+o4bI9+2GCRBloTyTV1kbKzOZ3dHf4P5sXIwbvLMG60e
5RiYK3TIOLiHXegXMgwzhwYMZQcxWD8x2T39OoTOhkZuv0sbC1SHCMMAq3EGIIlT
jvkG09CtRAcu+esTFGIhPg==
`pragma protect end_protected
