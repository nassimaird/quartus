// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
j8G+i/fw4/rmk6Wn3zRWhlJ7rBmdsywzvpqIBm3m0qTM5TEqPnZ5ZtB3F+73vJhIlrK7plees6UI
rp1pURm4SArls/+uS3G+vTbAr+XiRgTYulN6QJBJXOUgu72hhz1BmYoqsYQwmELyEkwv598vNaj7
YD4DP1Nx4URKH6bUKgVJ0g2rgOpcSgoZ+Pl3An0UbKsKEHCrisoW8OHiigt07SJea1TSwqCeRk+g
ANYRo9ynEHXBxRpQnNrXeMgwAP7bkOGSJWMzzzLcECsRmjzGzUaEr+lRfmj25NuSslnwIAbMmDWE
yDPRclac72/fPYvsYyfxr46fZERx+kJrNUg9xQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 35248)
ocCLkZ6lE6JHpChAzbJLiIsm9CyuqOfEA25T7FCxFlW5MKPyE+qa012aZ44fFy9kmUuxWRnRy91l
hBVM+OzftAg2yeZMVCmz2IyEc855Y3cKcZ6oxD8HWp1HxoG25jeaZOorodNPVyDB9/3aFLATBsaj
aX+Pe8zj2Gp1AbH0AKzAdfGXG9hHVfvPk7B5TNqkp6MT9XMf0wIUpW7jgND4kgohYJ9NvJobvIhO
iN7HIt2yhzkrkWdwuBidQHRcNuNgvo6Fb7hacSIwoAqfQq7gVvfeRiVVETQAvJ/sf2dUTem8ZHI/
cZ/hnt9Nm865lvVl5Fr79WiOwduIfhnMbhbe5c/XSB3lYuSBE7ASA0a40msZEkWUHyF98K6z7wSr
K/jMFGC6cOvxWhpoxcrdQTHhs679jtW0Qle+/41zVThu8e2aDbkmWqpXBNzZ8t8iLnlPBGUsJv05
szQQ95toytA1HmUOMLUPVO+uXAfo5pRW5OLsNYiyaGV1nLuQWESxc5to/fFWf7qiE6FOTCyaMAxm
VKnFX6oT6ZkkuvrZVslDcOpdxOMrdl+UnlGnRPo4ykRJGQTUcd59Obb090jWb8ZEkOQFdLu/ZSFM
GkopiIlMAzN28cT2rWJSDXIqr28qfphzM7t9q6fTRbky+ybD5YfQV5D16eYp87Hrq7j84vTrqbf3
KjFonHApT6DNcyjb0fudgVZzxpDe1sA7RIeYx+xdFqKPuz5lHQGUbzTEKZLhFm8QyAoI7MWWp+Nw
bt9LvJjtTxibzhG2E2FJd9B9gBV2ddqWzSnNqobtS8zWIQQwwB9f4hF9/EPwzQouxUgsizozqWxH
7/EUwzO+Z37xq4x3hTp4VnWXVvZBxnuxOnAkCDQEbHx4FED90IK9RX1mq8dxnlL3RqVbhaW/fs5m
RR7D6q4lOKpjIS+ySu/0EVB3gt2DyEXPPTJoV1zsG9zsE7KEkUQLikO9GiZe7ti9gxNZgVeA4bO9
d7cBD4Evj8uI+ENaNPXwQWHjBSSuMOkfIr7WjJHeoU6pHdM84NFI1gYKx/Ye0q3TAKiYa0UeI+U/
bqDEvxMA+UPd2hXEA9AaRrwGLo0LIqijXUY2/gCnOKYTPvSezeaEPiV4M2cTzmextcZUQNJlbvg9
YL0iT5MNxDZn9pDxOzx7xx8wLOLx3TrPnC11kVZMC1NbypyQ9UDtgTgeH7UO3zvkKDmmSs3SKdaw
L8qBeCzdpD+xB5gBjviTggbFN0LO5FOgGPTZNDgNqldqMMU0FlSwH93234u8L+2/qAmhQjKnBVH7
/Jemd1A6Waz6HfXefsNk38XC3ccOhG4D3/4PFQYvt6qlyCdvp4AAeXMlWqCWmwgP4XdET3fobc2h
SynZuy2YRPLyXKty3m0rFNloVl6ycO+ixBz8lNFEqZQhR7L35Rg13cSMUtm5nfvwSjT4AJuOu4YY
G/1JxfeBMcukdlF3nnK/n8nh8CYwQzi6Edj6UUbnIO72PguSQ7ZFbLgK2r4tm7kpncZqj0jIWuoZ
HT1Iz5MuEBLETH60+Q1e18vBv50ZzzvuWnmX+s8dRu2nMByOP3kf3gsW/YGMQx4CXTkW5dx78gkR
bdcA+lhGR64MnI/gqwKZO/X1LtR3eVoAi7AgnO3BXprcEbYMO9SHZsCDMqcwdwgn1e7as76z4isQ
QpwbOt/C7UP/JWIlXsO/a0AAFga+QuSsxJMOJgJ4zXvGPrz6/oJdWge/k7QYzWYMBQepN/MVl+dK
nHS73KioovujVmyoQbwk1sptXZdHeoLSrEOLbDDY9pwiW8haV/AXdpwXV2+GRBg13cHESw3L++Lc
+UvMydcAdefNhVy1u283YF+OX/w1vwJn1+vstHKITeJSvE4mOaPLUera1sTZpjZYyIJPF9IIN8E1
9ZNMfvuePDSmweJaOQwnbAhpiNPJDbqybtuoty90txCWSCng5+D9lvg5v//TbQalt/l6KGlU6ZUY
bac5ZOjYl7WDFuInL0uXmhROM7ZyEcfHKKHIy0vwf0LdMpfIwetiO533DMDC04LUogwaw4GYoOOc
+uUZgPoxtxYQ8+PXjzcKOtgjshzl0+5WeqqPTpYZD1u6wNi0xG9VC5op9URuBGIetiPEq0dJbaZW
TvOHGv6UuyXG83fCPBB78kOjoz7g0TGYazkfNelv6bTAcBwzJN1YHh51VTu9rROFLSYogl8MsxCt
lCuFAao++KLw5Bb9bZaFOnEA+C5L/CKBE2FgX185F1H3mrBWUU2H5ZEvbQtYqK6kShD9Pp33Uhz+
QShT0Zdnyi4JZhvpws3o7zW+cYoVSZ2WQTvd8XgopuMgXRePPiNKIUJarLez23gF0w4WZEajRA0r
9G0bygZ8P/4eyw0xoIIfxKDYXTpUk2G5iyurnKq9G2yPmaY+x6e9quRtYEbbs2zJQtBiSmg0M5eH
GNhzumnV5RRgr4T/NoLTc30PwZ86/5BQgwqUVeHkYluXSGyiKyjtFpkSg36icIyAB9tC21VfVk49
+j4+psqxXSTacgDR2Babzwwcslk8EoMXGmWYlePYKmNwpVU2dJaZcJSY6D65bv2av00pGGTy5Aei
fEGPPKb0NMOGRDiDZs4gO7M74cbntrPww13bvO7L+cCUEV8b+X3vmt3GI1177xSC/MxaIn6DYd5/
q1CS6g4c1lq9F7/OpwG1JkWrzLX0tdFDP1wecdQxEgMTuVDmPPT4Rs2nLRxDjmROXORHNhI7sKgv
CwFGt/HUo/NhKkrn9Mc7U9xp4WOb0oZW9jP3DHuFMg9MaXbp7U3WGRxcfjjnyOYB0QbXzH5ZoeSm
TdcWsPrUObMeS0TvIWHh5y6ieGp0cfngURZkzqipOG+QJcN1FkeESZvhYO7iBFy491t8PdXe436+
JhAbU99eFVQRQOKRRh/TSvztkNH52k9Pzy7rvbHFgoMkpDAV5Nf6tYlFcjnVQyvkLZz70amNZewl
a/jEiRbXqETS6t9uNknNgytcUmckoUyl4EqroH7U9LHnMqbPlLgyab1jjfwxTzMdKKP9ugZ1xRsx
Et1smPFK6MV1OnwKuVFYU/NqNnABBFhFJinj3LcWW0amP6LR5x3FO7LUzQOwaotWWFZG/xynE687
lkZcp1QS9JMv6yCLuVF8BvdoqsqLWYRAUD0xETwPWOvRL8Wr9YKfYsp2fwtCW4bAM1aS5VVucpmF
zM44TIt8rjejFcdBS5XnDcaa3c+JnPJ8NKhzyTTwUx+nwZ0jPBZBBDX1v+cSwnsOOCzu7qDZIPR+
+hpKXRpseFCbHUDVqHVEh8Bimq/cLMECATgPN7KhKMSR5ShRTbawbR6GiV241G1yPozZ+l0JUjlt
sVNSTFcGvAvPM/l870IQFvHlyWysHb4lmC9990dLmpVErx9sy2dQdRJ3gq1FqfoMBcTSWWSH12wE
JVUA+hTfd/yUUsvH/YrKtIP4NVwgkiB3cIfUt0+8LuTNVKpfPjbki8v2XwWsAHBLqpBDEZ08UfAY
gHUWpSvmgb4kDiCwjqqqjUt0bUBq5w3K2ESdlhInlBP1dl+BA99cgLzvc7wAfsBVJnWlICLH4G19
3zIr9fXQqbcB0f5I5aAjg/7pUbD+ThHhTbenY5jlhmrxua8NTMbjOPkw2f8FdldU8Z3kt0Ba6Fak
YqervYYIOq1A9koF5ZNYRLMhMHA2pFZPJXproqIKc+StzwRVQtvYwOGkLZ+FmUqfG6XIj3JLSOU2
zeb8JIVAQunej/DG+o6zR+y2QjnJaSR4Q87TPg0/i000JJSgM/Aug44oUItLLHGR/0rHL/1ZjJz0
jbiz27Pp4mItE1JVdmb7H9tE4B2rLoOVQo9rNbhtEHUfpXM7Cir0je1UMQI3NIrpCtkMWxSCZUTq
TMZ1Fm6QE8/7I6hihNmKSZfwejqNmBMm17qJQdsO5G43axAbbn/HDpSQCvNGzS6IfH8JYfTeeeD+
PxaEK3WuzghCLURWe6F2o5ZbuUTWh0qBCiznKPptRMPmnQW7MjmZ+MFP2IhJplLDA8LbqM6kLoc4
2YSW/VSU8lgL16NMTipjkcJeJasX4Hz4esPgKBmzcE/8nlB3+cz2oNjsSPF0e/6rCRtVXk3x2ieZ
ZYSKl5CKUifPX9m1knLpQxN1Iv6hIbV3rrILvBVMU0ChJDcnmtUxgZquEfZ6/JrMKcZPVulku2p7
lTtElmPpcpESvY9V+2EFf2g01OY39rGHab0VXgPXOX/6NQorgD00bipOZnaKloFLSK0yiKPX/avK
jWLXuZ/HpwIpn45tZHT9AGDOUpsOVn7t8KA7PNzRD7xVzvcsSX7oQ7K3+feQDFM9M5NPy9t2CKOr
bpqJ758J7o0WqiyllfDi3bWxdvP26zQGEcfKb2YNOqJ02pL+vZ5l4GSsltbm0u0a57srOmkkXRcA
yIqNjCdXMO1ZOWb4Bzch8ZSZVXXXOC8XS3t7kobLnZMgeMrEto/5cDBp+B4VrQti7jaNyhhJdSGX
dYYeLJ+OtGijJ2Dvg3ODyHeAVwBcbR7tsoJXVMEahi4d+r2olrGVUKhZcwlwZYT9qD9/Cjs5NgLv
cwMyFrwGVmULwnh9TPxjWWayL3R7irLZa7zS7xqvl/X2k452q6m9yZEBAp7K6KUmDIqspOJuIKG4
t6382t+81saORBSiY//AE7rtsBkLAPv8luHz+VhV7hzVPT7d09gPBsig/vADjqYUJ3MVkvCQUnBv
FReLolgFz7RN7t2QKsoO6aq0ZvAzHKWE98+ODRdumkgFW3TtvJU1YAKSDYtkVivwsSFaFOL9XJ23
/tXj7CEKSbJxHe+OWkbVs/Xq+DcJpFEx89fNQOVqmbvOOLWfO4O2f3/txMvak0rw82ykp7XQZRF/
oQ/ETQrqxpG4zRVKofse0rhajQoLzC5EPume9M1Iw+fMswnxK0EfAIURGtIF9da799Dd09TNR0ZM
m6YC1jUoO6LePPER2LuoC5PvtOtzkrKmByp+rcdDCKDgapY/NTDmhVs2mcXxUKujMngp46LPjBSy
d/6CwWdv0b69e3E5E0gtAbmXPwUyLu4AsloDWj+wEf5fh2NFo6JmzFGUUukHX9C2ughRCgdFVv3b
cNjmTVjfWrSDMQk57I7w4B1u+53L5qtr3oAo8kq96Yp5qLXxawh7HbpfgVqy0pxNBkHO2cUXUmOk
txbCevBZyAql2I+RXE9V9JnWprSZ6BU9c+3BS8HBpi7ExJSHT2W4XP8s8IAsNQ8mqDrnoONKTfR0
AaNpbRf+joddO8ICJ1bPxTqsIyqJJwGxwULfhY8g/VRyaQKzXLoTDkILf1nRTlpclgjVvh1T18n/
YyiB+QLjmHqiSaNt6V6rix6/z8UEQRv0GeGzL/qOjLo6CCnhE4j2VXBhybH+P1fn+e6CrRBLvCl+
Gdre+giGN2Rw3n5sF6TgDnzOa0JbGeg2tkXVMqjPsL18KQugDETT68xv7zVfCBySho8jwExgpPT3
AyFhvRyLMiO3kTC2C9ih6mNSScLlpfOQ281z8a5h286aiUOXCLl47dlaupNA7bMflUNcphwmAo60
K2uKGzkTQNHRD7rGTVU9gsVfKHT68nyJ67oLyywtuu4xQeUb8c5MZXy/wdsrp3uCoHcsOb1tWPPv
blY9643M26VR/SybQQ4zesDL11AAsRhbwyPy6jdvj/J0/Ly9IpRe7Y9rjG3/K3XxFQvhCqpSJaV8
O1YBIqad1V0ZbBw8zC7dE/T8/ZKgwUqEzTafUjOl9e/Q9g6ysTtMlJ4j8CG80JjDkvZ14C4UC+EZ
w4IMxVH3Q26pgImjV1pii2F4fkR+CyO6BfOrh1f2a8JHq+2O/KA9jtRVemrWG+KsXRYZMSNlQEVl
QI50ycs3mqhNYN+ZoEMoowm6Z6ik7yWVLniexOhgDU8waioqF9ScjC85HJJNl40k6taff91mn9Qi
mvRctNjPQkgdevlSZvNiBuvrpzJivZchSOaJ6WDFhDzai8G3/+1skpFw49zTPotTHN6te0rEYT0R
W0VxMcemjfycUMZg7wiFR85zx9WLvqCwbx/UVNso2tg+ZWbmGbP9ItCVOh96XYQ0YZ4gyu/FTV83
VQ1aFlaAxmv4TQmeMjFBLfAfB9GU1KP9lQODoFjElEzKYWMieGNf62TC7qYWWBZ09V9k+svZyMVT
zA3C8njnwBrRG4fteDWPc6bqTk488jet2GleVSm/HJExtpwCcm9A/1Onyfv3lfwDAY1XokmUxn1s
lNnFVI25Iwa0/PmScK9Q5zwGiUT0lS102vvgGznWlFWrHT7rzvVkQYlv73AzyOmU1LmJXbCJfwOw
Ok/i6bd9yFEE8AX0SwYrLJLmUrhSZq5sTTbjvWnl7c3jF/NmyVEZ01JljQY3wu9vKVtWg2+xflUl
2fkxOg8Q0aDzfbqByjLYC3rzXWLS11Mo/cxHk4KyRio/R/ehf4J2DMecQWCDfAPjfJOfZXjtKdjd
oPAHXDmSbjFIkj6c8S043cbCR2LLVGodUhjzyTi2SP7F7i8ZINhhWgeSAbcFmwwNVxxLLdXWq9/f
kFB6SE8xs/Mo4ajocrI46BpI5HhZloQocNG6D1Wuj3oQl/XyDr83LkXmUUms5hhSRNJsM4vci4Qf
lCrYGGkdSCT2NknsCZ2d6hOpONcYdboUcTrGzeIBAjj7ORz58TClfc543s5tfU9ljy3WqZv9s+CW
Q5J6jjKou33IF/xcJqAdXp99t79JO8FfpCV4jEv9VPED+o9UozKRFhidIakFWHOPYYXu5C18Qv4K
dNurEjQfWeRBZGkyDqahlrJ4gE29oeTwkgiX+nlI6aaT7vuwQqz2s36UDvSWs3dX7IsbjO2eDHp4
C+4BRVKpdv9Tooo5rgq1zgBrcxAIU73lNEXDpdFwN6X2IQXtiAhYQ1ymACSOJf76vSyv0b501Cp9
rBh70+X89+FBZtlMrcTfJE4ZikB/MgpvmS1I0kq/vomzF8hACVfwsqqQyApA30srwf8/lsxN3iQk
cVU5l1kZRTVd/pBHSAIm7lbwMYCAd/dBlECvpMSpFV6BTgvG/LNfUEw2eA7dt6udElaOx+vK3bLI
xHe/Z/6tH+m9P3fBsgaNEDTVtYxY75vYvWa6zJQe29WzgsxSIDS6n3EGw8NOoladBvJnQqPIFs5M
XNL/sbS5CtLuVUFERbID7jct08M/HV4fBx0HQ4h66KS/zpk9sRv8mqDci0DNjYR6kq0uSMQEwT+U
etK+pZciiHEm2wHwTq8JCziWUcE5PGh3aPAL3Xy9Gye0OYziPi5QyBrWfXg3fBdeHPvyNChraAbN
K52XJUQjS6zgVYmNL2VOOoFY2bSU00oJ3gT+Dn6o1E1lV+ouBd5099/PNAJcExGETpqgYj8q++eu
VPWSeILSYBmflE+b3zXLlFtOg99S/IXvrSVJ6NeSd9wg++cRgJ2gDQjuoNfxM0YC5iF2oh4P88Zv
3EDFP68FiinIYDbBzCkmePZPkhYDnRE1MBoZmbXDnN3q0uohguLbkm6O6zN9VbGSpcDEDw0yccpc
Z6nI/1u15D0sjn+8Qmc4VRCPeSB20YeuQnlBXfrSbq40/1jbVJKaUxgeEitawktpipTLYseXTQnN
0uIofWmP+JPc8rYgoGZKenTProA/+MxZu51/PNzxwZKezJISHLbg2lu6BNF6YN4zcI/dXy4JV8Lo
eXdit78o1K1nO3jzFQ1G/HDJvf6Ak4SyJTeyz+rT8tAPzbJ4oDmpixe4hxM++BR+8B6CPCR5NUJ0
AIFfcyGLAiSkNQhsQBagVyvQDzwzrK6CmC7aIdmgmL2gZZhesyFZYPQG4tXHGnRlxh06sh7qc46o
OLs59EdfRgYc+0L74jfOPlDbvU74/CagktDFb0UVvR0Jke/2Jo050Vy7IFLTZ55ORgFUevKpyimI
n/ZwqyTe6W99vbssjqdEcXcVdmTAzE4GQzUTIWl1JygEvCHKL1if8CUtyUrx+FpHjBD7XJtqzKua
o6V6kt3AAzVqICuAa6S3sfy/zGfj+BNFVWmoDFLiCI9g5PK5ictUo6V8l22E2FNgEQjugVHRvto7
pudQ8Ajrq97iifR3wiDpc7H9VZUMw8flw79MPAsAGCt7aCrA9SqIrxX+p2rwayS0Hg0hUJcSZgrN
cl7kycf0vQ2bRH9FSqzVnzL2/CNepo3pU+reVicDeVaZcgHXBjh85gqa0/iZnONT0qv8oQ1DHSkn
vzDV9GOfrbyygZcU4OFS2yi6qwQnWZdMyOCwbY+Zp1GlFvyw5Nk1IiQDd0O5LEUxV6Fq4T1u0S0j
DyTBorw6mgWGPXirU/Fjo4D+gQmXbLMmmsy+LxgbbXhLkQXD8IX1RKyGEA2R+KQGkbJ5EKvcFR+f
f44Nuhg9J1el7XKVNPLb3nZp6uIqU6nKL+Y6mpIJM64oNudum64fYgrD+9QjzTo4IcvbuQJ8HAxC
BHUKAcF9MasZuPX38pv3gE0hGxfBr4+M4s2kO+t0Z174rMOeBSdGRpmbWOytAM4pwvKYmLHAxqC9
hDWf7P5OmOVAMFgYaoIOfY0lWZIp+7Uftb8FDtKA80O6sXNxO8ngDJHPh2E1TOxeNDrBzBuBdxDd
xb9jxF0MwQIPSmfWuAszreyD4QjHZX4wEW3FgZ0Hswl175EuSSz8c1DeVzRT6WKpr8XQeJnxCuzB
CQlzdDw7iSPGgZobMofklzb/45bCNDY+prI9+nwalTq3nLOorTNHMw8dKjwjfZoNY+wfqTkNNnX/
Uo1VVY57la40g22uh4EFDHTIZ46R/EOljGmq8SyA/hzv7tsZe0ddIHRcDrBg7ByNCKdHXLRx7Pix
tVgPZiavFa562kt8/UK6ZEFewv5SLH/RJVsYDB2m8+Qo3shOMTEAzE7kETvvGcvJn5uV7bBpeFP3
oWRfcfPjmoQolC66GLJa6v8ZCNhdnvM05+dHiviIwrP3qYpUVa14Bt/HWYyM9232y2dHPULJ9Pqs
e0kMquK7mxebASSMBJlOFYuERkLlwG0NRkSc3q8m3vL9jdFkssNPMdVLYjFweM0vnJylVZNZ4Jrq
lc6Kul94ZfSyX2d+7h/uoGXTuiDKJ0ZfDGloBcBgfp/I7SNKiM3goPGIeSrqNivcSbEeJbuI0udB
JJQPceSLo6I/DIE6kf+4luDWsr81W7ozyy6QGsTn3XeL+tX66hOHW0d37OxE9/aLyLr8Sz9DetyT
RwyH1bcJQmgYTSgPvtiSZHOC8or951OZB4s5eL6G3cAci3Y/kDTZVAoLn20Iz/YCGZXeCSD40Z3h
ERWvOmf7FYkbjS+2jvp2VVCDGG3afavhwu5xH2TikOxlFEcVJZJWi+t/p59khmgzq7kcb7dOIk+N
bZyC9GNwnNtwCzKzqpiHarz7YHCiRnF3BtwA5g7twp2e+BYXDbl1cAdCymZaZ8OmbnmjaoJDt8uy
ZqeyPItSqrWKgScfIUajztugndkOnVeBTHkWtVXyLLO4vUx/z3Xr24PXY5xkEONewZ4NiiWUFin7
g1uJlGNBJsCY8xVU4oMzqFiAqYjdresQBDkkATv6gO+U2SNdlPFUAkzHQuxCphH8E/99Wk2RccbL
w5L/gSHmyPTcPWWmmEWxucRbHJYgJEgvdkbWF0uGxxx/GNwPYEvNN2soTaPslqdPOQoPuxi7AH4L
gKsS3op6yZbQYb6JUFjK2IVQwuUD7Cpll2DrSkcmvt5D7DgtZcqHvYiZoaGkD4AEhdimVbnVkAro
U7Hj/N9l0FKbzqOqrc6fKn/sAEuvd0E7j1wAyefyTzwB5JXh/EzAtuHQGxWYPzagiz7kO6wVZHno
LOVggFbU2ckKc1SwoSK8FoDu/oTNGBaW0P29jYarxCNLn8wuI0p5AUPPN008NpK6S5JWqrZokmZr
Upp4A+OJ/WXPxGGV8+2wvVJwi0E8pnZfgdc3t0+6pe6ODw4KOQt4gpvIfBwbfrfkSA53VWOqO5N4
leBYQ3S9CC8ucNdZjaDjjYPlultsYaMddxZiZZN84C/OCkUH0/WiJXogI/10DSAk0s4fXikhtiad
a5rohOmwfkdhDGIOqZUz2qkXPzfA3ygA9cMqIZ/0ni0w+k/nVliDiGnPqT8QjMIMhT7WGxfrdwdS
q1bSoSEjo+9eY/6gi1sse5YwZoSCy+xM/a5kFRNirEG/YQKY2atd000IrlGrwLnlAOPKMwxvn0VZ
kaJIf5eTQw6yN16RwwAcuBRXdV2LMcQfkpoUqFM3ndo8+kc7mcC3pn2AE3Mm/mCleZZw4pLkwHAT
EBVHVqX78bQIAgFjrURPmckeLJP8mtXhkf8qqgqZ0ksLKSuA0oIFvysgFL/9JZxoAXipI6PmpNFs
qe3pwcEXdP6da3AmlK7GMM0eGGYSO46qw85gX564KS/TEm2MocQNmKqGOYUgOAD3XH+iXApJSZoX
ZIIT2xd8mDQ8qY0Jk8iccxe6q1H6M6mPgZqbbLo9RtlGW+exqXHFNnmd4HziL2bZexHHk5+qhu7s
zdy697tLF+Gyw/fQG/YNecGP5vFKNmybGefIaMGjOVR9SXNkdE/NJhH6/rPOf0XB07mwj0IUNGZt
HUdsOqEheH5Gr7CMfM30r2QWsN9TPEnU7s1H0aTZ2INKI5ge1B/6S96xC5bVPhOBVo7dG6Oq6Lh1
olo2olfM4rDNQQT0svrJ0vc5chMcjlqAJ5kQ/oI6AgciRcPNK9MErxhGQPUDTK20wLNh8R4QmLoQ
OfNgpCUF6O+fUMlweRZAQTWfKlYLfigLldOF8PouVv9+BZ0GsE0q/CyRqMsfbSc4ebVD7IVCMmJt
IG2PmPQyNqD3iE9UVTvgKudC4uSonUfTL26iQBL5kvxcPgNZ91TSeCfcTXWN8K1fH418Z+0mg0tX
i+yqk8qs+DDTkcsZ4gKulb+kxip9oKU5en/JU0dBYciUW2aO9RvjIc48qwIRPk1PBJQXMOzKAktR
p+b0G3h5cE97V69tD0N9lYHCbzQ7Ju1QGvLo9UVRHcbBRIaob9RnlGtG04tYron38jk8lN67k3+B
QYgF/2XHdtkPZQCTpY4DPOhGY0X+70AYJqf3nLxt/h5eg1sfk3jBpAMQQ7DFABm1n2uCQuyGF2NC
m/awgEbwQm+T4w8YheP98gpUlOxBHVgM/Zb13Lr5kaKC8W0DWSV96HlZ9ZiESoyKCQOAfRvwC6YW
a995XfktNStbtbyOoyyKTmm2BJFhxlpNOEyi/wFOSlCYwjMiZxmCFjjWEgKCpqcM4Fe75/+WTUD7
qrxCdVxKLTJjUOuiCHKfDwrIJlkxhxUpupxNchMJgo2/gS2uvO/gf9k3GD7N/2R6G8nFTzeCibqB
K2AaT/RNF992m5FYh0sLl2iu9vq5s8f9uFxzPEmNnlD2oB/8whPlJBrRW8euCKnvSJoEEDrxvcAy
6b/nZW45uMhisWh4hESsSaeVLXDGFE5MZYMVq2DJUg838/DAaeinoLIrObgFokLkF3SClHC+tz1k
Iaxn5hd1QCw+zuPfsZovdc+kqVCEOUsWj7P2xouuu9QBp/Fj338Is9noGEasbX8YtC5BgbYq8uT8
65InTDU8EyKgG0wLAsbeXje3HWwRB5QfEOhX8PqT6Zg19ErlAog1tYX5uyckNqN820Vrp2YMOtRK
IfPI5dQiTuYb0i8uk6iMOWC+uu2aoVzzyIP4XofYJpysUUowzyBGlOdFTwfFd39G27klR8DIPra9
5rCt0PcBHPlqlX6nk5KcHqJsstDM7oAxYuJD5+ozPxKOevuGq32b3ZaiWCSZCUEMkhFWAd8u0vDb
BAi+paiVtmmz40ddW3K/iRxT4ez+cQ+zSVLPcdyxKVODzxoU2hdizJK9xuLCZnliOiUN4fhLAwNG
8SuUHJaXyGS/lZAhJQfI8lGLUp2QLNTPmMpHKk3nvIcIwj+IG+U+9c0lto1gZt+LetMeiUoZNlJF
uG28lzaOHEiRQV4YfX+YVzXqP4PSxbRjVu8xmFLR1hpWCeOOdnWChq7tA8F41zPnoCiaADuKB12a
UVfUAHFh38Cs/50zKVIkex5KZ7sAkFeN5T1yUIqLbgpxMD0SiGcCeiiwU4PyPo0cVw+ZRCnO07em
bGwS9FA5ILoa7fmeVQwV7fp+TXmuDswVlNUA/UenoyHDpUthx5x5p2xd5Jw8EGJWGtxZNYtTzTEw
tGe82Tfo8n1t29C3c2OhBIbEQ35p7aZo90rru1aHz12ot+Y7j87MSMEi9J+qchHXwIpS+aGKtsl8
w4C80cev3zUyTXgA3RtU2SY3X7J5qVlEcMIumSmf6kJfJYsZ/TCxnlo7GIk00whLL08+ODilWZsP
1a9cIGSox8NNx7P9pfhxe5X37IIFmTaX1XHioHNwLNVJnWtmKVZXOCWuypQJqKrW2hnjhkgk7Kz+
wOMgyxpTN88wk9daOqP+slITBtgNRVa0GPB/Qy5JPTsOA77ePMFEFGTwuOQ0Og8KXBpRCFWRPxTK
k0egb58GOPlp0BkLF90UhDqJ+cut+zcxVB95e4bRGBXJTV73aEsKyTQ2QHCNszzJZ7QMRoga0IlN
h0uKsi+gBrCxe8SMNYTerfhgt/VcDW3UzuN7O73BAXn45EDa+SLJ5vR2Mrb6LTWhG7wZbnTqF7B4
fWvjeXo2DP3/wQaMkNCtCDJReVQqXJoAZS5ewULwl/UP+xo4y2qTk86UcYzW5s91kOTB4BmX57o+
rnkrWi24p6R3AQkk6II9zjmnLPzEGE0BVjBU76HYYLT4M9F+UfNM+GFtdFmM/Ux+oCD3COne1Bav
OdRIIlnHbOIi8Ns5FJL9H7AOwq8TNjCIqG+3LnPv7nH3WGHgkL9sLnmxeoaeJlnW9iuhnbiDB9mt
7RJzQm6e23tr3D3+bNaJPZ8+zZ5lYFVy74WeY0yvarEGjvdzS7ltKqM5Fd2XV5b2MsHolUM1tq1D
L0Mqhkw8MnnpkTlV7N/+7hXVVpzHw/1IVxBQA6MdGq2fCHJoQC1CiOhigYid6wTX6miTTQhz5B47
v0BFMB1gVxSkTgGPrFIHRHVpRD5ZzTlF2TNDsBcItuPGiBlimJ9Yu36ma++f9mHb6gKug7W2fqw+
VEDIfvuDp1l9d18OjFQhO78yfEyVUC1ULLKEeWGoAse1psaAj5tOfPkQmQTC9vJl1NMbaeBgMdBM
IvdnF7BvkyDoIGeVkNvRHrAy6J9PUJHDwariKGwjw1c3gW2BZpxARUppt7uyGUR+IKNnLDBGCuT5
C4sufK7mTBGItiP8/HQy/lthBFaex2EeqPZrzlO5OxTBSk8/r4Ehf/sR8PzbyuADIOS8dT87WF/g
u7z1qrv0OZVZZMcwtWqPfJ5z8a652lWpKorPe9ZV0r1VxiuF0Uqng0J62RN+15TmutWW/zICRGWy
JFojkjxBdSEma5bmj0fknwoTh8LRy+RQDQqkylwE6Ta65OX1kcI3IYBy0hGNvCnnksS1HrOo/rWr
T8+mBNGp1cR1wR1cpmtgZ8M/Q68/vBhDEsBMDDAYYDevaV4/xC/mpi8LZ9l9JA0eM7SXWvR5ghot
hltnV+EDyFit5rIr9ayxrSjFrIuDd+tlbmfAYnvZp8BZeaVSle2cJKqrQ9+WUh9eY6aW/EuYPPZ4
Yw2fshI/ecsFxYJGSSYjDgPSB/eeH5Vx+wDwjCPEG18B5RmK0nrkWbBujKUoueZGJ6O+Sbn8Nuz5
SeP/ssf3vViGotrkwLfHUgZZSSBG042C5Xb/qPUyz1ZQPnTLwJ63IjpMrwx2mHwiVPIYOLu/6zZ7
/aYDV9vFQarGTyE91rnuLaMe3MVWEy3yilvQYGl5xCxWlGZzCYR4JINExsXeoHEVGed8YzCLEgD9
WFq18Zd/a29UKLfH0dLwQDtOZu3+lVRoyjSSSitPrOS4MnUYyrHVXu4msrliTYaA2kC7I84E4RyQ
BrJCKhq8C4pmzSiF9mr/tNyznhDdG6pIdOZo463hfJgL7/Kgn596voRKp31qoXDZjChlOEJAaBFB
gZE4WAHHtJJ7Q7aZsdw8ZKvZnAdjbH5sVmCeTft/KFRKRW68mv+++PEYarS7KA5VzRn+lUh7Gcny
Kd7ttDZ1Zs/LNqwqns4fo7bUkZKIF4XSM64bpwt9n13NK+/HR+RWgWIARFWqDcJIsB7/ywY2ncav
/7yzy52Bq0ufwM4cWm1RG/HNFspMKx8mAfrkB4YcKyn7UWGBg7Yzsk1tT9406Fv4BsFmdKUIhR6X
wkWQs/hizFBJ2wE5aTllKKpFRlydXCDrXaG+I64tQgmwVcJWdeni3i9/5qHItqBYjzQv8XutR/Xf
73qB43ooO+CVoaNlMy00LBXcXfOCVFk0EsvWPYIpKdPewfc1BDnpol4SCd9LXpYrhRqjyYnUOdqN
imvQ0QIH48XZyLiHGazFjk1FPuS/9JEaF2qj3rpRWP6yMJWJewqRkXDqZJIbRbaRTahwp9YS9/Ch
9Z3xw6Wt0taic2TEvSAkqwsYiXYOVu2Vli8Ger+S7fTCaWwUK8gGMnkyzo1NDMY2+hRg/6e5n+oH
n0rQNGz8XOzyohA30T23Ej21XAwzTmHyZckAJR6fDKRCjAp2fJglwWuzrOHHCunNdwFyq+QgEVVi
2OoFNlSGzQ6EQiCa7EYFdhBCdsIEvEcFZ6IV81WOioh6/PI+V7GW4lUxOQiQyWnjHA/0yy//Luj1
JFHXqtmjvPLALc9nhFwV4cwxIOdeKn2eL9BlY7NWL0jxf28QbXPsCoRPZX569P27D0EVz7pZPOTT
tjdrHfMs5IbwpptooAlo1fslQ9v7WCBnJfoJgw8cgHLyUtVcmp+JQir6FyB5zrlqLAi5kAEWg9LO
Gvy3pXv5tS+zLTBOlf4UbVpdp3jHPAgbzrHwVh6bW57VMHAD8gEY9SPvYSr3UsnLFufdhl6ZEHs6
+Hwo9lyN76OjD9XxjDAXWxDbxrJHqREZkjO1VGIFri0LXtHD8d32Nd4fKFr5zaqXBRI/oVQ+++ky
5majiyJh8FADNlhIw7KC738jIwuBUk/hiFHrZ5drpdVgooIe6v+xQxjkCEtDc8myw+fT8LovphIW
JnlzbmybOt99iFgq1MxYs/bJj3WOf3bGMn19eWY6+3gcgLWY8NinXcTvcFmRgYBH2BaFeZHdQISJ
TzPEXcRmYgA9JFIkqJVWhIeiQPaRLeVFED9b1J8EHhFwZRIL2pUOmjPl3u1hdaH3KHisnDY+UKul
AQwys+Y5NlhwhfY9QGWskZ4UsulBcgt2/ypwkW7Whlb9g1btvfZluzn6K0/DN4GTGgssOtv8kzdl
SUAFk6oVQf3k6pLf2FZt0nqMR9h5UGb+iZClSo+b/BOdTRQevgxMPaWHxRkO9gcbZHhW8mRIHzqP
qljBwBtSvna9oxdFNScB+A0ZutA0u4b4DnfAKhtwC4VDUcxXncvhsVQX6eAPdx14Eex3LGwd9NG7
E2S9+4Qd9yt9NgI7VGDdP6zC0VeA2/Ptkoe73GA9dP4K8LfCbDZMYLufHXISwhgdPBdaSSQCXpR1
0TpRRbGoLp9Wwj0DBERKsuiAgetcb56f6sbY8mC8euEPWy9dcjlrjOnYGOBdixCUZ6Wj1tGOL/bV
OTJJY8mTu3G2A8sN9qqvsqecB3Wm/w2j6ddz8JXpHUr4WxLzddwC7kbuFgRemrE5qNv5TDREWrsI
/44JppYsdbujB+AaHavpHy6SSJeZhMEHAOZQNVD14BuBAP7yWDV48zvTsJFXjFmAe3RRmvVw6AQ8
8igFOgTErcqmedN4xVUNpHRosir7bOeiDHps+LEXfA8tfuE3cKAdg+wYvExylIfrHSwHyPrA32n6
kxa4JaJXptii32c7+Mft58nxRsdzgGZzLWb8xIhRab0DqXCEM0a1NbPoOqCZxNdX4/BlML/KImSM
hwubX1MdqyRh8qyrKjRZw79wDsCOJR5CAFe6EBwmCSo4nUXKw2gAI2NNU7gSm1k4Rj/fO+e8I6b+
E0SBEyOHpcUtfjEgb9jWKBY85JoaEKiAjb/28GPukDY7xD5HK/S2gfuwX527oq87RlGmhd0vEn9t
7asLDbysDIuMK+/Fmd0Vy1h0qVxWV4VvVobT0b+HkA1R0KXoiBvMA7D0YBxOGswXy5w/WtcHHDv/
drpmmePTvMDVqXQtdCUnujf9JjdIg/PZs6t0STdUQF4au7BQDsXcMz/AlJUApd9dsFy8Zu2+wJnC
+kNEOkxrdiUhPJFqrsgD9qQJPDtjQYtqdQ3MLZcJU2M9DvwqXEv8/U1Y4P47S0r3EI5d5+r0PNrl
OSzj98CRT/8WBhT0bWbbNmNs3zlGPsXHm2PDdflXOXasKRDV2DiaCWrnmYE2EUBiKkkVO1mFCnlZ
+STN8llK1FIQ6l4y8SBOnlgpu1W79ALAZIgcP8ZrcniCGex7dXrd3xlPvjDKs/9hgmynIic3Tc+F
lRjNw3WGmWYD1tFwodNKt9s5VekVa0J2MAUFDvabJWgoqXs9fmECIN2GKcjrOsYlzPn5AyBBFbKN
dJ5LIeV4+5WfVXg/DxsxgD88aIgH0BzXhmWgq7o4EUkoW3hv2frFhRl6EegII8xkOX6ea/w6atHP
IOmH+9NJtZpgKIKlBFsoU+Tf5KmX65MJYGEaWHwGaB6ZHH7LO4ON6ipqhOUgs9txEURk3QoQX6ba
NwH3sDnUmKYfBAFktFYfj+e0rJplMjofKotRFernSYVM+Q/xZATNUTyuhXxkK7ehJsXXYSyj0x4Y
05hKapFrMXEWAbXkidPS4yWoz1qfkmdh9eq1mURXcxc155fCrcLCuaJ5EGq/QGtgjs41JncY/18g
KxmHK9xpbd8EbNiB5HcVARKbuwTzHZdJTlVMujquD05bAg97Y3Rp+fjenoUSUu4diNonakuk2HsG
OSGCYkScnxgk5dH6q5y1TCuAZuorx/bswXwcVkcytZZAVbFydxhtSIsZr/p7hADwKHGxDAr5q863
JfPwWuXupaWNNnZ2Yowdf41fzsWR2HXtDVIt/h4ao1EChQsgc5lbkPQm318Me4cfA2OjxWUcm5m2
8HP0m5XwUbO/JxRjsz5NczGtFE3pFMSEylQaj7n+kECz+xS19g10MjpSrC6ZbiLHdhFzEAYjCn33
/ulMIyeUpfpe86zJujk/Q8Li0+QZtP/i39/hNUMuXU8gF5Ml4LwqI4rLvjXCzknIR2g5HXjWDvRI
bgZzaGH7fkaDLwatC3RK5Pkn4HdK0HWtGGc77u2cP2jHo/XgYzDFwqD5BvcG1nIBmR9m/4x9Zivs
kCQcgSRVdv2NQuapPdDzxWi6xScedJ8d6FS2k3ECXzs9YRy2S+yDliAhvwMiSMnlLE+5lGaeKZbt
IUDT9OoOmVegIYtV1eVTIWxfUklOJWhGxzZpW1510JhfmIwtdHBr8tGgrCum1OKdyzLeWFRAZrKo
Pwv4eZzQkS9nusL/qY/+Vw5EK8Z+GGn86Ria9rj5F1qbYIqlVA+GlYyHOWiTKKVlzWu8+Gyk4OkE
XHiTshAa1r+CHjV+KnF5zGd9Jt6zI8x6IiBnDX/B9aKw8h3pRkg/BJzp/K+frBKpNZBa5PFc17Ba
AcZw2b6tYrReFdveDNAWMCWRXTKtVpjf0QZZcZ5NzRAPrMJTG//TG9boSJPLACclZh4hLUvVqA3W
1oXeZ01zNSTzPaXtTaUqLl3zj1e0yIeRzDgBqvw4HP/adagFPc4PRNg9ckZcjdn8gQslwYYiynCb
nr6RxhChcrO90Qfi7KzYJE6y/HpE+oL02OU87TukGKGqjrdRUdDf5rPsj3ZPHigCEEU8aDfgkPJd
zlI+29lmdYYvsw+szxLM7pKNg5u5SUUZ2ZgHnDysnzaKQGIOjBe8b0jUs+1RadTn/j5tenOwu0Ll
xyj491qo68/mSkl1igQHw/BRC/o/7DhcGv9pOxHWNyzuDrVOEtVCd9hymgpnshyX18LvS1kVKs4C
W1L0XEQCf/a1T6J2aiqAZCSFkKC/U0D2fTJrMX01okn3BZuu09hc1j7fyID8ynJDKmjCS2Xg2WKb
2tbTlnRC14Q3ixAr2DSpCPjNMWxbA1Nmup38fQU2nPY4ge4Aw11DhUPHWlfcd2eMufhX6nJJqbRn
eKQxITNeP74acE08/xgPATq0ivHDa+AtcgdLpKy6CPj9oewFUwHSOGqXy0qYtHxXLhW8g0CO2VL6
rSe4ZMX6XzuEgLFe6Y44fvvXFXfpYfwWfgrcYW3NAnPhzw7OIxM6fEtZTb49lMZWS1UjkSk5MA2V
zENdN5u15caimipfoQSr5V8Oco+WxLAzF2dBgCaN/94C5o/CXA7NxLBDoLian9F179vMNRePMcfx
9cu5OiVaI328Balkq59+LqlQ9RVv7jmv2nqvMIaZnfm7blGgoVdQjgK3o9zqFqPSx4ue8f5iTD5M
fGQXwP4QC1ARO7gU1qCRa06EIz8f9ErTjNAsKkRtu9wy3DD0HAOHoj6dU2B+CH7bDWNLA3TSQXNo
Gx9eu9Abat/8WhMCa+IcMYvlCfbl0sOs6DMxytSgFd8mULsDkes9U/QVhHNVoSbgsk2Sy7kum/MA
GgPV63cUcDDo8VKH/E0nv8BxmPyTT6MEu7iihOKw/VjNE4p8e2mZIb5QbHcVpm+38jk8N6RpYB9u
ewlWwy4UF/tGSWXhMrHRnkQMM69ZW0O3uej1EI+xTeIhc8GwZX+LidkpfLEEYyN19zlb3g7QtqAH
jnr5uovRujZim1a0VDR8l+zFyxmkVDm/IZJQgYTFhVtNZK73jyMNg1S8dZeUoFmkspMkjEuY72cp
rQ7NX29sfgh2QdP3WytwhpK2iKNA075UJUMk3OD0X1IxJRR6eUT4WjWBtQ6UXqS3Ir1dauP4qMef
8aBl5rU+A++pg0Fj4Y1o6k3cdSKxUPrlEB9u4fMODDfGmHxVEc0FjCqthE5JHJp0Fal+arH/UFBx
qyFaiJ1U0tb6NgcGO8t4WHhB+P2+BJb3/Z6DTezNesGxzKx6WnXSGUeYeXaj+7LWSxujQAHeiFVJ
/X6t1e0NIevWPtqB40Go990U2UagIhjYEIqMcLJtMcrm4Y6uL1iS7vweaFylI6CPL9UuMbIgxj1K
HztebaDVTbNxMOZrbPlYqg4QZI8RnNBrgwewf9I4WhxhsBUcNpJc4Jw2lP8poXDHFfMzM3/RWYXt
E0B8dpg8PaNbRMMLJZ66emhVKpFU/xoORgGe2jIGk7uomM26H6INoBJH2BY0okxNv5BO6CnB9Pbb
ZkXv3atCYeM5596uAS/JvBSaQz0DAEf9zMxlzDJw/cAnXa6VGbeQm5+C4ZZLHyzmcpZckWRLrivP
BtDm3v7Ai1bEvqyyIMPEXylJEcj7JDptiovitLygzDFc5/USMwYk3WbSYl9+bubVEcx21m+qvvxH
ycgpxc3OxjrPwi0fnDx3fYNiE8NnFtMAjHXmoMJ5q3ZNv7b+oH3AdDKi7M7Km4rlR3QY1SnYUrF4
6lQTWOeONRLWFoFtoEN6PQstoddHXwp+rl9ZIyGofT84AgoYb5GlUjzerAT25oiwMmpMgoFVmO5Y
bsvqOXIeDYYkwu0FTkubqQNUBYPAO+yU4lNbRshUMMsb0uvlJdNAy5Z0fc9DoUTujtnR/BuElnX/
jK51rZlz5eyNP/ZiCs5eGVjJ7EaHdoA34CgUGGzBQE9hKr9Vw5b+mpbWnfpHuu9ODjlbwkYgmbdO
BZIGTAjOa5D2SGocgIKS+uVImY0Wd0vtRGiEhFz2/njMc5iBj01uXQ2UvkLS63dvL3oc3amBvc4E
Y+tvsmztjAjSHFnk233BHB37MRQdC85Mzw0NfOeKvZo5px3rBqLaO3PoSm+Gphlq+R/BXnMCWGue
8ws1ixUtH1dsKYX06cG43bnLXGKN89G4hKjISSCezZfnK8bYqHifB6BqZIWgJvr5brrR2etqDnnu
DmqF3w4o1p/O4Gjt89uuIXpmbnIL3ynSsOaAB6NcRXryO/INJVXmJTFEeRZuS4btM5OFDPTEbvbh
AtIT3e6q24lC7esuK3EulL2cHXjUsA+2oYQdEuQOCOhyje6Lej3uiFyE/TtEUygjFvVjooUgxk5w
CNfp9QHOafkHdiMDI4/KgQTiAhs9+TMzcyqWXnn9rkIHeVqVnH7ZQzMjTKrVXTlOomL2zg1dsk/j
XBWf/XpoT3EzMT+cqAVINpcAT3Na/WF2HXkEvFIo2wcuBYC73goBAplCbxkOe+mvFTYAMvXU942Z
SyGU1FwRXqNQnndxFomF5xglgUoenSabg/27DmJSP1ptp7+FYBbCZVuw7zHK+xRygrmvhtMVwUeX
xacaWTWgytK56tj2fMAVSf/05f5Sz3q3o8st/TJtnC3DJuUs2HVrYCYs5cIjpITnZ+ZuypCRvgbE
Lxi/aMRh1xHflj8ND1X/B7OR1E1TXeeiei26hZtmBrl6EPcskckd1Cf4pDWoAoTa9LxRYvFt16mt
A6bx2/S5G8uGSJQhZk3IsrT8hvBCgH8qHru50WQPvPk8B7X9V5Z2ytnQ/2GDVRfNAoA03gFUH37u
BLZUlQcAfBrVVrLeOQoyhCWuFF642jet4yh5gWB80dGR2WpiTzEFUdoaqEQrHoMDf5auhtB/qDNR
N8fPSZvmE9w8hh+xnYHkQz058UeRs+OsW/CtwZkWp2TfVeGcTE1mhMIsZtHVPGAlMvYNiml9Y/e+
1UbwrUs24VzdilyfAdr1ur6f2ypyRp1KkNSgXfbVFZwwu4+JA5fd+hK0dy0PraOC7W7Iyp+NZDl5
Bb+ef2IT/hdZ9JdY5ZYToYctEhCXYYjkHkAz7B4Hjo2KkNG7PKbxXEgCtEoPrP5IPDiipYdwiHdN
1pMtriqPF63oatdiW4uYk8MRsy9I/jF6y47/KIBZqHh1XFFF0clj0JmVGgE27BeEE39sicHlCJhq
26YpVpOLWVy1KjUJrNkICLBdXcXJJkGZszJ2QDL2JMamEK46PQJDf1shgHcEGlV2ZBXdt99JKSuO
ml1aVKI312nYOPIdoyOYozNv1lBfrc3wYD6rER7YQnYTWKfP/8qR487EU+TF5O4Mwsn/bFqdZmBK
dFeUJPz/sa7ar957RjXs13tAf352ENiIloN3TWI1Bex8KHJgvlJTWXpvbkVfYXYGTnEIXInmsQcL
5vkV3THHNbR6/d+IIshNdQHB0UntE8irLwySzmodtHCYsEIDZwbv8obTBcyhVk5pS8r6s8gn2lr6
JOTahflo/okuQ28SjfufFICUr7300BzbhmLhhPQPgppo4483AB3Ur91ZTTDr5uF/tMQ4lD+B8XFQ
Ojg2EH3O5aXC+D8ohT6C+8EEgglbgRwdtIA+UW2rtTrbaI4+CmpPCODDiCyj4k9LG4KS/BNZzlPY
KJjzAtvqEP/xYKQbDcWaSuhmMTwCfXOB8tOdlKUozVxLZH+3Y9OPbgXkyM8ZRquXehQ6qrGSHWbb
2npl5+Nl0sTZ7ClWjKxAXdHOLAhjl5WDeldlFaOcu5sHmV0Lu+JXq+c5sdUMPNMM4hrWbazOky8J
qUmZH4BQLk8ht29g/FgF33ABLIrwZnmChN8XgkVew42/FhViEMIbr8mvTnlh8SXJ3fD0fe6i36Xu
AFqzk9PGF+OTOdfMO8k0N6G46uwgXhKyQRMbYWIOOfLVKw+fqcICG8x6A94dgpDZMCMGOly3qsBh
Y7B8ZqXMn71Nmlg0Hs+l5Edvqtf9CI7K7gN4ZXxbWEtHWPXtVX3F3s63kbvoAnY3xBmFwJlggEBe
cYGW4fUuJiJcDPJD9SWTTOhYTpUQAhRMi5jOKTWjgCYOaRWZ7xhqmS4Di/9r/as2VlW0aEDNeAK7
xwC6nPqLAqoROWxc7c09xgSbM2JBMhSyfux2wxWJkZQaMIa9a1qe6qVEdS75oc7Vp4kD+KTG6Ynw
zpokP6ZSHOV/ZBivt8jzzn2NhJWrOr7MZOgPFjo24tODIF5BkFTFW1ErZSK4TDN+cUzqMVw7UCkm
r4NkjZdRtVOuGT856/wBCFvyubxhqHlW4RTayI3LqJp6DlHGp0uc1YctqVvmbZZPew2gFxQr+2cY
ckc5JHRR3fzegixQiNQXF/vBzo3TclIs13fer5WR1QVPIVtLF3SLzCY7tyCPYKWZE9vvxytZxq8W
rlXSCXhxw3dyWh1lNgWkj+VxUxYj+6q4bEC/JxQGMEbrHLu2TuYh30xn3tT6R7tkgcaFtfK75Pjo
fleG1BVIQkJrxsVrUn8kIOJVgomLe/dgIA5GKsikqwHCbBdYDst1yuUH1MeEdeRviS6WDP3pEeqI
ofUbj9V+X5fvf9yIU1B4gEyeTPzzLjZTtxNRVrz7Fv78htPVBlMOsfOVAdc2vyn9k21tywhTIRtv
TZN0EyefKRwrAShH+HWGylu18gN3tLsmDcwcbG39yFFsZz8iUTdRtkNATOMxyakQtduFmsfy5vJV
zsKXRx8SmS7UKSVuK89vGSBoKLvibqHY2huhv+1udqPs57y9XNiq1UjvTrs6//Jd3z64SUSJOgpS
XQeBdtTuPbKL7np0PdI4jOrtP7d3eT1DkpShBwuDM9MchzSjZ6WgzWnkg6DeUQ9CsXZt+k439lu6
oxO4O8WU//5Ngx6AQv2Pvf8lduhpuNbja9QqDeYUx88dipBarq3ru0P5dQGPnl3YcFjXo0tns4cT
DhdDfYqeMOeqSar3XL2/iEv6xJyJKcAHaa3DcsiWqlKRuVU2+f5Mv/S3iLE6irD+azWlyXrmmP72
6povRaf8MdK5pyeAypb9aaQ9GSKWw6dlSkI4RW43RtWSFseNBmV+obaMOwYKThSpak6eXw0uI7yy
SWNUQfzF1hbCV6Bg03C8g4KbYn4qMshc6H4unJrOEJCC+ZZeiHsgfrpHFVCxwAfipuDzmht0+eMt
FO4LrTFm0ahFT38aXa+0d7SbrGcm71DDXsEAoEt1tMG7N23yGhls9bvwnO49YU1GS1rYObvEGihV
D0VGB3PV8lFUp/j8f9oOqQTwEPWkZOdPXf0VL+5neb/PMqmhEIzxG8yx901rpVxKi0akyPMvAIPw
8rOLSkHWglkLi5/ybNrYzLNSiCFDlXZ3RwsL+UHlmQXx9fJ2RY167fcXIhRRY68e/m9FiBtwRqc2
hcmZDUAzYTrXfz2s9jIoDLneD0QCYYgB7Du9d/6o3XDhIOh2CkfIQ5ECOUdQFDtlQlQaX8x8RcDB
d/YXAvAJxy5bvfHFJD7Ce+zxwQjsDgJHJxX/FkjeTffLFwWO1LJ7AJro9jJSuDBJUTM6Y+HhagE9
N3V91BpTPF593d5ZiC09xaMW9QsBee+Y7V/CEg00OU+Nje05Zzr0vt7FpsoQM9PjboEO2WfL/k6s
5gFNvbZZP37mY9VgHsFQGwSBiF3NeHouqRcNnT/KJn2Y1G8nlZuecD2Pg1smG9of/jpfFIXK14oX
9S1HtPsvCXHt9uHHw5mzMaV6K5083FL6KomNq12mXXIqliwIrcwooDNuU22bkUjGCLVSppnHoGLQ
COzdQDUW1z9AlTMJ3W47xHKzUcQ6e7vWek6JzeZzO65Xo8GhBY2A0oxH/6CdICgeDmyEu0EhlbN6
2uWjwK73gSHgdNORbhjqWQ8km6Om93qOqRBkSj/kwwv5WPA0/jZI1wqWCeJ7eF/IxQ/aFq5I0WJz
ELLRu9SBTlvKIGYP0KlXxCsl6JEiEeTqknQ2hrFu1RXZmRIH1h2CN8nF2hedM/uKDTd0ajfkAm9z
jKzZXk7j6KAG1bTnwWJQ/qWTZmTnMRTF8tgi3zp3DukNfxbt64A8GTwmfHlJa3zVOoSxVoDiJC4W
yCVIHcpeQECjO74rexYGao/sNYgIi+RpWKwhLXNyZj7Di0VLH56SPQ5tvxDu60P/GAbIXBFFHvT5
4q0q+Lvi3antoukZH1YLokXMRVOIcP8CMdMfOAZa051BWJNmyWRc8HXXz+dnfnBFBL75C3QNt0V/
d+FduLavpVr2sTpIXOrGYDYs4axbkD1j8AtpNu/swyjkLMrtsXVQyjs3yt5h/0iFPAwKUtsQ0S/u
xP96jhgT5tdb8KSadkc1NIU5YAnh47b4/CZKQJY9kTDdhxZhrIwzEE3xGtuLHdmSTB0Mp25YpA8n
DP8JU78/CX2i07xCXJkSKhcNGUGDWmd69qEVt2qO575J5F7LCuxI2WvaqJ28oC8nOZzLfg6ccJ1z
KoILGqNwOa1l0+j6xSwqrGV5MxJnw+u3l8wRby/FMynNexkGAyj0YGG6j7RPyFn1vRTbMGA6/DN5
1INMH0ODnoZqIILpWQzDc1A/jUI35ofCxu/iNxZk8FMlVl0bZS1Ov/t5QHISENUSHM7mEUzvGOaR
ck+3EGcP7QJajmQZf9BV/qV4JbwlJ6bOFX/yhhn4aHza/X7Jp1uzYL3eLHL6W8fX1KUcWij297Ny
RvYnTsXxDo0sDwUU2IhvLnmFRaXkZQalBqy2ToecPRiDuEYsaaviUeBMvie1Qop4uBHdvo+8Spc1
otGaG/paqFBXC/una1FPbrPFShUW/2DmSjX8cPqpN0s0TivqKuxl9SdNgxH81neIuKFsdAUx0Iv9
SjJ4kjmWh4sFyh0p+ct8SQ6Lgp5Yd6nme0rgTwl9Oe4OptSEWVPIcYzOjtACJE81cTm8TlZJW9Ng
EtDgha87WeMk8fufksEkwMg80ajpI6QOks1o7Y8iA4+TiUQed/ZzjvqtDyBgfX97SLp0hhvmfZMJ
B90i/N+iqZU85stHstHaWKZ0j0C2P2eIk1f/RTGu9WwneBlYRtZN5ohBwmGWXWQu2NrTBmvVaoMr
koNlUeGanfj7UV/vczRR+/xOySXzDlKVs09piIPYFyCglHmKTePy+y+18qvQNX3TsXOtKOXZMkvo
XLj5OO43DagzrvxSB/lLY589W+3s03lnWux1+PCC9rKoNigVWZpV+CZ7e5FXZbXVcJU+6q9I5H+i
Kx5ms0LzLsR6CwdYqDzXF9MuYbneSDot5L6j+Cp21jFF6hI6Jw7sKfdZgKbXmNdgzWmjnNSD8wj4
G4KdHRMxHPY8whhBvN4S8aWA6JKHSSeaznrq8Gr9n5lWjJ2M3Ett+7E8/QeYOIGYhGqlu83KGMrb
+Tec4pC0o+u53dME4ZYYauTY5OIMynyEgvoZ1ZA8pB2TjbWLdkbjp+ctaQWv+FN9FPstSQ2MGF5/
JbjYXIq6+jHojAKoT9TvMEumaIe5rjH276dO2eErVdpvv1kdAdVkF/Cy6iQSaFIkNQXNmTjqjPNT
gbzITbhcgZjvG2vF1Nz598PJgSY/CjdiQjRD5PvJczBawlhvKFVvsfPdG3iC13MOQf8SjElFzJ4a
t/w6t0HvtfMeL/OezWmY51gUb8ZsoFtdajvP18mYjon4wT1COLMnfcoeIN0u5Oq/hdajJKQ3p6hA
mQaKuN8zGf7/fGU+9nub3vhYt5LpbfTr6GekkRQUJNDGQmlYJq8sxX4U16pBHkyB+ju0wvG/u+Y0
D1tF0iT2efaucom9Mjs+8ELLL6VpM72B1gtQfS138hVIuoTYlECdGB5Pw5bUSdapd/OCQ7fVJYVh
BOhad8liLkgucLoKpuOt++6gLyx2whJzwsn/N2hvsQ2TeOrkGHqckXPCu/WMfmUWJW+rLTiljtdM
dYnU/tOk8w0xFuI37O4OMIz3GSAnpcRI5gyTX6AWFNIMQWISi05V5rrFxqtfXbCkgvL1RLTpipDR
QP0dzCMYqh8etCL7WkT8OlOIAgzEWsPNhf7Iq+kYkJF2v8Wp6re2eoDF23ntT1a9FhfY5GEUgJ89
UjKpO3LoXXVj3WeM3e0t43LhXohlYslD3wbnzK6vX2rtsw9YoxJlZbGp27dHdPqe078Iy3/8ogge
g3YuNILiu8KyWmx6++2QdkI7J/tT5Uz6eehtX9zoqjRAsoKtcIm67U8EIVz69gpVHi+dBtEpPLOS
A2tVpzqycTZJ6vdRHifh7q6QsWh5WUFc6pA9+t3tZyGkiI5Vz2yK/Oh0/aPcXzOgbnqCIEKsCJws
wtQZ5zCdNbipSMOSJWPOpNgFqP2SE40+A/eXuzxTGxldElO/YDEj04INOukm7hQcn8pGNMri3paQ
Nw9u2J6+UpgpIOJlLBASjacFW7rWJ4hm3E9ho8N7BwtaGTkx5xqaWo8uHMxTMmV2Iq9OWoFCPcoC
FUHDZAzQRwl3PMJNQsIlPm/KCCGcHQhvgEfR97ye10gkSs5npuMYEnKpCMjwWkJEu03Wl2+n9L+l
mBv+MMBbJ6Tp+z+qhqHz4QjPui7Ov0ELE4rwRH0mDk7Kf2C/qj8DyOYw19rjQ7YxXSBbdMtamy9m
NjEZA1l+itWoezDjuHJxObOC7M7RfVYHbmXeCt5QOvs9cjwGVnyygoCIMKr2YE+PeKr62G+ExwFb
3utvSd6zKj4U7b4K3q8Rod8GrDsy/zR5lZo5Hnu6HQq78xPRkgecAWwLhxsSPGrUuze5HvY1mP2e
xDdos6lj+OU+c+b9L2Qf1EUk2bNKka6xHUbqH4d1ATIozyYYbK9fDJJ87GZhonJrcSh9yaiyh9Cd
+LThP1KlXFtFXRAtqbra+UpQ8t5ykhbw2vLBSsJX5tXVIk+NIopcaPvQDR9bYeqwurMYEkUmc8Iv
1r+18lk0aTayq3VRzHdHWlEWO3vd0R1mZib10FUERMC/OPbfEcAZjmpY0ZYLkA8na8yoVKovUFqA
hdJtFCA9HarB4rDPiDg34bREKmck34T3JQsFsZqRXptx2Xp51PlOnzoZ+ZTQeYlB7cF03HQWmiC+
xmvyFQ8/LX8YlAAtALHHqLbmqCoyriOZTmTX5kbGWMDkPDimpJIrbNPihFFZEKSZOF49qfLfkPtf
BJ7ngCC9Nj1IJfmJ4UIFLlU1LuoqzJ5ZPx5k4hgBlkbLjTQ/gc8gs/mZJ5Cdf+ukJ5tIdW1jqx/7
WThl4eLzUyt7w/HS4ad/TSkkxTXYRKLhrUMZb/l/6XGsOC5+Eo6lLDJj6hwddf0cPEpIzzzNPbCv
5e8u5ReMIIj6l5AUTN+EZrwQUNv1IlPb1oNqUT3UuJHFi72LVuymCXhK25rk1T4rr6My9gek+td6
LAgzyZ47hbH5ZOMP/aB5H7DCRK37juj5KeARBXXQ7keeoQTCnZt4X7hy7gKyijVyDn8MEZhGce3O
bT61dW2H74qdgQ/rR7w/ZunkWLT6qw2V/DsyrTAqrXzNv6PoiMOMybhtHsRqaqWBoDwNxP1EBSd1
cCElDMoY9HudXhS0gD4F+bdF0CgeLJ2NHT5XbNkv1lvn7KsLMyBTkMkXIc5IR3xkKWXQCiIRqrJD
zs718Sts4rntuXROCt1d9B5IOqZtBMaRw//+FkcV5RApbKxyDU+wjIgkoEBhPUuUp2KBhApjrJaT
V8j8EVX5iHXATmbtbAMn3deEbMRglTLwLNAh/GOr3fgK2AaPZfWhhg33GZtDKZqFlN8QT06kFo0q
WXVinli8vEnkcgLYzNlq9RSu7bUUyVQLadttGxxZ6rwewd/O+67CcDA8rQHzpuCMrDA02DtygcqB
mlDySC5YotTQrtNSfFrgsk+ZxR2U+/T7MVjTG0tVtJj9lPWpvlgfitjT5SsVv7RvLf77oh8ef/n1
N6KTAH0OXrVNlkppHR/17i/7EJXU+O/nQgY6haVavI3fC/bE4fet9FJgsC4YvtC82pkCQTDAundX
WxVBieuPrN/zBHxrrDil5WRSDXR/JyA5tnbTaokuKJOtT9XKFFVa3oM+YXPYv89vdOxPSquzWDQc
a8OJYl7P5nJvumFOd1b/X0KsT4q24r233K8gNuhIH6M45UzxcZQLLrnUsR9iTSGJ6VdMMwgy6MlK
OghGGHy9qGZNOqKFAJmi3+Sy1DbjCIq4QREkcTm34LhiA2h3akiPNKDMSuT1l4JHzXsiM6DoGiFF
fGqVE0uE3B9UpGK9gEgjJHRZSuZaljitEMqOYekrNPUs3UxYNCxVLC48KZqG5twvN6YaUixmSCmN
04O6tv1XSYkOFmzmLPAq9GnWy49tPWRBh7+DQDJDdLmJnP0u/Df8zq5RywcWUsyC/vwPVixLaiLV
Kn6eO7k0DIVQZqxtUFlbLfWK6ZldWSldUL1b3EfpPYK6aKsq2ZlWJv7gQVJCbcjBM3qGSQUnD/cp
97fWkrCVIDKqyLn+LDIjr3YErYCkcGdpB0TVFU7zRuKxEj3GDeAiHRpOjzdyk+zX8IcPDCkulM+D
ycy7I43hBkEsRWM3z4K42kOg8cs2GlKgvlSz5D4pGEP9cFXk0gsW0NAn/mH6h6BUGUw+zpmlftiT
QR5+dVhDgyn2haY9Nl9PLDBVVv3JNExNDspJjXqdOO3fH9T71IhJk2PuxG/ya4H9YHPBticQ9Rjx
vMRsmY8ePNf77NIyVKtD7PNuw7API4pn7SeUgfh5Lg/zVJtv3JDHoDREMXOo9hUM7Yax/yi/2WIl
evHCtg+LQk3F2fJM9z3bfQ1TlOYZT/CHLHURHgYtxsUIDP7xOCO5YeZlCCYSeDoFS05DZwOPnK5z
HEnWlMB7HHwwtn42UDP5kfHpx08FyHgbxX86AGm1HzuPoj/Y+OoYXBS9XC2n5QUSjqkHtq2li7ob
NiIHke6PMFtLKPNKoo4MDRQfq+so0e+fecmcOAKEtfj5lkwAV6AHiqeKewOQXEqOXC7If6ZcDBTX
Osv3Df8at2sh9DKe6xL/2cDEKBKNbtIixwpRYDmbcw66yQfwUCzIkfQQDuRppwkq6DxUjDvF8EV1
3BGLsIq0TcWEGC9x5VtV+g7k0jLwM+z/zYZPH//+yelqUweBrz3cWmmzvvL9l/VoVOfIunjspYfD
mLwuOcmmOUzS0mmfhhFRWL713GwMslvfps9BAJeCuGJUAtimXtpLonu92ctCKzpkb0Jb6fDYkzhu
qS3SbMD49fPACWYrVCI70sEkw6umSknGBRaGZ36fiRONwf4NyCM+xaGk0vxTzAGJJZay9JqNqs5i
enFhItU5uaSTYS85UQkkx7UzHXTPQLdiquoUo06FSS5700ITlZTtfv4w+R4aAgn1CAwTuqEVO3iC
Tqzb7FlSuLeN5nx73q2cdb+yQFq/tsyNnE7z333HvXMaDV4tCMm+TsvXOu6X2RbYVk99PILdJ27D
zxGXD6f+6fWtpeaMLc+MKoh84cp6nEfOGfebBlgNdTrcn5OaoARB2OuViMQ9zoQViw5KeMN44EvL
2zPX8A4/H7SnLWL/hbZogoElHpc09JagmRhCbu9vOvC0hse4ppKXAdarzVK0u7ufwxw2KIhJKRLR
T2B1SKXOk95rAoig3jQU89ARi90rbjOfNjflxCqLGr1by7Oqp9Gm47M4fcjQbLqV7GviYcAl1vKu
Ro8bBDxtcfz22bAX91Is0n9dQiPSAkY6z9LYWjpwgGYjYXjDdGVGfm2v0TIckzOfhDbyYNDtkZgc
7FYImHWn55Wd5BsKelsBPHGKEUOLKrQj5CAmUlz1dGfe8PhZVhBR/K5I1fs0DmF477n4Zdn+JrOb
8IpRfMi+uLpHyiYKbDG92wcBTKHZYhwU29aajCfPk/3bsi1u6Q2ZvKq4RYhn7PvUs15yz0ktpkkr
oRun0GlpzFmyOa+rIyInpQ3XvamjdsISHtkCRlm/Deo2ZYKseMm+9IXuCiGaibnQd27pkYrAPcI+
vOQDpkKer622qR2yskm5jqcn5ySD83IhVO1T+AhqMKdGkppsmsjx/jhjypRSJXPKXUn6gUxyTnyW
vM5OeXI6/EHcyJvMNQn+Dqf4FGi/V4NOPpkFEp76hIFFpo8AkznHb6fr3Co0zQe7hR+/W9ZQOyID
jeUh/M0jT99AX+SxgUtvbf5W90Yfg8me86Dj1q605GHRFeeo3lKigjKO1gUUXz20ydoqMoB05J1j
YVR6tk5xQ1OgmOJ8zvJxvneWAIbgPgf9lyl9jFdwFEbCyNDgcQPTrU3LAlLHlH+IUNjTqPCqfR/n
gzhQNdY0stlL1BmnvpFTNbx8XMuhRm/9WBVYMEYoXzNNDImCR+5XFbFL2AEIqmXk2+1k2940Wmif
XUOjemYMzv9DbdWGb+w5J1Cw3s33IH2Qe8UHBMyyi4rBjoJ6s1avDOL20p6doRTJeRnrU5e8dNSs
CuMk1fJnqk/9k08/gmUr5gVyL8pQin7exNU6Mf/oj6Ep1o+Dv8s1ZIPjWBjVwI90aKjfZQHRHZE4
oUEzZJNU2j6bIEWWIobnuhwo2kKMsNSYLnt2IDbfErMdA50CHWtiqN21nnzO/NW4bu86+UsI9yFh
qSzwTvpqPSTwDhXnu/R2Jnt54XHX20b34f95+tkmPGMvpsZr2OrBb86HLk0fgQu5LrHkY1zcR4l3
SKQoJlfcTN0IEwb0laV7NGE7VDev4h+r3rM2UCE3mxboFHk+pylETWFTmQASby41Rtvt3WG7V3Ia
EKEjNf2jX7JoxPzMUuwU6INpvOt2WwY2hvkfXPganEkUOkFldy2KJ6klPR+08otDS8MvCcOoSeaE
esOmEUJ6lYXewWQT8TWJeFJR3UVo2mbj3NSd/P6k3UAlVzJS7JL5cS2Ej37Y9TqqHyE76/nte7u4
0MmklT/5fxGkHHDm32JcE1kWkuFQpgRW0pqBD2z991SqIrpnQxS4RZwtFT23shy9Rhi0V+eCRwH7
zMsJ+N5yHd3RzlifVwarsROFTFOr+DRbDCZCRTY+lMvcwOB9gfblyB4p3cVySC8jFARk29QG1dcT
O+hAYMdKxaZjvqwkAzVc6wedHkVySoSy+aznFhQSUZklzTkdykkETwHVmom42KOXrD4odfiCdGgo
932XtyMstYRN7JvKzhqTRjYDZx9mxlw55Q9V5tIMhhuJ3j9o8J0snOZ9R1k3MeSReugnSCCU+4lj
NQzLt/CPIkgjmxkvFWB20YKBDDvaTqw7fsxCm/Tl7SJ3d5G/uTc03/zylz9nFRV+cr5zqzfW75qT
bv5NRZEgocwhflRNwDXQLd2MRwj4W3u0pf18g5IXdlmsOVGiuCAa6QBybKlJpPNjsqMhEk6g1hCN
b/0UUFYqwdRbluWAV4G2XoOX1uoPC3cZCUfdNwsjZAO0HpWYzmdxmXlkVkSXqfK9SaS031mYcRbL
6qOSIdAy28k5Ba7Z3q2B1gWHuHqS0FJvzMy6GdoMbj1QnXoyRDf7Y+ablh7xWfbyKeobat/pljK7
ItwpGUhjXtdSxNiNmNXIiFRHZwvjGJ7wWOEkK/KqFXLl6ZsdFmT4dUSuaOPhZ3zav04IS93QiEsa
+178PSmNwlsCt2Tx4Kew6l08I86zAB8XXQAXXPl3D+w7UfpG4jj0N8HSb/1Ckd7vYYcphskSoCXG
rt8e2oIG9/di6eNxnty5lTj12wZF59wOMIQD8ET7N3mYWYUiuISBft6iCcpqcQSNp2UvygXt621h
oGKr85SNyfT1w7oI1LxuVPjgT/5sBXL8TmGoqhkpKvSGXAKKdkYTR5U0vXRh+PoH9O8JzLroQOEj
w7bw5vWoJevnvlguu/7hXilH/8VTqjpmykTXw0Y5NKc4nwVBrVtBPxQi3dk3qZDd3GFo8i7z0gwx
5Vc9XrjJ35yKQ/m+1k8RSysf8xBVFQoskckWZssRYVWo4KFQitIlDeA7wwcgpWAYvX+93feI+azL
dF14vH4fGzH0o54IKurfMMv35jfY0fYJeIxEfcsQ2S13oXrD440bkShCAJ9pLKa6Hii0CYiKcev3
v3CwnEwvsIApiiFULhC2aLc4bHln9CFdtPcSghfUe3YDtObiJ1aF3lscVVi6f7mJvxFSyYdlFat8
hugcBBKB3Jyqj3N0bOrDYtmwcJcsreW/+ZSziLH3nQOjPKVQcA+z3xBFBx6EndouDHdepA6sfb3O
mgW2Vg4jJJ6PLLo6+U/nfTLQ1SrTfu8sA6o5ByoMQmM+d+jVTnW86g/7ooKiFdyIgbImPPOFC3ZT
SGws8xtcL4E2/UsJX+oRFZnWlu1ioP/8DhBFmAVKtOPoJta/7ICLnhoPFxu8xZSxay1X1tNdpQ8Z
G/Yyu7KhFLhqMGnRRS/bKGJL6ESRKzGJLL9Yx8wKy7ZdSzrGhgRB3xw+32veOw762OgMe+asGljM
7PowQZsy3tLvWzRhpeejzGu6ZhPib+x0+HSYnOfSmLaBk5/7Xah7gy1XYk383CAMQCD8HyAcQBaR
h8ihyEzuGpCoTmSD1GIBwuMs4WWYkwW0kpjEvhDapnImw3ZjPlcKHlo5pdp9CAiR9faQvuM0ih0c
LKChGDS5CxnsEnH4SqiFLRmo6k0scEKtXCg8iVc9ljQSEJ09HitnGavF9i/1qpvtqp/9pLqWy9Ps
KRrAXXnRsSPTQbuVFsVcfWEZOvGl7bI2O+YrqJ2sFA1TacUYILNWBtnxpitZQ6waBb2u72bmIYZR
YSwGth8RG2ao0EHV50kVY1lFbzAcid9zDPbilRXJU21LXmbJ8F5f9G50mSDXJR7E1u6/wBE8RGCM
9tOkNE0BCJ6mJNcUoU1mEfyaVRBPL+9XnCtiNIhtvKKidPyTSSXkZbmS5LOWy45QE9oQVJS/f4Wz
NJkk9ZrRgdHIpwVY9SD/eAyZgmRlEr/ugw1TTMH/6afH5ItRzA2yCPaqad2X+WdloWDoL+mWfOgL
U/ugHYUFOr1l3yZudJFKDi4sY3bAl8GrV2yBAgxXZUwyvbYFZ+s5LB0wS6aoD4abMLr11YtBH3PI
le4cDX+AjbO3bn/hOxxtM3Zk0ebIsD+3cGkB4dGHDU2iODsyR3DegZCV3giANSU00RyOQIthc+7q
PsYQzz/kRpM0cheR3sqHmmk7M47FowuRgtZ82U4qYBYpylmGoEHehLN47LDsPtZU19yyi03OT8q7
ZXw+bc+hSx+RUKIdcjV4l94KvmcLksh6moi7JNOuHvy1Ha7vscS0E2IC2AN9YYWbK4TORj/hsFY7
lsiRNy/4Iej3SFPL2LrBBQ1H2UPq3jNgDuNQUJ77moPreXKKjUn023xRoQ09TalSEAiHjD4Ic+f2
Qi7aZO1zVx+vuRIwUmKRVPLs3hKZFTw9r4QsXPfGzGlLMddtHEIusypCJsgmFC1cQfjtQsRDC1i2
PExdyLZy7PqlcYFfv9MBKl0GnMjOd7kzRp32fTYUvpxJwnnCIWblzPUc9Sq51fXqfSCCoJGrzI62
swjb4/6IBPp8hR5XPqfVohIHvHvVXvbRvyBCxpTOankKCKVA1zfZEm3IiMdf0FAqS1dy8LrPrO4K
W0AozUNV+qSEkK0dxIrHCDWDMEGWwKm143ee7LrJ2tjgCQUM8FCkZHgXBXxiUd4kmlHa+EFcgxnU
gPUa6ww0PWGqlG4Jwn8jiXkn1JBxKgev18f5Pg3g5Ua/fsgJO88y4EHoYHhd26qPyeXC/DP4IAOI
o9pBVWdCRim1MrU1SmY6rzRCkfe4fw5dQbg/hQbxDM032223puNpYbsN46aSqWPo2jXJ9VAZpic3
VmUTPYEkiVPzi6XSAIf+4xELXnqEQJCkEe36TJ/rbG6uYzfg4sM0g8l8Le6YGRcKldWelI/+KXci
WSnRRJ+MhT7vUGgZDEz/SoT4ZBBSVKTK1xYcqyhsW8tSXantgFRGG/+6ZmD8NHPBXvxKKAhKcsjD
7+LcRBXA273Lze2yyGALCOEhTr+zZC1Jer6fa5hYL3HcmO8Absvnc1IEDzR+GsDncWuK8bVAOv7K
0/CdkDEHmdwC23mKLH5oKNyXJK0LCfvdWyvMjEBLcq1uliSEO9zgC0RwxkUt1JE0qWfpgLeyZ/21
ypkCay2KXZe6VP72sYA4b0NYXEIab4KWmpIfVZAsf/xrZwNpopoZ0YCULswgGDLMU09fMCs6rb3p
sPf57+xLW1V9YsJRm0I8YmrD+i7fA83xRR7+mYTNiAWt2tEfS2SE3PwM5oCH38OoilbrsQLbp6Ac
stnAv9e7OfxNYifJo/TsxQADIiM8iJilAl4uPFdi5I3o3164q/U90T/bbw1vfuydzfmD2+SGarzc
HJSc0IC/ieUdoJwHRXU49DrXcQREu0rk5zD3goKuEbydmq8H6Pc1hJ4DSjMWioUYFatVGr0cdt1n
OmE24njit5W/jKaSpthyBjRrdwgKaaJwwiHntGEdi43EbTlvlximngeSp9WYQ7PwjpYW0SBjPGXl
Qrv3r/xD9aC79xEvnx331uG8kRUpOQxmDdVP+KY2FQynTnKlsi2rW5vHkSJEaMweCVlyjXKDzwRK
WlD6RkXunufTms7QwDvG4HHn4DlNs0J1QOp+fnsiUy0FZ7BQqhta7sid3/gfKoEr+VjSfbRDlpB+
MU8YFrN0VgCXov4ZwF45wjsUlHlbJsQoWWSz6M9vTHQUWBuICJIcYn6kspQlB8kNDquwB1xMypYF
yeIj5aHo8QcQm8u8yFsfAYjgkclf/n9bxlcScYDmEKaozS4YevEvGmcxg3pLaOhCGDvaEf/lj4Db
itK4X45EJGpCRZBu5czHDQjHXhiI8eh6YdfIFTqCSSTXGy95gvMoKFZ0ZFOmKTJSoSWEtUBsXDUt
K1mtaefelqaLxrcLAsHOJw+gUHTn5x8n3cQ7vi8LJOIRlVp5ID2Xl4covIOLioU9AnazFHwI/3wh
cUuCSQdpBao3pWGFrCCwyY4J9/meUmML60RaqNyDaZUoacjkco3/oAh1dvP2dYXnOx1/1POJPnf8
GHzAEwTxH7kVUgq65NJR4A3eAbWADU4ZKk5oPXIKtXIdS+SU35r9Z8X+QPrSKKlAw3rThQqytZbs
eoTlwQijhxQrhlsXs5g6ibXuIvVKWFhjVv8m3fXMw/uMGSp3Tg5d+8Dbe9UBdMuffycqw1ic/4ss
SshHe2i5wu0F8PL/OmlZ2Re7uVIP9p6//MI6DnZonjLajVqzvScOtqxz+DPM/zMElnOPrFJkpH0n
MLEYdwQ7UlwWn1Xs9ovIEuHvg4uLW7tNhsKblOPzTJNR9uL+Q8ETn51X5V9+ztk1wWOHxzXDA08I
dIqzGfx67A/Wmn9YeaN7uJqoj1pmS5AH19HyzQqg9NkvqnHXrMQXrniiS7NpiTEvvj9TpSfJB9jP
6ddwM5Z6WWhckkxz7yPED2V4XC3ExCBmq9jvFW3TcbKA/nCM42bN9VSviRV2BoD6aOBigMHS+yxW
4G4viDHRFlhIGA14JP43QMGMBkgF1fsvagtL4/zf7ljhYgG3rWM9vvvqorVRg0DiNVQ5FtVD4PFB
AoPuzmTl/NvS6408Y80cKx4erf+mRH8nUIWAnDsToNh57V/NUjxKT9TzKcVyPn54EAhX7HTh7Hpn
oDCbQt4hgvJpQI9UY7F0vssfOMGJNNaAb9ufAy0unlhzWxSqg23VBf6UGem/RYiNR9Y3DC0lk//x
LOS/tpNW6+Z5rLBDAa/ju3/FSuhBrOPnbAwgd48tp513uzRRMzLUNytu0nMD88NncyAe8XSL+62k
A54DY2PQU25XTz2Aso3u/QjUJXoIWd975ge2RjYiFYCVwj8bGqedrcbCo/lQW3TxVDrmRNQEm3lB
7kZg8CdCQ0EXI1HU1d/W/aiAdEuBDegCQd0YbTWeXIHioh8VwIBwl4lwTasrLE/1j9OIEIPXwwEa
TqaYmB9FrprlsVy1wmLhrCC8v3Q6szjkHoUG7MEl7Z/wfOqxxZe2ZHwSzpQu1Srs2i43///PYlHD
gB+ivZ3svn3Cm4jKhu9CzQ/QfMTANZxI+Fk4FilBtFEXj9UFLdDltYRQrn6P3YTVhwNVigI9DNlv
Au0+2ZlyiYR1N+WfLkOIzvJuTxJGOiNVd1ROaXLbDbU3doqeLrp+M71AK7KK/oKjHlDCbTOo2kZ7
BEAOkz/VgkQ5dg/v8Cj1ps1sGVT4zxCaRpsoddE4Fxzoxaw+njfmsmLvY3WJuN4Fve6YAu3D/6xt
iuDB/hcmUVc/6gcr+3PpoDNsfbvots267T4D2NEF7tw39rjcjCeZ32CHrATnlSbHt9Sxs+lwKQMA
7pdoeFER3O1qsXGIANRE6a+TU4c6jxBeJBCjvJ7tQ3mWSpZYCTL10CzGyxyX1ye7foo3wcBpUSdf
mTaO8YX3H8+RKIG0PGhPAEpQ/KSsM1Djcaz/kL+u+iOsYGniPJ1YnL5jygI5fVVqiCds13cTbmXb
yIaZ4TAOJWxLoq+p4ZIV6b9HYFy0SDHgWr0MdenZA2KXRz430+ahHWL7wmyHIgPih5hHsF1zzco1
gs0E/v/Fg27Wz4jyL/gEd4Nai92rPT7zCzAvHgvpGYh8TWmygXzAPypqbWXAqV44yOqIdg8KZKu0
M6ebiv+Fe65qc77kQaNrrhQ68LrtSaZj9BwTi9uOtaGHptRFGwMfq+hSpAF/aDiToBohUeb0lOdT
rEWaayvvCYKkt5tpaYhjKW9jLsYLbDQ8xAVlOTGtQP3vqVKjbasTFUjjgD5n9e/Xl96M5chRNbsS
dZwTE4uhmCs1OF0oGLQG+70N0diRtvXxRsTM5ntj3t0b55PpbrEDSQcWS/KAHiXSARqhaTJp49HF
xEuyY+mHucLODTHsGccowQXrBUKkBj9Kp/E/Apo0217ICQHp63l7QTipUk2Mhfz2Ir+4pfPbz3al
Y5oJVJhQtbISJ9tcPVJGJDcwDf46gsPrydA+8iO7Bko0pr9A/xHUvBCM+jLFZRSxicsH8aMHTmwm
hUV8n68ue0F2xSS7oUzQq3iC27KcRLwMUpkmixCf7feSeWffeGVQxhhjZvHJu/qf7QbV/5BnIhR6
3N6GM78IhMxJ1VRz1DuxcYssO+zqtbASB1IWyJ8c359gcW9VFWBR3OmNCdhoMvcGtLd4ra2O+2lw
FNqO/KgnGkZAKfPuFIy5MljLdQjpit2e9Zh0GkJUDdDNkOMS8Mty4qyKJYz2kZ7LuhiPj0CeqoUm
pZ0iqQPMyZpN/FDA7JFymg1RhJE7+TSr167R0zyZLsk9Xz8MVMnJVTUwOW99F1/pgjr5FbIWDj37
nX14S8TfApWZKUJkjhMeFFKq2Qdit1BFTeIkdSr+TOYmD5EH0PAkH91I+MfGjSZ7k0b1sDp1Cwwg
+LOXCvDTe2el4/25GdJexTQmAz9qlDcE90Uie3wHqAjWA9T2kolEySTb3u8TE54hdrG/IPDupxT1
f/Z8qpKs5kbIjHkQHdH/fbLzve4AQ0rjFhOATnZyiwagCDoX6IMFpB9EQIgxzC8TLhWESegbXkjU
/o20v8427glVjho3ml8hjjm2tyuwiurmbdMEkE8xP1L5MPcVHgp7Ko8ord01L0+S9HoNmVWTXkC3
JZ0uCED+tG3bkN6eER4r+V0oXrDjsPw71+p7aqnsomMOR0Ov032WT7TZZv5M/p0sFltD/dkjBvW7
6mbtnutTiBNnuM37mELRZveOQ+gsRimdzDwSZg//NYZjxY4JyCGll8sV6pt3g5RprfPI7i7CloC7
+WO47P8yVjZBPicqeiei0QD+FWHfOceIjX5QyH+ZKLX5WbISS+4xuVQsNLLVqSv+1GSCYT5c2aDY
LJbRN8j6s2AGWE+iUkYf39PLmv5IVbSfyCPU730oHbc3IVy188gCqe+vgkPRDV5sAHeydSOefVvc
ENMKgyqbL5306UZ8V4pAoxlXbmrKcT7lcS28dotNlFU/LBA8WTC/ob2wMc/MiDKo+EgoU18Vn7Qx
e+V5t+c+wQkWWKyYxSiPR5SOUXwtqSaq89fDGWFbzZO4vvOvTX94uu34P3XHdhrNCegh72bxIdAx
rqZshhjWqy/BF1UoTpW1PRqE8X3VTl6q/LZwNVGRIjGReyyU+ebfNGBCSnv2SRXPsy4uZgiMDxsh
hKbE/5JllJzsAddpXv1U6PMs2xmfcmAITa80HXKUrUFUEHdbDIN1NZd10zOV2m8nSfHrLXYa6Jr7
hpB6J5+5D5DgLuKUTOp/1M97zg2CmM0Dm3PndZamyrIcbN9ghCUbEC1E4pEutloqZmoVdILyj9rx
R8pBrnmIICtuTcxkR7MYT6fNbnTLHRyBSkF7yJlM3Z7sMRgpCFQdV3mBIAHKHo+NNm5mcWauC4sK
0q8AxWw1qt3UySsP+8WIOeHY0SciGo8LdppmO6WIoKRzBWzv2K0k6DN9kosddyheRVebtplnWovL
gk4u9ef0rdJctgl4Q4xBI7cZyQF3c0+O7M0mUJqfmDwDtax9++BVpR9Z44UVHwWF3FDG+hvGv9Oz
Ryr+fdwa4iArJKyY5YphlwEE01vH9Bf4knvp/yq2/UQ/pnk5qrj71UySpgzt1xMyVxyklCiLlzpk
Sc1uAhWyK0vmRMiJVY595LMD81W4yqiM9QQBh8Schn9qW5O/TqikpiDFdvX2gLmT53bHF5WC0XaU
GBBpBScSsJdmxYg5eliXNZuYI9/pN9EU3EacmfNUayOPhnzRaHKKxGrQq67vAdcFeqefSwICpGzf
fXwq6RGtaNmhnAZMcbAM5PGauxacUHMHQ1j4U+be1EARPj8+4FOYDm7agaJEa5VACVeSlgd/uLKy
qk+FeW2XY8K2OApZWuL8dlASz2AwkvlmTbxA+JP0h/UR0FWVXeWXNk257FcdHaae5ZfbZaCXCb8U
cQekbZDks30k7ctp5m4TmemR6XrWMJjYhC3+hIfNqFJdDDZWOyotLQJYPo/hqRc+LkWn46bWkN9E
QxOyuFI5e0SJEUQF+S3hVtnyPgRkRfZvjNPTaNlqCOWNeGy0jJsWBzbTgQIXk1uaGRX4VwVeujio
iNForOSRhsm/ealHPm3Lfn6o77IWhNh5cRo4nPWaXJoVWHfjDyKSlHelAnpMBD9gQTkD75q9DPUU
fU0ubdyYwFa4lDKrEfA9320Pdmr0CgCbN3V4SERMzt/ZfwnT3WCKIcpUyPDT12dwg5f3E0LeZQif
HfLR9Erw6k+u3BfVG6Y6Q9/QNOyYihXGEFS7jklcgMCwW93wp6gFBdYOPsKEHCIlaD1Sri6PD25z
tvoZUE/Re3dGSeLJ9zE4o2Q5EM8ffzeIMdzazru0dlcysUN1f+jmuEBoRURU0LYpw4ZWWwdh+tE1
LrZ/D65oesi5MBPVf6tpIBMWDKScm7JvjAbAurKiYTaT0MVvDq+QAs9454Wmfve36KCt3EvQSlcM
CKtqSIaQLq8sarGcLSdYNolcsz1iHiZrLHmf3seUEkdzjyHEzd9OdcOVbN0VPN1jOnwCp5f4LCym
3p9kxDHMWUovCKjv6PJzjikG9vuK/CtDdb3upaDJKNoQ41LFWRf/+1jy/84zl8KldaDDPU+M36uR
udb/djG216kp5njtBhqPUmOnFCmj8DSL3pEzJfzhi0K2kuGrnS5BK/EJHbW82K4FEbM9XrnqCMv0
3rxN11vInOdqS4hcEuMtfiOWKYpr3kf9DpYymr+nnMnc7vtlB4/0N3GeexY1QUhSxVo9BaYdatm3
gPeTnB4gtexR8zwQNlb0vJAs+EsDxbeMD2OvezQH0hUInDKnZdm0dkoPdpvtpDGodtK8oWUTsG9j
5kJl/4S2pXsi0CffYIZfg6K1rNOqMOYk2qC7vpZcozVtPHwiV6c9EZo6M58eWQ0t29BhEBHwylKk
R0ElsqRsXWPu5mlgvHfkUOJNUI2XrItsJmRh0PTPbGalWO5ENtU7Rv/Jhv/wChXj5vdHDOFnr9z7
KKfaJpja4JzKUUA7YRl44dqKLo5iD/cVmt7HBuDC1xJmrxns9mmm/QhBzHd6QAqPXjlhMG0y1yW0
iu7G/j2eIpSvrAIXbe4QoXD+02/VKedKqgGR1DVKT3GYifQGWpGribbRincbHYuSqByB95ps4y3O
on0H8ns/ItvHPEhzpMIOVk7OjJLgo3oGBV2QtL2vDh7LN/lCtYsdtr0A1TxJ6XAUTWWtzogAQUUb
6nzNSJjzJQGa2vlocAYqWYmTdK9vN5AAiUm6Si3OSlEDY1IixcHEIlYJRarWLFQinrGpc+/N/zsb
rzctGZt48LccCCXkMxiq86G/FcbxTJgO4mP/S62+nrcrvPVXPkzdFL7TTcv3GGeLm08LmHmHvyx1
sUZoB/W34N0HwwVt7dlGBlzFft5qu0e1l3MygGSqgYZraFE8voBZ4w4v50lr2oFrbn5FYby0w+2Y
aT9nnMQhaNjIXPsjdS9Fy8elibPnppxTAYm4d1M1BZ540ggHHbKFgekfY00GfVTpnvgW1wOnl/Md
+UXN/VFdnKZIdZyDB9TQbaejRDXFMgm5RhIZbHDu/OSf+BMXABAvo4jBMsbDLBfkz6Cw+fVM5tNa
UoOZAbKuZ58C3u9D8XIiY3SD0gzfjjqmdLTorJTpDFG7cEgqEqZaN0T5x1AcIWNAL/ybPkKCbQaz
Dd6y07mlitN5If1cymvPQu0lYkxtoWK8VbtV60Nmkxo9LQaY4xJNKvA16na7wJJ7CV3GVPyMFhlQ
VpjmPzvxJ+sv2ToP0iuO5b8ZyPH1CEFHSiDXCvrEc0RebhQ+E8BrRDXHDo/fCxovoRXFem1LIE1x
52AqtT4/qGObh32ZEbyD0Acz6nKeJ8SLyGVS0hOvUsSE+Lnw6EyxvuUuWr652zpy65Pc5vn0lcsO
1M2k6TzC2jbA3xwteM9WYhTJHcdmVCyMsz478C8K4q1k+NjT4hBepLnUxl8tBETU4m8ukixca+mW
BmN/WQ3ASgm0C53t5dVY4PsHf+6r20Rj88ULE6M3BGk8UP0chgjLbxlytFP2UAoFCOePRDdB0So9
u/VJemQ45gf5Plq2xv8kzzixtl0t0Ovil9AlKQtPPey8QvFOR1VQuQTASttq00w4BkVUtBTgt2JS
x5Uu20xSa0VDBAJKBNVvqoQ0N6JmTa6nkPzC5ARYLuOmKETAABP3oR298PvBRSSkmHOb1Yo8NwNC
1Tq7hq9zXyUvfG52AZ+C1L0464TJ2x59tHnIu3uMQuFsN8N9OsoF+mHs2rXbwi2VXHt8SCjeb9vv
r6RAYdOyUF5yPcMB87ngxu1xUAjmjxVZRRm0TcI3HgiUYS/uBICBP2Xtd6xdSCT3mv3o8Q3virpP
O+oP4+Gd9osao6a+uAnSKYMDWJID4ikgtsgsqt+mOFXjWIBRddP3HagX7LqQwgxYjThiVKZMu8Ax
UxVyOKKwFJCIjLBSqIsWRXEWtLdjGi07xmDAvotdm2r6uGeuBvZc15N0Y9PKTX4MdKUd8GFLBVKO
FTD/u2V+WcZmGLdyyIZDwW1lrnOVz72JkdNx/tQpJOkTlqJ/t+96jMO1JH5G2J1mNrKAmmC8yq+C
fiVVLZcnvlVXzXXiKl2ebO72UY8brP07Zhqr/pDZapcZI8iJZW33fzjkdBKn94WnxF/HzdLE9lPg
sL2TJwp82RsZAT7qfgRZ7V4tX+Fs7eDGW4MXtwrNNnNj4s4+pqjFZKf94VugkKoKrUc+s0MeCzc2
4N5wS+yfAsupHyzAIRMP31fsHelc2bbZrzfuvkLnGDn6h4uW+ysYma1cUnlyYhrKRHqjiw+J8L6z
Of/biuNsI0N6moZL3Tfk94obMGLbp3BR0tNBwiNhDaYqevTqEOsIyom1tAMTC7CxUBflVt/iJu1E
vv1G/pnHJFG3C3vpeEvwgVKVFn9Ofj6AJCQHFpC3go4bQT6tXxkiG/W9/S6DzvJ7u9R+/fgdgZIX
nwrchc/eIxNZ7BTXwRfRkMt4sEn2vjOvm1XcD4hBy6EuZDGoEG6Mg1WIDlRMq029XiI7wEvZpw+E
CWXC5h1/GMabBKDsBZIInbXC6/7726SYrJAcsC1A+Jaq6aUDrZ6LJbn9fZPfHnNg4sMymqHSHo/O
XMWDm8lLR7fgJEB3aDQgb2BLvsxuTuzpTiENSFf+6CVHExlofm4Hl2NpLEwhykOq5vIoaX/CzNB5
7jYBU81jd7B8c6fWwI5vcGdpg/+yNYXhMUJc+e9x6PGDUP+ib1mSZ6ilECxa2W+cxvXyXPXBQva2
zDoW4vlG4E6D0WxtOJIaIX0rMW7wEErDL6OqSs2ET2UEGeECP9CPUtQmt+UDoMrzKE6jyeSgjfOE
ShJsovIXwebxEcLFvX9FUmLyC9DvJCY/nCGfhXjNFyRueT3JskKiKClDQdDBJcskHVTcyE6XmV1h
5LeD8y+9Dtr6mbY58CWggRVmI/Ogai9qw21J3pjodTX/YX2VcFzKskuJxCa6y1M+GpW3aa5VJq38
BBK7RMzNv0wSp102cd5psOnas4i3LwKb/c1+OQoKgO6DDc0wLxZTefv9eyaGTKI0d16s2mqiHXln
N9ckP7dtQQDocsM+LB8fhEpUciUGaOExdSxkqfr+kYmId2DX5AbO06L0/zm39iShfjSBa28qpjaz
l5Vbq6WUU/VUngI/+SFCG/6P57XAZ8YiBi4RBDjXK3XqwdrOUcT8zXD9+gPPhicN8HFHQkHTx+cX
MqE0uoJW2oM89bSjQyvc5/L0f8OK+d+9b+Sj4I23huSs6bKCEzRnCDkhetTvFLKBoNN2Sd+Uv0Lp
f/TPjhQNvF3k3Z4qCcBHx0VvqaU4qtNE10tbLq1x0tRxcKOcGGCdaJla0xv2LDU//RPUiltB9XaQ
QhKcHaY/2UsJoj8zaVxQ0y4uUy4dNJnuJh5Wy2/kcrWBc1nMG40QZi0hwom5KNJCQQlte22TKvMZ
jWoyFtlM/WHKFFdsXSW8+i/15eE4TEZuMtx4n5W90d2w0NP2WvmGFc0LH7+EufrWfGDzoIg7Y9MJ
r+76QfcuSRSl9eTNtr5NS+BA9yXSW7E6lRS6hIaxV1nTW+tahc+TqrYPNCv/rHpdGyoQ/W2GP1eK
jZ7B1YBGELEJenyQEjyAyOwnUL5z+htaFkgHlMN4FIKEV6mqXEb/QgmmbTJ2WECIofL4G7v/UGHx
e3OEBzLDp4HunRN1q4vZKq6MH7ajNPv5M7frgnQ74d5MQ774zfacegm/ffteViI5oWc5zZRmV7Ys
7/qDjLsKaNCPa3jWyp5s2DDI+X5GF6fHeVA4ON3HayDxB9UkBoXqCq2XpLDCYgBNSc6JH8yRgdPC
bq+Y/PY18w4P4K9kqABj0F7/lKB9KEB45nnUVb1xSdubOzAUBSvdk9Zh4CzfcxilDbks3VgvMNXL
3/EzkUEeEXdqrgvfiLrursDu/jeNz0JKQjq1atjFkc4x/emXXoVaseWXDbBHgJBTB6uDXQgvIgKK
MNPqBaMVqBTznuZi9finqcBLXtcYJqBIO+Xrz+iIdJjfrMhvhW+7Ixy7DVXeSLeChFswu4sQL2W8
LhRLhkPhobUB6nvEJ8GG68x5b3rljAg6sizUCh3tGEUs4TI8h9XlBflCKTtbHbIzU6Ns0eUxwhjV
3rqO/gEYfstsGQbE9I/T3h/dUn03annTO0wZCNMqTr7qdVxk7PRRDu3OH6sCI+FcnKtiuVYeZojE
8GqpOGbSqrIRoyim96YL543XK6B776vV3p6VgRDbY06QkDPTd2i3ow4sOh+ZTwBlGOXby0Q7fOGN
yMMwcm4tjlSCOrbtSs+EWkzluRCNkV0yyfoy0s1G80DInud2DrQuI9U646QEiD48KVZKojJz/oD1
FSLmcwG+beiQuWHD182B5DJv6NhIFDw/aWoxsC1dOiJBOqM6FP26IMACb82ctU07dZaNpd7cvhRT
X6/eefGv0c2N6/Z97aM3BAuAOmnFZ3LMSP8Y1UZaBCVkYBU0ogU638GpiTpf45xh9hEhZZoAZlE2
Ln53zf9xns+Jdqb0ejOP4LG4tQZ4JAgKRKLAwYiB/kKLCLZdftNIgT5yANgvpIj+BBjLBuUWhEcU
JA9S5SRF3pBbZiSQZRYzo7gQ8GNK2FmQjJeGz+eBoqUXCsJ16j7c7rCa4Vos/67whGI4svWciliE
oanmvDYtfjxubLpRYbZ+1JYtUgqG4+zr1SpbtZb3PEljO3T1b1zoNmp8ujVofld5j/NxWeDBSTUG
shAQyG1YAuNj7VnFSVS4oy6Xyy4PBBWznD4eSZVxOTQaX/keOW+d11UZtWeLWAfpwkXHHkwAra5F
eQno0JlQo0cj7iVq7O4VQx09snewuZF/3KF/R7R+oMvOirm4+MOcDPdXEMHSgWfIo/qIdtouYWk7
JiodFu3IQM+9CL5cnRa8mHpaSWLtL1ijPscBLZ26Gc8xcT3LovhCfFUZJnuqC6TbatpC29fTfGcM
INHO6MiWRKyaRsBC34321p+E2sejq2WtQE1UwxLSdc+LKYi3MxLLc6XPPgnzhRm2AGJVoACmxOmn
4ALPiMKE1zVw8fHAVllpdx/o8ttTRdruSK48MK1+TUS8xaAmbWNr5TN12qQgKSTLOX2KRisfA4NV
3aZY5K9xAfeGAlUBki0z5SprbZ3LMWaSn6XCcOhUdtT9RAMD1i6M9QaIU8+/po16lQVjVX5Q/kcx
5L/Dn8JmMt/XSIQ8coVcxomQycryBA4verUe4mdZbNSlFirzjiZXko8rUkfaP1xiWz6HAoVBPl1i
UuZufpeiOfnjTnhFq+Bh53JWiAzIyOGTGKuO1/pHZC7ZjZlOfG8hnxMpVGE3STNmLbZFjdCgOqKr
6/u4wOb2Lm4AOiga+P90noUI3vPAzA1v0s9ScZXtzCDWm01jIl7j0dt/F9FyaH50QLlisJWMNlPn
MNWtMGUJbyv+o7U/6oCsvfZ3Qc6hTshxWDwCL9CIBrsM85F0MQV9jpPsEy0eC0y5yQEYijorA0Xw
ISqnhmBLFk2B4e0DQSpGJnZn26kYR0O5rqJ1NbngNCwXQR8dXOnccAKXGbHfcH1P/Wy1qorGydlb
2aqdIW9cEkvKy5w7cgfTuu30EzmOuQUHApjujAYXyniMFALX/ecDdEeabP/GRvhRRoR3s6yPssa2
nDTSqtL2QaDMgzV5gPpsdRuFBLFlxA/r9r6a09mNGBugYa5beKcx9NobTnvQTayN9tA6HRiSEmj4
BdGcTuxEvBAgXoJweJX57pUuX5bEOGTXiR4QdFInD/4VdLgC/xL2YnqcV8SdgKCJ/siAHSuG+wvr
eFPuj9aNBTnawwUG87GeNOF21ns+dKZrnvzmGk8keH9HalbRFQgAnw9458a0aZ/snardeg4Kh7Dj
DjrBBXb68Fgk+caYdtGcxptVWU9VcOx/TGvhg1SfW1ZICyY2Xzch7h81q17z46nU8lRbikgg2ete
15QIDhZoY0Zx5FU6MtDDX0i3IMB/C3Pdj/clueCdhV0YulEMYV4rQBqyjQ5YOZzOWMM5teW/mH6B
riWhLsM50ewCpPzUiJ+gauVZpBqvxUvEGn0/Ci9tErDmz2cIOXkA6Mi5iHgBlO+O1e1TU+5VHGNR
ZiobDIg244LuTJTIFxVqbSHn0+UOg84cFhllhesqKPf+MjoIeqBidJx/Fmol9ESR302C+N/9TWAl
8i4XEiY1XB6glHnz458kB3Ny+94+AmshIse2Z+qaf+/JW8RsUxYLG6UjHXbsnpe4hJUzDbP1Zt/c
BZP4l6X3mia3DjZUja5zjmSyXORwWz4zqj7BEavAZ4j+NppDkSRT3xn9LxWM0zLRF6oGdgM74P6J
cEHPOjOoypFEZ2l0uWQSIAS/u2p80IKUqwHldTk/IWLWqjPvLbD+Cefi2Lthx503ysXft+MW78Kf
QdBSYBTQO4TPeyuyij5w9zh1CUO/l4iRmMr83xrVNyJHk2oiomwDCBPKj9i287anaWXf+hZwwbVd
qsRTbFp3/9X7y2m9AhPeXCDDCDcWkO6G1f5xHMwQdHjPvuEV0BioS8ZeClpSkskHn+dtZ0+LEHs9
RbOKxi8fqEFWNOEWxXqV7h8aOltk8Gxr4ME6TFOSdbT2/AC6AkrDTAInzk1XMe4t/rGAGoDeoAta
bwdeDcR1DXpuNOAQ8476qL0vgXEjPxgkv4J++glLLdbCvyGAHGtTzPEVL3wI3JIvpbOBZRwNcLqt
0GJau9llLMk7wyO3ZlUp0Hcg3jjfophFGOBt/bo9YIS3SqenesraOy0+v2pbSzBQSVyPfA3/q2z3
lfE5dzbTkx6nUjkLy8vi3tyDZufunay17V2+dUq5LCLvHqGUlCiMdTJMnOiGMSKXgKIpo+wPKHe0
KY2/LCeKUtWgUWdqFHn5C20CSkqDnqHuYVOLo/Bjk/iJpo+OLyfJC3nGxxMYEx9W5Ep/bGBx+Yi0
PLtdNlgUfBNp69nl/QXh4sAXcOaNkMnoxvGrUd651TedKb87q0PkVqRpp87h2TGwhh5ikutwUR4C
Vgbk1H75A1cCR3W9WiHDzvsyh1mNNAxzsSi1GSpstNJURsSC5BXaD5O4ma9ZOTO3jikllgQcKjX8
30YE5DIReEEc7dRBMH0igdR6CsyDcn+rsSOw8oXVh6O1VoGsvNZZlmiHQ9F//oE8IZGbwzkMGZXI
00EAOHSGbfA9paDpwWoeIE9zNrzvimUkuAixDCvKVyk6OAA/EKrxYOF6qyjmOa5fOeuigbezCkUa
ijrOcjTmaqqqAFY/ANKxN9KLu/wNGKxkA6bMvEZ6cI+u/iidOm7Oub9xzY7ku7w1dXY5MJP/6Hd0
WmfiR8kkwL2+dviHxtIrArmHGL2sXDdxtFZMlv5yPhx9g0a0yDDG1jdhQ/cCsY/z4z6RR7jsRP4X
lmOn+JYlGaTdZ4I8ZXXEI7AgYYzd+E2BVg3hvwoITyuPL7IbI7xrseLnWL0OE1RuKmzsswN1fv5d
UpBTCzUcyPTymBgA9aveJAMypWAR77+EH6mQLfZFRKVVAarYIf9zv0bGg3YBsNL0KjOR2EjWG2Xc
mhoK4Ts9+4PdswjsHtJs7xMQAFeyDo3RpqgVg2U3co9vNRiSck3nbMEJgWC5xFJhz3Rg7STbb6N1
+ac4M+fMppdnIQFYR56MWUyyLUe8m2pFSEq/o9OSUrTKydNzja4T0/eOzhbUQwM+WHj/ak4QJQaz
ZaSQkD+AprmyasR5uBJw6rwFSldE2WIqUB+9cfgvXkZoE2d6vT/T0ColxNW/8hNMtcFaX32A7FXB
jFkvM/gyeLnL1CHH85pUNj8e4vnp57+/PcmawvLlh+nRGt2U5/bDWnXVc4eDcNjM8mQAx1L4Hohs
Viy+ku2HUAX1VaWF6dFYIMeE17v8LA==
`pragma protect end_protected
