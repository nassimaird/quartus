// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KlPrA9m9uvbVHYFtTV8Ypru/rVRmjksapTupIMkqPKjHn6h5p+OZQ0mENSy6ZhMx7p2+DxD2oXAY
+64qVtDewyAc5l3vuWwBKMh1Hzx0JeO5wY5C3pu6b6JzrvNoj+nByw861EI+K2qMv1TEcTkREDjD
7u/ccCQS9kSWa8QcucJVHik1I81o8DNpm/oPrpWk99b/z0MTTfYc3BZGpio8T8iSMGImdQB8lpQA
O1ablsZfPbP5LCaM01uc8ekkHeC4rjPeuDtd0oDgnASFkzvENxzvqLzsm2Fwzl2Th8lQaxp2wrZw
AdXINMDlLLWwQM6zxJ4zKE96hvwatT4RNfR1JQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 109056)
mR1GMv0lgf4r7xMOWwdGi2j/rjFzEGZOzcc9gKmMQOTf/W8SHWHXEFl1EftusCX3/hgoEux64VwY
DuMdLfeyjPXIlEuBkFN35/fzG9N6vpUH2ueXS0KUdL7H5q7B+Uy/LW9At0lO8EZAxwGjhiSiyC2h
ruSUgcG6vCxX7g4vqskTLYpO7CY2yU2dztYrHq7sfwldAd1kukYTn3FVrGqO4ES8qV5SawktI5+2
ab9oqYkebf6V/00w/RW05kze/CvB9uvdVZs3onlWSa43euAz/GNA7kTG7qPzIo5Kjc/ivbUCSEP/
Ojk+78IgwGxKp8Y5Ir5AwIlnZkip0m+XyJKPdBL7IsdnFB8sGdN9MqurixodotL0U/0rVaZdlkYZ
fJxbOaNOPzzUADo8/SyrLF61imdaV2l7K6KjU7qj/+oeyFGw56kKvRIsREQHX5GmxI9e+OLpw7AA
g0/3QXj5Cfh0s9eG30/cnHqhD/Abw5x0yhbdV9uAXWS3Cf5qr23cfnlx5GTaplJH0kujjXFshz29
ZN/G+Bta+9FT8ZgX93sWXv62E5S9UUio1B4p/KbBzZW/1toLfVjCYmhMfpxN6VXFKD6cl7AGr5T4
8rZ5gY0o19ZUZQVDr3F50vb6ZPVCijYn2YrbbagrCS4+KId6xr0RcmtMAzlmm/RonEuLWuopmx2Y
dqQFi+NaNofQ0kfjy00YCmQxuYs89k6/7h/fpWLNlLhzzJflqyIrO5d5jQHfxb0oKWMx23CG1eYY
+sCCNiWMoASFTjXP2omJJt5sPh0yP7xl7JjkojMb+Z3uKC/HyH0ycCg6LOudZHB3vHMTB2nGL6eo
LlcSC4Aky6jAQqJ/S4NpSdXg0ak5gX080yAABYo/rvmh5ixr6ajtJpArng/H/DCSOSlS6XGonFYQ
Fhab4Tw8RybL8/GZYdgIcxlhTV3n5PLuckqZV6by+YDg46Ku40WtgBFt44FFa2VtnuLQqMxacpTq
xEhaMSyzoL7vq1DYEqnuX46GMsUCX2jdmKawv/Pt+sNXWtKCzzeGlSY+AHdkd5nAEm0QGnl6YHVt
ozY4OdyrexV/dVHdTocFI9ocy35HoMPneO1rfanbHV5ECADoVj7/tfL27ExvM0L8yQ0lk/00yC+L
AhL8dnnSq2P/MGZc8hQrkdhXuBu7Oon2+VlVKEK/+mvNa7Mm1kf3+TVTb7GjE9EtaIojTDeom2Fw
QLNLzc9lJh7YSwqUwBealPBbbTRmZT3kfKxWWqcdPFSVcxrz1Vd1wYMDBeCHKrGFFLuTZFMgKHlx
/MTt46SoBdE/AWRxMby04uT6h/KmQxixQztHuIyN8ncwpUuWxapyUlGkgilvCYtZKvZ57aiSXPLm
k0tnRiHGCciaesmN/oNUbTC+qJtj9K+CKwsVbTwh5NkmW0ccL0NyqV1W+6s9E9NPQdybTMSb4Ch1
5Gzu9ABC1w6C+/6GJ50me2L66+AHnlwMi06AE2zCV197zDjtmBK/5d5j6/xopBoplKqkO3y4FsQB
HEm18mImodjxwW4wWe+snVM1CufHpV43ZTu2GFmWrcGvHuUlQsAI0Pc3FWjPB2H6F9VNEVXX16xW
R4Tk41jaTIYpLEIYfFgKFADpNr+2N5hiCrr9TtYUydKlC1TxUHRf5Kd+k5TTSqc/3mGfPwbA7jf4
bEeXsbcgBHjqtCosOUDDHpkEd9BQl16KDn+UTpO1vuav5TisPYTTvpUyItr3Mabb7segEiDRqclq
cvkfXywHXV9aAKhtdxI9YpIzaZfej0yW22CYdYqR1TaZCTIanNkAcoRNvdr1f5vldaGDojbgqf56
i3pnrPbguujxGq+EIhY6tze3ZjvcaWeEHPX/69K38zOcnEMkf9WG76RPvn6gC4M2U8QtmuICkxTt
vwucud4AFzsJDuzSiQUBTQNEPwr9t3pAgTZaZbDerPFi+XBoxon5PqlU2IfVt3jFnR+afzN/D9H2
J5rwWEi1r5+n/wl+W5zjzNc7v+lrLjQATFnvOS5ocaOlgfNrMqUocPpTvlOR05rFNvUfnw8mmTZ9
7ERD9CT16CrhJWHDHopawT9MNvfRq/Ip2ngC4jgbdGIlKYyDN0cpoDgmVSy0vuurVNhewr2ArINv
T/8g7DvJIxEsU8lp8vlnmPxQhfaXCVfkG/5N3D6hB7/Dun4urFfKTsstd5R7rR2GUcrX3lnTPa7e
X5stCFkd+Iy1YyOJQwF6tc2YYR4inVIZtX4wEIzQLkHYTRzi9WqW1vX+4LJyDM5DIPO0vtC+41ZR
78Bx/Wk9zpBM6m+UUrQLKRUbzZakmj7hqSJzQmjcn/BJOMTtIJVcHrGwOlOaMjOotObZve/MeM/H
0U4mIAaon14+lN5NNDnIlJIUg8kRtAb2BMzVdp+SnL76zjrLdcujQXK532N5rXdmPIorEGgP1iEs
fAQFnFqkX3jZI1bXDK3l/RSx3EXZsRaeDEsAqtqTajuYKAeU4c0MxDKsdZdXGjr0HpaHy+uWmB14
pHB9AtDoS+h9Cnpofq4GOwZ1FBCgpXXwkqMEkAel1k8o3K1rmpFD4n4Rx4f78S0Yq13iVh77YvvV
gqWdrNTD4xoz3RRmghX9JlpQcEC+d4ThFXUPhKna22HLP7t4dbwhOU6bPwQ0O1cyF/mcv/XjCPTo
hONiG4rgYASaubbJrkXin+NDFDQArDPHt35NxSg1o2QpTYTaEu8FIRgc8tsgX9ZzpbIVoUn4bnp6
PORxuPVud0giS1F6wM9c582PUX8o97g7gFfkijPwPGh+5MsAsCgl2xLMX42Ibx3ZIXjFvSpJJs+x
skg9Goq+htU9mYe8ydFgH9afdVT1jP+jf88fUa6rvKiy6zQWm7eJm1x7rdOsiNERYQrOFJcvY2nk
Mg0Bi6rUGjDA6SUpuwvmj9YHwO5MzYQO8OHOWQ4YMliNsijqdfYHn4U8IAIgjqJv9bwiMFZGbP4x
iAqC735lCX71dpCiP9MHW3EJE1El/Zxs6r9sueKtSeNjatOR1OiGQOXbLjihy465DvxhqKC6jH1O
yHSHz5KcLcNJe85PUZvcFHaPDAN2n0gZ3b9XVdTdY/0As6S4vQX1fQj7if5uEQi4+Y1nuHcN2/Zs
dHpxVH3ETd+Tyl++7x+Fsj3KRAn6xEjW7MF35WjM7b4oAiNfT1gzggJFvbOUWwxBG8wDuVfVIbqk
f1i9xCHcgrUf+AK1C/4kie1EkzwX3gznq/PEYbkAygMhQALmLX9T+hgKQ/JCsMPUubn6mDHNzQfm
idoaBRgrXrzCaQcK0SHcEGATyg6eO/8LFItkExwWOMwyUMTg8MYGUrMhh/0Rbyo5KmvYqur4v7we
iBnmq2tQ4OkVDD5djEQIC0n1y46ch50RRlO+5Rm1G+tXvcxadsFIrRUOYknea9Uu7mCu+bkbRdSJ
sncS9fIzPQGPJzC7hM/xpYdOZSv8X+Gd2j1Pf5cnHqq34vmTkntIkxyE64DxyNhlwgDWMKXpA5mR
sSY4Cabf26orRN3NmQKZfuwEiKtL1z6Xs/L8Qxoc56pjr91CQIA5Zm6PjzKuQ7jnnCNTy2/J2ywy
aIoK/ds9LxGRiaGb3QIHpOqEeGMxkz/ClccpPuhISs81P/m8uSpDm4wwp7QLdfaMa4cejlQkGA6/
yGHAniAwCHujlW/DOuiAhcoM9bPr7U0Tk0yZILLA0YF+3JJnNIpGuo0u9/CcZlXqdxw90ypePxUv
OfDsqGjtGwv+LWBMU6fGf2CtRCt+6GTaPrjLZqwinqk+ooD/eWoFRSsLCWQTRghH7AEQwXt0psBT
ZP7muvlo+YuCfThuy7Yok+XN2GXU/NeenhYD/gquScZlodnmafD5YgN0Gd7t7D+TQM2c+w51DaFp
qgZ4wD2fWtEC7sSVex2brDXOE9NLe9kDMwV0CQZuV9ZFjsLru/V6D3EcExAAfxcFYDLom86aHabu
d31ns6DXjrwEYpRAFXysApXUFexo/yTMnZbHn82U6MMspk+HnCq+zphpqHQ+zF9WotqZIn/JQKnJ
81R7KXlhQ9J7BjBXPAwAcu6impI//glkMhodK4wu5p0GMu5qLQexzPKeoRiSGNV9K9X2q1Nu38QW
YV39FRJdruVR0Dw1oqFEOgn+IbxDnWqEPubt0tktqay0p8CFi91BD9fKi/SPHswum/Qefbp5t6BJ
LMvzDGECbxL+nFn3wHrhzMwdJT9kZkcF8G9zE99LEx2LGUo3TFKScCOdDFT+yDVMzhjCa0qiwbw0
r3kd1miF88l/lFEfxroYCwl1AKvNeV9q7LyDrjg8svTwQeV3vyxBTcn3UWOnxVYEz8VauaClqQPD
vy3qzyM1FF1YwCP/5wrWI0ad0PSUBMSX78TSrudT/RseDUvqAX1kC6ELvHYloQ2W+3/+7jKozWRF
/ncesgcRBfg32Yw7Ul64jqAbeVCBOqRqYr3YUBzlHN0m1ePIwf16EQ1x6UBbevJk4wGkmzvU0QSC
zbLgcfn9pACpQ0uvxK8C0+wSPOh8T7vcva9RAqHJXetzBw4L/CVWO5t3bv/6ypoii9XiuR4SzLsj
Zya5VveY9ngkrirTbDzbqvscY6a3sSq5cTxzhsvTm3aLK7aS4q6jWCPgTGEvYJKkXtDJZr67Jz41
cnKeOSX3xyQQFNZnq0vAh6Pd6j6vzl8MJ1GfG0h2ojcOy8Ci/WlPeozRGHtl2/NjKGnvTOHfHwGG
LJ8BH5RAidUEHsh5ztlBe0d+/I/UwaCeK38cK+a1PJlDc97WKK1vg/ITsFkQNTdYFrHvXVKiuUvp
vsCE7Mj6ocl0z/Ex004xcn7TyQBgUBqGjP4tI9pv//rK9UCkKp7Fi6TZzLpJzVpnDUlhufycsyLw
FNANu6q60AmHMGXtluTvVrVP/AOKV/Mzwz+8ztIhoj0aRsj0LuMD9OP24BsUF8NL43RB+2z7MYYu
abWYkZ6J98wp4bH71slMWO/bnmaxvbY1/chS6ydP41d35Rjgn8DvPdskDjTQNfoTEf+qwCuS+JHV
psiC+mf1hQCHzxCSzp/haogKv3KFGWpHoWLN6HRPosnajMarkJnl80UzmVjXa8k70y35jPv4Lnrd
XnCHBrENPydReL+LUKwaiSxzmf4ylW0wRY0DhZt5GNlLap+A8ENGGGejgLNxf6jeNw7guat18WgL
pX9/Pei0Su2AqN0S6isSsQrI0E4BVu6qV4nXBu2wXcoH8ocmWV/VSnYkkL/AE0s5egTz+aNaKKtG
RTc7fuDPJzGhwR127qVCZSW6k1y5orOqkp95qB02XSKbgTQ3YSJG9hoJCK+4XLhazbNHD1YhKbXR
7ln3x8N3e3IRq04W3JL+hAeSEi2YGLEaxOEJx3j32QOQ9if2rD1Wa3jzfDm63PsFv7pApYNrDGbR
uFwj1Y1KaQr0jUJiNpV8hUXIEHdvWokSeTqyrUXq55yUat/Po+fBB0xdQ3iLTx4OOCkdmi8iTQ7v
RmVoCONqH8PXzOjDL9HbkrY3TyTmWycn/X1Z5mhdnSE0tSzwQB05AF+UJFdU/uNe9dfeeNvcJYlo
t2//9AFiE12a2jpG3ApfBQ10y8BIR1xLvPkGPri4E3ewuoDU0/qvu2G8UCvUxeso2buxiLx1rZJc
+aNGmn8SirmUi7RFL0rtnHRhhQlQOY+nIMPwob5RDuO0A4m2R7j0vWkOgnnNUi33M1zFa5muBZav
mfGURNO5jGokOQLkQBIA/iSs6mWhfQus+kqW0dDuLY0O4FyJLu+GtAaXYE9z5KD7VFJTbbGs460K
ZuH8zIxgrc6KwsgdCE1sVa15dr7cHAh7/eBLQGqyfBzlRC/y/JiD2xcI5EjSeXKojHon5NK6mFCU
BtjcqGzRrsPiRuJYULQMshojJlCTwx7AcSjfQWFYAYBp/+NduQtiY2SNEvNgiyO1KOsZgu3q6VGw
FfXRKaEUxaBI/0zwbMM9kmHgKwQSMCAcDrYq5V3qpUcSYTQMzMMc/MgiXlDX/lbtUBQA1/q6DKrm
4373JISpKWgJzNo1tSYyFqiV2yRmZAPe+bHDU59dvTm/HhWxgBwXUReQX7hhplr2+zXKPg9+Ytal
UtvsO2PZO3xCYl38NCRyrV8G2OQmmT3ZxkmBNztBe5lyi0u8pv3beA//OAewz5QHERQKRW9SWjlH
9CFjeJqS+gFoJw0xk5Vl253zG3ZTHJA6j042SY0mXNSrqjWbWXjUyXKx31IgB7tDx8lsZaxizoJx
1FyH+QhhwVWNYzJ7gGCFaAg4CLY35q5mmeZR2jsAEnpu+rpF3wJrGtPTmCkUQk+dW2E283PfZIZ9
IE80Z77OJXw7fcuz6oVdgVpheARqKnaeAIEjOHXtTTtl7xu9u0RH1GsE690xWxPQVWisYT3Wi+gB
VE2JkNseyvwp0Xc5VXx2M/PShfQ/d+Oer4U2BEEFG+8rBHKOYVm/SCl5Hiy45bkejr5KwgrC3Yck
VMLI0HA8J07Az8K1K+emY5fUEu0zp4oK0E0oyCZFzUNG4WhKq0cbL7o9FvUJ1hT54OT/5o4wRZQs
uvPinVf3rmJMM2Oi4wIpQQwYO40auJNjn4qvcrbw4vIbYW+DFGG0x1wrvzOn9bCKDFxZMaMbaqfy
psQFIJdexC91V5GWFHixxTfRYWSljsQZO9FyR9fSM1ArhqGNWGpOBSY+oKMVpQfNP3eyNTTF1cMy
FUQh1/NQb1rbeonj2zXuXnasuuCLYBfrr7tclmjI0B47J9vV53TRFRSiHzWJq42jx1oNWoKi1UJ4
U30PGcEjDjs2gPIIzXcFfH58McnYyTF80/g/5GGs6Vo15bA/o+c7xHncHh0LciTGz78E5/Nt9m5I
IqcTFcPZf8pyIIGcDBGvylyj55MXrjcO9D1qcnTLg9W23KyPEIWmHlqQRejHjT5BMz6Dy0Hfl8hq
+IZt3FOuoRACrbgaCIacH9+KimYdQbdlW1gqK9TjXSUjqAdQ+KXL5ihpjYgMpkvnkzK0aIs6GPzI
UnGivyUtsdeqMl9CkAURSr0JzPugvyHvGdbqcQP/z6+R4gCiafOvGGr/Uj3jfXUT8DzceCOyu+jM
PVxMLUpKhgIGPcdyc+CsxT56D00YwrKOQO6fMqC8hQxyHYz6UF9+f/U+NikusoM0CNxWyPRbh6+u
d39PA5cZkDW5hTIZH7EMaxd0qotiVniq1xluHAxX97i6Xk8GeYIi/azqi57EkFKjIpVbFgZPb7oP
izEL1aqjYKyvIBVDWNWyChyud36Br+WohWvbkw5D0rC3jwOmAVShnvteAnbYDkWtUmXXy3fAYuB1
HX9507br4QEyfMblFhb/NMH6gsjv0IR9SewO4DFkD8Xj44FkfP/NC+KLwuIFDqSj7j0yCaXn3E5r
fjmOACIOPoVVJEspB8uftTUGo6iqqdIUL0k+0Pb/YYzQz/9g3EaSuegUUHXv9h7tSmWSH3xuSrhm
1lbMpw4ds4nPdfBUj1ea9o+yOKhJgRL1Pnp4/x4TgzMniRAxDW5q/T1o7EwQUlHckBaCtoHQcy19
s2nwMfc0talB+fDP6VXO8B/kFRkaciFtsrNlf+HWefN5cLPyUbTH+dltIpbiB3ibWC+ZjlYqok1B
L4S6XrVj29H9yAo+J8QxinSk5lEEqbRovSnIQxvZwTXq3d9t3PPVfaigfkAXHI3mjEOLZbNfA7mL
BaH0Ux0e3n3pBNAjo4Wfb4C0Y7fcq2ZFtFCpofbrDrCuHOLTWIZKlxVXdqwJVYtDzk7krWjWOlhU
M9itT6IAzd2b9saIOVFZyyPuidHN8ewmEqgocvlr0evEljPYoXaHtXQNNjB2k4S9dMgYXKBITGPJ
kOfzBzDaaHXwXqudErxT2EgxDLNIMOKMIaqC/MvPcAyA3rLjNHOxS1pofSF/K5/78vgSfyRl4PoZ
llQKzaZcLWifgAP9Cy7EVa6B7cZ0N9yb6abcOpTvYHvYUZiyX6GuagJ3p+EVb1vCtOjoqbsmfJnX
hvYpThaD5u2LmHYB5PVZ+szsZ0GQNgwE51ODvVrNNZTIaKGlLS0WI/dueFLySacAUKu5Kv8TK1eP
PxB9diGsXNWqxy6K2amKWs2y/VdX8dmL4BUnbhwV9XfHGvQ3hzmog5idFZdwwUPwZUyxpe7Kc5Bc
QPJHQxUgoGS2IbkpPrEXdNzW6s8bwZ6l7AvnhHIHk3UHjoWFQLPx/a8U3JyRmPkM5FVZgCMZ/kUp
lzDww6cZzRAxEDjwfgwBqLqvkTCUr8ssfO3QfEjo1Xo5pLMYXeAZA0aRMZOKSuFDrbGtKZ5BiYPo
7qNjOKJb34EVgb2IqiBRcZBZkQl8Obi721pokLofteyZGRDPfK8mE3fropDU/VdRUEDcWKipUGpZ
yFViy7pz4zaHaQUjkgX3ma5PRRQqotxjjO33Yu3eYvYuJ/dDpCEWTsqi7qNkQeS+ja9uvhM3KHhz
Dz1phcXt+RLOIaXW1+piU9S8ecnTmevvWZ6lpWUb43M7JlJdnJZgdrpMXVWYXAQS5+b8MfBd96hF
sQZ7TseaYmWHczGfx/hBJ/zEgvfb8/W6IXO09hB+SSuQqeMBSZ2tEUv1B+0fbNERj8YxYc4jGrCz
3FZz13dkbZgvTakHYBWEfYXktYEoVpVcrhi5pXKQTOl5HrMIOe//sTddSrlFkUKhsxtvpi04oQqv
Bc5CpMhwoSw1NWzgSzwlpADdKf8jkcTBNULR4tkOABS5y6Qvf+r9WASHiyEDzgfcLymdl4bxqe6U
mNtUJ2bAT8knhn0PwEsFRz84qKNqrdKbWpCYcZ9DE8k+WSRmpsHX1FiVX7zXDX0JATBMSoRImosS
mwTJEBkd/eT4NjmonQFm7tMYGXu4PcKG7wKIspJ/DP+cdownD82W2d2m+4nq/NizEQNOLV3HDnbk
PH7j41fVgk5Vjrx284wCfT06eXoXXO7kmhL7ntSXrd6DXR2cq52XPVxrFANLOR6EIC1VVU/H8fs5
NN3NcDIIqptrSP4YSIWBEKE4tacpndthBDHeq9wkd49sMMLCmLMDjsdQ/2YvB9JlnQ0DLDSFgyPz
xKl37xjnfW2xDmkd4vklRyK2YResaiPjgE3sktc0bLMXaRVlqeMSPJzYSj1eN29qp4NmJnrU2YT5
73LJ4mKJ8PGDKjJqafw3qRhRdkz1bmLf+oSp8VqSxi2ZlR8Y1uveXYg6oUD2gxmYnqhU5ABadvRZ
eHh9sZEbOW76TClwkmYt5tIztxt8r37AcZ5FggPntxH6uI60G0rOLM1mFkM9QR0Bt8ILtUXy6hUp
1X3YEFoON50Y/KIwaw3F7r3Zs0JaFrVtoZN4zkJrupC0sshzTnTaKQXyhyE9MdoEiBTkH466mc6O
Pjju2mCEB7aaGN25X8w5qw/jcEYNw0KpjgTtRDKSNQN+SQRCuNkuB0/ppVfN/3QqstPM8Lvdq3tE
doCnMrbuC8OaCqWPl2NIWJlN5meVYgeCdB1kunjq5YoeWipndVuOpJjDUeT4FdaSzI8HXRnSCqso
mSkYYJC8ebdhE4TIxr4n8dVnyUSR1R7IaRJX8mIvh1byL/GEoYYewIEbD7K3A9dGTFsw8gJZXzQy
X5Rdm/j3twZodA77+nRQC8eEMdJzT0pS9UdzDmaBQ8KtuBie+Xpzoa77m6qh+0QX5k8Lv0AArntJ
eyRBB1sif5hz/+YiDH1I0GGilPqcRqPpNFUPT/fbsyMI3J5g+nC9AaaVzqX9edU1d8ow+zJpq8dB
o5AA7nVBRe0wPxFQgx2YO9PIT68WvRYKKKDAWCDumgas/00GycTMqJWUgn+i//5Ba72Vuvua7VsK
tD+2Tk09iXQqpefB/kPqtcHbBgh7Rx6L9JQOCJh6bpTSZ0LGRNrsqqIP1+PSumeud/IxDzStMuED
7RH9Y6NbjN1dQ8+awH52itlK6LnzlB8BPilhbX9eZ6fkEW2tgWp4A3cjlxEso4miQVCrYaEd7bMM
PxH7BGTqKIrCiTnBCTXPkTPsZCktR0oNt3fTir3N7iXNZqiAPTCSpob5zwzEhpE0ySdeSGlk5W2S
pqdvkUfx3tt7vFYD19Dy7KWDbYNbE8DsJjryrgr//ZS+XMUAmbY69pKKlFFzip7Cj2jEOWViglK0
sakXl4b6GRpPn+1PxWTHcyFla/LjuUb5suKD7p/XoZK5j6QLmaoYQC3K1c7Ufsqv2v/IDcbMa0/t
5YjoKZn1TYY5FABrXCM1kt1oYLzcb6WRneX621OnLxeyRZuFjkViF09TOSWF7teSj0jrvdzfIXT7
Cxnpl0UJ/PeGKzeDkb+RcORrlnbFvnvpWrBV+OaJ9ww2yIhjK22nDKabkZG5RV48xrE1SSdUjf75
AiSWstRADBV9B+Hg3gXOM61PsM0BAnMClhuymuA1YhNcsWIJ9AAcutv5TbXsVvAxGdA42ZmSYrSJ
HT3LfVV1JSB2d1gd38OAjdW76vrbUMPr7GVpy4wYpO637Or55WxaP6EDRDbhRPfndr9yZVOByEGn
6hhItT8PihR1zR/5iJlOCnzAuJqbrDNWznTCjJx45IzlyyfPhKLQ84yzLmPZ/xvEgpkQCkvtOo7T
/Brwlg+ZMMl1utiqVGC7s1BRenopZ0bBAd5EeG4VlCVzc0FMnSKhVz9Vems4F9Iyukf+2PfHLAAn
SOLLNWOR8Yd4LFeqgMOlaYWgpiLdWEvL6rlpFhnKGEkd1JboUdlwk+v4BtwPMMwlF+7I/F/LPzTr
R7OXapLKK+k5/g3TS5/eOq393AQlAZyD+qZYFxsb8EAqhLuOfcTfqZGNO3pTD6apfEAHzLaut+vd
LDT3ozC99CNiyOnMLHzXJoBQ0ctDcqlqnFMVAjDSDtR9hJ9M01ALOpQ/DtyhMZHImnyK+iUVd+1z
WWcYWOE1/bwaDhcDFn1x3Cl6qEGVbgTYtiHWoKOAtcd0LEv+hlJnTOF3hT9Fw1c3U0tbAboOg7QR
un5osFCqUaHuDzvOLI9P5Mx7b7HxST5bqhO6OXbQWTrplMI7/XgKcYyPAqM6BvrkC71qJpr746wS
fkiHqWutDUcRmFITTIcT7WMop3avis+39iraqLp84AcBM62hdmsKl8mKRO7WSeHEBj/E4E6b1mm/
RlkFMeMgqWF+Vjn6oFoMKlQWVOe1e26aeQZTAq3zD9AmpoReV4whV1asCVGI+xlfOJY6x/viqkda
L1pLCmzan5LFZURyS9Hb4VOulx6bKrNsphHIXg6NOfWDOVcHY0aYJlDaAYGWncquo0DYGqnPsngV
3FZ57u+TfrdsaCKjLt6QKK2wInrHXharlZxvBdC94ljLUR8gz5Ll61PjrPhHMwtbzhmGkIsciwIa
0jxLxT3yFNCtqOniW7u/prGxakdCEMK7thY4qTdE9MyONOt9cbk+OUX8yF7Y7NXKaXh6jjwsZIeE
1sqKHDgSDyEVozKfpghU/zwjyhD8KtNKR6CRD48VWMoU08ZfLyCD/kk9Qyh3uxxbrGmibY0dsAaO
Ag1/C99mPuttlf78mkqEom8Nf1ONx1a1CoabESaANKAjU6Y42IwnBUGrtHb8uK1Lqzfs2Dzto3YZ
R6kNzRQrwvbYP8BP+7DQ7bvI6wbYmOJR7lVOojJgbllGJI4crXusDMaIEpocJQ7wxReLqwMOLZ0n
sSvLreLpnYWM5HlYyeNtKjDkW4N2nrJdnA9CzEHIRnesoIM/temfy//1fv0FPrHOHfHIo+JLgO6u
7iIoy286N7WNrzT9EA0VNtHGTakNjOHS2vsohftRhiR9tZEvYdDPJ99krdcbts2wwP83l5jbR8n+
CK7CVUBR73OBJAjoyz2rmX85Y1q0eSaegeAJ0f13GKuD9d3iIQMoSlHGGof2cfDSB+zshIXFB/1g
sRCev76LM6RnUXxpnib7tw7hl5w2CnhdNjH5+w5LxIA+bUXCJXcsWsuHSgWapoQcBiXJzO3Mvj5q
LkactfG5CtKfScGvjmh3+KljiXo0pO2zgXVw8wG8Ocjr+pbhcACDooEYU/DWSVlUZNCOZhZuLo4v
5FISoYijFcL4wuMXWS/OSMngsrAkZ6FNLlzomtC8tslcJTXptzIcCK2qPQRB2wcHGM8EFF8wKp6E
rQ5jqTBPtSz9tOevCrbYvlRI6DNwqiFAYbicPbkxhnrSU3nlT3tTdvptdSSKkKvVBWAPIixviWJu
gz9SzoxPEuqgbWP3TrHncudf+qwvNBgzJUQOxYSDsniTJfXhi2RSQufzu8aYsdpLaZZwahMJqAFw
rCETU8pCez9NFOGypo/v5jtoRRrzPrONP1/U9gMWWKseDiZTJFEAWT6E8DRjTdinWuzplo+KVVMV
mbYyMOWGMYvtg28mnmfYbf6rToAPSQAYJF93R6A2k/PfnS/cIG2t3zCjvcFZJjr+wlSd5OyyPE6l
peLHdJ7PqETKh1KRisUwnNS/rGr3uJJCl+LBaSwVkma44+h19jkJZqZxWa7k+s8MBZrtqB+npPzn
LNSAZbmvXjhd4IZa9n8s/pQmAycMSJ0jdf1RXjC2GkE8CMEV+A9zaOpJTw6Jgf7pXxMPo81oiSMo
Sg2cIaDCmEbSNRnhg24pFbpFBueveYG82iGT752aElroKRg5c5gFH8906fwap79P1QhG6s2ZgT6F
MXq53xwGCTmgphfqOUZGwJa5ZDd/BcJgOOy38aJLHBjeFsOWCrO5SvnT7beD9maBrW/NDLdkSnbl
ogqL2/SmNA0uEX1ST1/dAJRe3dT606x5dQTRUMyeoZRKQxGZ2YtLTA9rdbUKz819AemYdWg4XWgj
wW5L2LO83soTUfcO6w2czUFceFWd5GsjftAtQ1AZHCc9oV/jIRiRYuPmPrAq0uCMzfOwNcjwAXbf
9KrgehjfZTmhquZE+hd5xOj0gDT7l35fE7ERiLhi/iNDReRU2uehZ2xTplDsoWneETx3mmv6kXkf
Amcy63lGkHP0uTtJH/x1HCpYW1Zorym0WFdCA7geaRFfWdVSp2JJweDCGZcQ4IvTuWY4pbuvGUD/
MvfFTtkR+Wg/0OplYDd0+XkmITw0tf1hyljBxiP8gChyQ5a5HFGtoFQJaGoqdo0YDxIE4M4o8+3h
QRcP9OmjWjBFTdSCt/YGUyjvacJ82oMnpJz8wSTxzIbaF1qAN4W1SuLuMgPxgaVGgONL6dRXvnxL
Wlr9a6tMjjXtxXUV4QnDLzSr79NMPfsjmjLN1Z/aSG9RFkGU/oQ2cTmhRTjsx1Pc9j2jSvS23Wid
TvvJgBjYHZWjNaTygME1rdtQ14i0ZK/1POHhBC9EIKBCYThW8POIyYYsYXkCFYK/heoUQy8tqi7a
zAjT+FERfleIJvBf0r3K111X3OJPP7jJVZM+c03P7Zh7IUrvFtdRQPfQjo3ruwVxcgNtzy8cgBBT
S0KjPZwaxK1PJrsv5Z9mm1BpV8aDJ3Ub4vcpNsEzSkYfX1J5zKHUBFjoYzusBsRJVkLSq/OIYnmB
X0NbaNpcY+t1uhBAMIBr6EUGf1RHugekjkmB3lIUp7w7u8D0G8UDWikoI4MYi+37KXF/LreYLmbY
D5684lnaI/2A9qPgzSlY+mpgIfFzsvWOxjF635HMo48xhf8WFptMlvtvW9ecLQqPpfkA2/I9MeMr
sfEnW+NO/fMZNFJ/caosZ9/SvP+kALk1vV+WI7OHw9kXmfot1prpvGJOsll1vokFWFLSJjgVtHcP
q75H56LcR79A3s30r93kAHGc/xai7Kspi4P0EQOtl4UmzVsFSQqtja0ukQs7zyzzL2SwrsnkTkZe
gn60g2kl0MuNGgMHUX1tj2gXneOS1NJIbDmjqojUPyoeFd0KKCE1G7527A9F80hiwyHGx1V0aLv4
1fU4wDjJV1iO2KUzEswxNMCI+pXqK4p2SU585CDI/l+pjvsupiGsGxETGZLxW58sB4NE93HjZwJk
cbGnZ71LCYHesE7EYp0FT+5jtpVHsvVK9wREhRJZy/Re/NVJGYsZ0q2TrKf0xYzbvAcGpLhaHPYl
eg57s+ZE0vbTSd17YID66h1AXjszL1Y7vvvPiaPjbmaXS4j1bbgSCeRrfQPjIxszBaOd7YPvrOwk
3PqgyCGEaklKspSNnsy7NA7fJGKdPcOFk4FECHHvIx297dm+a85criRQDK3DDsbIqJPnCKyhA6Qv
a68qXd7hsDyO2oIQGitsShbCP+RH+68tN8VUoe3ynTtBvVcnsILN0+M/dElE9lLMBH3uCpTDyi5J
TGyFdD5NnSCm0XQ6SX8F6b+X4aLdOPIxtGFHYi8+YZz5eyrKpYunIwto3gOIdv/rSrUd8GciapPA
DqkbKj5YSCdn+Evn7JS1ettjH24yC24dEtvADsLdIQdOp6LWGKmZq8QWM0D3ocOlPgNIvJ/HpuZn
1IGHiPk3xa/ZVkyN4R5HA/YLBPWVqbNL0oEDzlSZG+siG7VmSy23AozjoCArxlZJwSMBeQxdJOTL
n1aJrvyPtOQ1WLBbS7SGOsEng+lBP6kxc0h+sADA+aXLcv5PMXcL48JCJLbHA0BcDokhu0tB3D/Y
Ahe9cxCno+EBzVmDXEa6gSfW4uyyIFIb6pBfj46Ko82FWXzRSQR5/V1kjUhC7/gX+nCrCm0NLrSx
xCErPeMadyRevQnGxDLlGqq0v5tGzTFHDu4/CUIgmRtInfO7F9cigVaxPWgLBLDdyVDHVDUUCNf3
dsjMa8K6s+6x1H7jGLJC2zuvPpATYCTP+PE/7FvB83u3V1EIsiZoIwhdGwvPuFrE/7vsLJyqw995
9K1q0U7AlLNtOzSwa+4eURRTLYIr7nHbQpFDZo9gvCr3EeNBhysUSRT0u5X53ABFkMN+9f1qZ7SV
MABhuywmtnTtY6MHbN1ft8dBXa/03aRUrDX5Mo+uRIGykc4INuW/vj1M6Cj1H2UZrd072HDSc41Q
pzWQA1vrVlnBdL7S8QCwsXvGk3QQroJjdnuo/7fz81fdPMIoilzEgNnylSry5STQJALr15Yv/vj4
1PyAFwgqRnipmNl9Sho/MFzDPxzzJ62b3HPhub/ruB/HAIKmKLoGMl4/ar8WuLkdlf0L8hjUX3iU
sQ+elnA7C+xbfUYZMNmgmOEYMfmZIMxwPLI9UqqU5okn9aSiv8e6oWPR490Wx79QeeFB8+Ss6RlS
LX7NaqlxZD7c1m32YXXHjUoQfl/T2F4+eQc7SUQeAheVWtuUGDKMoIoaLscRNVNxE/JgmbbdQvXD
Cse0rb+3PLOgk8Yay/b1sGSvSWSFSYZ676D7QJ53GE/uaPEWnhrO5I7NaU8JOnBKftbqqdbtctfv
XHXF+yNUrqtkfnbI2akjw7ZEx4GUGOYXqz1mNsG/RATVaEVM+hARoe29rumpKE6uY0VsCiYWxSVd
gq4QlxPsJkt0DwUTDLF3aTgqYaUd7Glzf/94kWnlF7e7P8yJFnDfCS1Rt9BAn1LqlKzdNmftWQSb
ay+HVub4BH+493a/TQKD87osoVYT1jAeYZtpNWYsLdU+FhYQ6pBTW+Yf8slebSq8xy0lxsxCf5oB
FsjbqV6b3DdrZVaIvXxRQvu9XSXLaT4pdTkX8Qn0IGv4Q1I62YP3EYaJeg8khUX5xZtiwnRIoXxj
hF7rj/axJwPNYY719j563NCDGvNaSiAUU40uw0wOyd7vk6C/jgvbMI7bI4O5tDZ00Fxun4FadKlh
jb0VzLcQ2Woa1/3GjWBlDoAPKDjV3NPLxOPWR4Y//Y2al3HUSitncTrQgTsg9mjF8MuUAetOQvt2
cpOU5M/d1PPlro/+JEhvtYY5OkF9tfv96Aok4HJprpBmh6eLUzhUmWmmaV4gGso2c4WPyKaosjps
HA9Jfdfw05/J3FmNNoioBRDdb7eMQjRF/Gho+MA9XfcRj6+3rjQA7ygFkmlYyNIAXGlkNsGqUpIb
g+sc8WV8gVASYHQgVhYVud12kPoAkoaPxsnyfatIBWIDZ5JfXj2zzBGtZT/kMNzP6omRgmusEkbO
RyiwPTcJOmqQ8D7VlMdUcziOWKad645+SUEIOHGmdsi17mL+8jThDLFm0eHMl22rVFwb8BRAJ7jR
voFNCDSkE/usNjOoBoZyc8SpQ9xQo2cxM99J6rqn6yy4o6mfUam7kxmsCncRW3ZWlePSeW5DLIs0
QrLjQtWuXbO/4ten843X25S9SkaH4wQtUtD0ihSsLNp5ixJpqRJUkbWEosE1cO880VyDjSA9lMe4
9Uv3ShWF049el/LPcI5/Hkl09bUP8dvrukiPQXLT36j1ArizAdCCQjPJLZsWmG4CSwMGYREUsIT4
zzQU0gf9rGqHIYAiJXoHqsuGQhOFKMkrAAPJF53feQHG0PXe1Zyagc+TeOLvkZBWy19ft+K9h08n
CF60LyRKvg6v+RBDBOa3fSrUlRSu8fuVDdh0KJXwKH+iTGuld4UtqNlLmWJOdHRl18kihjaGzKr6
wfsjy7W7tNNqmnpjrl3g4i9cl9cOoADQ4go5jKDU2fd6NsYMiDHDpzd2WA21FoVrStISTbU/HLWt
TqPGHMGQlmbQwe/z1cwUVe1WP8MYS6Y6vMUpLoefu/DwxRH0BoxOgLCDM46384bFtAd06KF1OoDc
38RHdYqksEmasnhtF2BTBYLUCDFvcR6aqh4JqVsklX/kRJuTTh3joEgxiSylbjvr+EKXMC1cwAag
Ngswe5rNh9LhS5uBTTiLr+If1cTvTIIdMljeH99KL+nslPuC87rKbd2t6hjNuxzQjRI+xcP/LmDl
yO9+ydaZR72/HKu42Zs53JAEz8IV9Porui1Xd3tBrNA/xUGhywC66s2i54GLcNapOGrZO0ErVh+k
bjmCS5FMf0bs5KDSvIC2bTkYqgs2LoJf5ATQeqTVrFlR526Xo5nnO07G0SB9fPeF69YYqSXNAs8Z
0KOAKKoW4sgtXEKyxQmBGAF6WO3Zm8tevoOtJEqAWCBNrECTSZkNjOTFsYp25uQC739qigwqiuqY
vOeoUjinN5TG7UvGgaVWboRXJ+QWJTLPuq/rC0tsPqvil54rdp3UVBhOFkGc75AiQAdSB57Kg5fF
Zx1Wx4P1Ihw4Lgu07Hn7BC/wP7mfvV30iW2vBXIxgJDmy5lzfKtSYoSZmv4+gGyf4YahhlljpoB8
OsogpC1FlVY90lFT4DvrD7bKLTuHARk65szjrHx9tyqfYQUQVbZmaeB6xYB4HPakQhPfvviZJ3df
vYxJs0QdCz658WTuRnLuELB4MP83wymwY6CXvHSz5UrCEHd2Ax/RYbb4/kRf4JB80la+ySDM3QwT
wXX2Gg+oGMFt+ze/6H85e0Uj2DToIgGV0RdKQI6bd5GBJc9xJ5G7pEAQy0TGXq2r08pVnq1UnRfo
saYTI3/XceZIQQyE4JlA01tBwXJxXTUMT98s4SY+VGB1L+3/k1PmcMsWf3XeadHXoxE4h+uI5719
vEMKokm0JN+dYRk66WYJIVKjqGBHfwrstiZPkh5qld6GKfflJRcetzrN8yLUCFwWfLJPptEkTE+a
lElhql5hiHpKg7ORM330252+ADhXknDoNEJvfreTJLjCt3szUMTnZEiBPTCSOlqprq3tBveIpfAT
2F8G5e6vzmYrXuHgLYXh8IpvzT6BCNVPiNWdKCIkG9fuSDRhZG4zz2lpd3UoLZbymioUkx93yCDi
pyVhU5jvpfU4TD9HG9JNZhOggD6ahfgRJS4MQpe68ivf7rbRz1odxZCYFo8HEUY9kitK6NJF2ZYZ
MMj39B12sExzp0GBFUJ0DAxbuFPJyl7rTQTHXls9Bynh3p56DWUOimktXPvyToJR5wp/VGnwLwGk
d0LGnESwXsCs62q6eE6uE5adaC/Ceo3KmPCNCXKQfTcVGliEdfqTWsKqCjIltNDI32crEMaMYAkK
PQrjxtDljUTK68GEiOuI8vv+9SYVVaIn09sWgUw1HPM9l1T8VI3Tq8bXMfrqv5g5GDZqBylVINIz
4LEtdqJ7x1FKLjz0EUSD0oAZOKZZZpZ4GqgjOEf7yBWOs0OaMm17IlKRRQwBhPot2VTaGj6aYX2p
lK+EJFqHihRoEzMzF6drgP94rbDO7j4YmpPoq+E+LM5AiEGyQgtdJMz7BZtpwEcVYkcgzWeU93VO
3boZV5/JMTTtRJXgTyoFjcvFNPeAg1gz7D7lmwTeACOPN1kMZa7OdFnQ2pma2+csYnlKonwrTS6g
npGKQ7sLAU2IvKDG5lj8OEN6AS1ndnUrJq+6ZnqbYJS4rYO7l2YE358SiNzxRhnr7k/dV/37BmMP
3tHxyvbDTsB0A6ZkrBOok87W3Kfo9HiQQG/EegQREMJ58tGTZLzOIe3aw0sJDT3gRQe3XnP+k373
/345ktia3GnrL/9ZLaPiywZbJaqL/54XvChBFTFZMplcbewIPy5/wXMOkboUdVPLqeGfMSrVwPgt
TBzcR4Qlzh7CHL7qCbCjKh7p92em4F0zcXGweA2X7h+ABF2I8PzD6IjBK3Sx/zIP9XxkUUWLpBMo
8lkbyxDDHuDF/jx3EqfuGaYO2oNOEx72jJVivo7wSTF0UeNW+yEZkOsQW2qaRZ4Sldrr8s83rXI5
ZYdlnd7enbDIkaOvC/clkU2Mt1QW8YZc/7luQWOpvxIifUx7qWdAy9RkfbB5QakVXD8xoGjlJBe1
pLuKA6+zJOAb2eSf9LiRmnIzsAjZWJN1xMLD9Rc9W0dk16EzrGgRdj3yZDErsXiHPRU0Krg38jXG
QbHkSON7OuGo+fhT4m9Jv89OUNt2VeQwF2ZP0CzEcYnnZPqBGr41PmcMr4PclWVzhNMCJZh2aSqu
GqDlKJa4gNY9iswbP/0FgYL/7zfLVfNnEu4RkQiMmlOim4hlgnySwE/pVsIi29YjlcASC+wjbTN7
wws7wXsAdjIPb9KDpF19bujlVauNDs58ppGorirsppWp+2f/Ybo1v9GIOgHSlAUD1q5w8/Y4qClC
JWAt3++ayUirjPABn4aEa2XZDtHrsgdzx0QY9irjLDCpNpx8Rn7dZmViCc5K54Aq86Xzjz9kikU1
1LknOKSJ3N7+vwOQpOjByiKmVKBw9KoHnsNzbaCT1E2WsRRBXLOIe9nKGkdgcB+2df88YYZgNC7Q
RcvsyDGH+Rgb5xznsL3Hr/WOULck3odx4XhpoisnskFbrU9S5R7wfF/b/nUI2swtvYzutr+DJ9dp
HwTIGsPupvSL9ntiOi/G1XA/hYAFoXUZE50aLFEiZP7RZlpdBDVL2KLGbDsIFYf3UAIWyAFiThzg
Matxi7gUi5mkd905OdWS3yxMncW1B2nAoqqk0E+6A7/bmS6CSxPMh2sXOt/beFiHbBzGyG5Aip+B
083LfMrNH5OUtx9c1ukZB3HQ4i2STt+IwGpQTr21G2wIMFLBFaigvfEjZosohBYBqdaHx+GAFmRA
tKKd0FKV8fhSMUPD9UPeYsnqbPXL3eAzy5vp+MBNIjWFdJCM0mcMi5WGvRqT72w6bahlOIbswdcg
qanpwH18HGoochxLuX+gieiRRwNvxIMdfIGmsc7AW+c3MQseQDsO/gmvHLjNbWIl/kM6tz9mSts+
GOZUV2uRHboVsErhhYFv4PNOQafNHuJi0s70lvaJM3/Ipvef9CDKy7VHfe5MkzPN5J7buJNpleZo
cCzxOfpSGNAaGgV/AjIr6OnYtQ6pGaaXqq+pwysMqC8BCBxVz/zh/CQJaoCrm9GqLHikleJWBkcL
FUdkVqlAVC7/V8xCuKONbwNavNEH/YcXAVJDBpiNUA2EB1LW5jETzxlC/lWeIIUAeXm2/obQwAf7
iK94IQs7rXAH+oI3qfH7/g48Wor2JFTxxzKQcmBETjvX0v+SAzaRm0366DOECQ8wxhYc8Now5fW6
zE2e3+Prhz9cRyy1a8COL0VdqzCtpp+jnNCDjyobH6o2f4o5jJF+ArXEzkMdyc8SgehMBAJyWybE
E9sWUH6Szs5Ced8QMpylbcgtTyeJ1pf/1MOVLoCmX29xLKubLo3MX115bSyv6L8Aja1WBPzgPJ6L
o8Nxe36r9xx6MOl5S0X+ABP3A01/u0pBAnR9f2qmKDq1wSQ3AUwKl6hrrIOFwqu+UsD58Xlq/PG+
o94Oz6flZDZ44RJLX+jNVmLjrMtAqhchqmGJ0cnZNaIM07M4MIkZ4uj2YbPdpQjU571D4Iq64hD0
Phgtab3UAn8y4RSIOhGsfjoe3E9+k9+TXP0+0uRJBitMYG7XzUvxV3wicPx7WIU8CKBNVQ8E12a4
Z16VkHr5H11Qt7hCCHr/Hlk5EXhE8riS4ytGvxhaZjo/5oMUT6ofC5tJ7pgv8Bkob3FIBmD7ule/
I61O3CFE4nsqmaP+9DgdNTvKHOHtabPakx0xQuBvmjWZRZ8nSnUNIeJcyJe7JU0xlWmuT3kYXUgw
KMqV2+sTFNzbdRd0KdRUcfl5adm0DIvEk5iaHZ4lnAb2R0u02EBxvJDFCz6ZqAYEtviFT3a2NYBM
pF0G1CYKv6Jwx7Dr5TVMiGdlQ92yZt01+1zFHhxw6iUMokjfJ8XDkBDJwRE81W7HkkG3QZ5aTMKj
Nt8w0Ck/73+5HErMFH1OStpJNRmQSrUKsFMYZS3blNspfweZhSNNxkRCe09I2dXmVOzl8pto6kRo
1NrwsAPT/ft704gVHZkKALLO/mniCZGMRn7L7ql7yDGnY0ZLuamJ0qAktPU/4k0c0LafwVHKEIqu
UhJ9aN/+LFhQUcuMMeNxuTdo4Ii1nnqhtGTnHYpTsfLrtvJ/qIvwZCGqBYXskLGjA5YpQ7aTAgdq
MzOttIaa/LkCUMoDJ7ONA100UzZ4suNl/Ibbd+RExcper6qACNyukSpoIIZqAbpBMDrzQ2mbsUqN
nSyXEGBNiV7qZbb+EEGXRcwV2A1k1WNOL6ZlxcMRA4TU4MirgLUAZwz0CWj/9DrgUN6calbAm4TO
jIKPCi5P1GA5wJW1/k/HI1cqcY5i9dKEZ9YbQnKi0L6/+Qqnp+/9nwDBs8wtQ/2zNwlxkQZcaof8
weTVNNogU/sf2S3NwlhPxsfKS73pbxBjGTbUdu8q7ggAl9nalNICH5ZmJM2nkkU8LcFXSLv669X6
qndcZHP+FMyE1rgO53xvkcoMWPMCMaM6bewtwel9TCNauPNvUo5eoe7U4Xv5fS9d+V5Y+86Np37v
MboNNmN/JX2LBPaT+pewvIEN0fvwaMJqLNMMyLVHBGxf2ATHQDVSQpqydHbsQsu+rHS2cGAGWHBn
QgfKah95T0CBxNmLEScgHY/S/ICxxM5Uf3rl91FXzHftv9y9Aug+UHRz5DLshpA0KUfMiWysIl7/
NSojtSbO+TCQJKf9LQN0E+5b7ZLZKuqlXcQ42ZDsNUK7J0hCVi7oW2O5Jqb36uIST/nsAGzkgTJd
hKakIgQu1fdii2V/S7j/GqskfE3cM99ZvpHrgNsq5glZOmOiFWh9wJ0UUIcayLnXy6e0HpRoALap
+ev2Flw8BbTAazyinMtyhSa1iiGRAr6H6VJ16R8l23S3g1Tev9UXxwsSvpWH6RBvsUGdAKJQakpM
td3I8onuFzdLqQL0u5v7aUeMoR+5Fl/EuVKr22/lA12QebvnUReTyLNpEfes/uEU/GCzJsbivHT1
SaoyV6nx3dK6PCh9DETzK/nf8GKYDLzIKJ0kVo77zAvmvlGYQPHbBsuj/cbo7OC4D7nPTsI9lsjC
6sDZjxTxwEUvm3GzY2EXjawdkMoXI176u/LHF5F1WVAsRglv5KtIX9ZbkTx3xa8bIt18ZJhjBtG2
8I78cZbOGx1IzLsQXWSNM+5pTwNKNgu1u1cZCVakyW+w5ekiqE1UDxUNMfUYTGH0HwrwQN+/Usdq
YwE1KykVZFln+7Z4xawz+fCHERGRhiQWWO2Blifn4gNkobKyiqvXUp6ETkXdjE0cWD+I4sN/X7To
ALrpDla869hlIBnn+K1hWSnWMfwgaWGtqwQWFHx0Ux8gLctirHCox+GzSgBzK1DMFDoXaugHClha
7rghvtDWdbdT9NwTrK7V/lX3dFzLmW3oyy985O+X3BanX5lKjbW2U7G4G/gG+PyF2Cx30s1sxrbF
qxcHjqojYGlbu3zoAFWnc9FUFmb9Z6ThU0V0Z4bHnVuz40pTHErfyrDqKsK13rusrBbLyRUdf35X
+8ABzawliQWmGw78c31DVJ6JMGGQd32fzn5QGHY4FbVBmVltyAOOVEi4ktumGrmP+n5cpVPXPT0u
f4NzhTVbtuqXIO5pOqqnke0QQ3HyPqvskXUx6nbrNlNU0CDdnSdClQbjiav/br6AKtbojU4F5mUF
uTsU/6wGBhuz3tmjeCd5vOzPuvd4KXSqmYjwx9SXe1uso2fYGtS2kuxqYYywFdM79196knya2gOM
MhO2VWjYMIR21x8Bv00v0321xpydwfosQWQXeMOnDGtNMcHaTrBaAVCHPUFgy2TstD8QO4LrH2db
P6Xg3OAzeaSrlvWrXN/YSAbQ2VlOr8pJsc+/mEthmBfNNJCt1AHkzl81rVpmEmtnJxXAajKtUKL/
wc0pV3dsM2AORwXyP6Q2cM5La7a4CLwACh1kEO3HnXC0xdz6z5Dv0ahjDhjx0mXodvyVucdtcWiv
RnH1ngCu9UNipEEnOroCxbXwC2nd0hroO4iSc5gG4feRmtpcpOanL1V+UK/2qopYCPAzO0hj58o9
BVsl5f+uJxLD6porl+6IScl4/eQHrG+17kq+A6Xtc3S5TSBLFOt9QRsyQjQf4SAeBDi5uWpNCldv
+DJvkilfaRAV8pLrKUuywgIJsRkDcXYrvjuDGuWZNNM3LTQEfqYim5X3qXhZuv2sfs/lXPR/sJww
bA0VnippKHmcts9BEfaEn4LTgkkEQQKOtYxNm8ABXtMFPxW3mm6yBDvGi135mhTSDMKEhJY4SR5h
KLuVhqNVCo4/be4hdqMZVRlqLNKTsNw8cVowfnXG1pV5BfR4VT4CWxNRoDvI06XEA0Mvm/WGpZ/n
F6Bj2Z7Ar8fBYxhxpT8VQ0evpUYzbM8a/5BZ9pZTptvGlE/YFr+HhYes2LMY4QvGiCY4Fo2Xvvmb
oMphjXnH3rcr8abSFUjaZ5y4NQKS6YI9rGJk4+zXsMZWKyyRsOPSQlvNZfQCRIkhTr544cyNKmg8
iL7zTRz1xVGK8FmEt3F1nwUaa/Fx4sfdNsYK0oixTJafWTkppJSd6jhoyQwnNiTRP+jCdH/ys81W
M1JAuxC3VEMNe2pv1hoZSLNDVrD0TdErsm4vOpmPG7SIXbsL2YDO8ZIJSD+AyK5+rmMGW5fpnza8
Ffk5Dp1f1kg1Pkk5Paa/Uwn1PjTnAEanXtdlFhPTgymbMn00xek2oIMRdGlVpdm/NhwbsWGa46Bu
fLXPsnD2CvJ7awtIb5NEi9IZiYyNUJ2bBOprlqI8G6MXI839K7gkobIutCNfEmpnLlADCnqlSS65
fg0pTkq9Kstpr/aO1uemN5BhkZjyHuqp0u0KDXvZzh/GpYfu7WfCIvCObuHt4OEq4uutRZXVVnwa
VISwyFpQGEixOlLtKXayyj2TnUfkov9CXZNtniiy/zvTYjxCQzA+kj7l9/2DQ6wRftbNnMBS6qdk
7aZFn3Zpt5R3oMndWbmMjSp4vkDC7VVNmYugTDdaCamNhWULYvUusI6SomvE8W3YDf4K2N4tFlir
4ReHk7zK77kG4oQ9gmkNO2TJ0XsK9PhO/lOjwvTme67dvGr5j5n8aRO8TUF6SDsnqo2kKw96v67F
ggMniumBQIybRCL+KtHBDFb+As/egGa6rdNOWcoCXj3n9/RIq1u/UZKQudyBGedy8r6aOmoTRV55
ZhbA4YybM6lnB5RkAFmzVY9Npx94+kdFZtuS4E8afAROxi36ml8GL/W3WI7PPlVbGqJ6FYLKlwul
WxIhrO7Z1+ZCsjBIbnPmTWvOTKUBBJ1YRMsFVxMtn3CTSI4mS7GD4ewQgYLOast6bujJh9jHAVVZ
eaJtCWX5MN+xm7frMKpxEo4YxLe23cNt1LOpYxTQ104y4U12PBrDQytT/VklPlYevaOcYvsb3qat
C8C5WiZ7pnHsc6ln+rNXKKspBUFCjH8RhSX+2xbiIE8wdLPgKC+5XnQjBM/cIJESWlNb8+HOyasv
t+rAtjNjd1OLwW4boOLX4AaGtY3BJzPpoDSbC230AV2Rd0EayEBWDjglGETDpY8dfik1yE+3ol01
LZULaUvbrZnMeA7JxY7JJsu0GWvy7ubDPzeh9a9wSrhCxyEJiUR8FcVxmZf4SW5sf9eUeL1T8P7G
mXEdCK8nHws5rBM1VWfCq4hVKKwuXDpQh1Gtjuis+soLosWK9FwJJRlwqlp4PG5PVhulz4hiYgUU
TzsZlNJ6FH2y+z6w9HeZkDOJSHUAmaRjG6NDQH/iwBblQm8YlY13Ff158nUcWMxEOw1KGL6pqsKC
7VQZ42iYlkv1N5aFSIzvr/0Y/IXf/GtU+7jEkhwHzgEV7gL4RDZ8Ys1Yt3s6N1mpz5hMqOsnTfk3
j6YpVONU0HHjfPgPAAtFHUEUAhZc4ZeGvTmGLNjhTTK6dazZlGQstPRtW4PEuFC8uCOofvvvals+
ggKdq8dXasQsX9GoM91gYJxlTX0Do0eyJ2yy+yMWqATWplespt/vL1wdrXCiuAQQsNfMaNysbnA6
beSvbid8a1OMcCF5y1vBE+K5ZZeBVo+YgUpn+LJyp9W+4RaoG5I+RrZcJS+rDiWv73fBzSA/+UUT
lj+QalsY2nOvVg3iD0x73JjmcYSVMwGw+CsgAY6SNryVWDszJ+SmvRu9zmxuHVd0b/GE6WvlmoEH
1hSVB4ZlWToQYQ8lDRFtyI7dU8UWzukoaEtQ/hhUxuNmy5mt80qyEE04huaEAbiQzrcf/XhcKnsC
HsfltHrzRlA6vte8HVA27+ya6xKBbugb/tsyy69qCNT4ac3V+a6PNbPctzs59V5zKTr7O5SzLye+
Rd5jns4hM8pGptQVonBndLj4k7G2zfplOnay+ZGNetDkIX81pvJH8ZGXt4hkePVWeX9Y528TY5rr
LocHrM0cRMClgbpG3bydriouQ8BrqxaC2IuK5+LCWIwHE3AsjTPnF9D31YGxT7OeCeDgvuwtf+Nj
5u7NJI9EHCWYRFnSKzl6iyESuMjmRFt5RE8HnHPin/vREt+hjC1PvfYVO+bwa8iSW/931VfLb+qa
yrckyerOecb1lidBdzD7oMNNMc0NKaZU084/yIOVmfJLpkplv8qIf4837k8e8oZ9GA5EZLYTOZuy
tcM7QWvDKxWixnxQIkjxt8esltrSg8wxAkzvSlmjAsZmLOp6FJ3YmBRJ43xukiWBn/cS69D5c1v4
j90fMqszIKIBd6jG8+b4pMTNf/7OTygr1FF0V2qusDoWQFbjmv+rWanGkzMKgb767YPzDTNmmCpn
JpCGmtsCjprMVw3M0w7R03EUq8PsIC3IS+bMZ+cIKNcsslzSRF4Bdhe+PGY9UcUND3XETvGF+HuA
l2puoNGGImy4RuaAs3p9RngkBU8nSh/ru0Ent8j4BstDAoM+I7Zk1Tce5w6RWgURhrkLHpdXefFq
raNblcoq3FjysNA3UtXgXJQ7Xt+hHP0lkqKQrQEYf3/JU4xg+P0poE7dQMBLPc9KPWsj5ka4Ki7O
Vy8x8RGj2gJftzcwHQvhq2Rf+uBgGHXZtQaldZxYKA5HkzRDH+gjrd6n6J5ILCBBvuYDP7Cky6tX
/s7K63elzzQxgXXU3yzi+0Nas3iG3BWMZPOpnW34lFqKzFZ0NKT0DOsVQgDc2iOfDxwHEHryqTpx
sXwvSQA5wIrtqNSYzUd2+De5F+psPq3OK928Km5xKifF6vxFhma8qNAJkxoGudAze6QxzmI+akkd
0Qls/bLuTM2u9velfTo9TVrk++aEi10RqL0mHpV9G0dAFr/BnX7op+nektj2QPs/RjefKR5gF/UY
i0dbGFYjRvk73khap67EQIXSGyxxpVAOwvkjiJwaFT2rohESWFZPPSw6woXJcTXgUTXBb5nh9/Yc
ONuevbdIU5a/PkafJGE8FmvaEe4aUiAqy8knzk33Gk9Wxaq2hs9IAFHWFlfg8sr8HotcvPyWI3NU
HzinhMNIsZVAwGKalmbWyVv5zOJ7qe5GR3vQBWireTDQu/sjuzePlF6fx7m5+AubBWCN1ua9+nHL
vFyiiMB0x1nlhRGQvY6OcBez1OL0PfdgzV7MkI7dQssBd4EMXmD2ILLxHWkJtTHG7V0CfCkxP0E7
PeF5JkVPmgqpee1IFP++UageXkC3x0k2WoANo2ZnjQk4trLqHaalIxH0+M7Y1Fj+SlK+7Y3DJMUB
YlFcxBzXkfKmqR2txk1RwOn11BN3tGu+YRKhDxsfCiRPe6AMgjk4Se2Bxd94omeFMZjYJa0ZF5g7
xd9pEZkd8W1YjE0tmP6vTYeWj0m7a6CCdPZSIpJQELQm27TKX2YN0f5p9JksNyXknRHEO0K7xnQB
Qps0Gecw7X+BMd8FSJnLunuUsYsNjnPYwn3vJ3DUu0Ku7SuEOA0CtQe6l9IiEwbkO91Rgcu+G2ci
ytIhRfvd6bExcWsvNMC/g++dRHCW+tfnqNSHsLDHfu0IbTvjpQYD2oxPMi2hmQ0XnSNpyue0PbfP
yfIG7HkAHPmQ6Uf71N8fHk2sVab77cYrNjNxnD0nrgagF8PpqI7lDdNhxNyXRkwUQKAuO2CtAeKF
HabC6EGLiYgAxLQ/EFiIVx2VtBWYQaBixCjNBLe0deoVXh/8APAGlQ42GPxJqZPRnmPCh2vqcnVc
BsuLvIsxWbhWJOs5evFJvcb1xV+uFdJKc6jHlnNmxXtEAV8HfuElhJmthRaCd0TjkQmCtDuRkW3s
5g7jF5juxBuCw+1LdmSYeh/vH9q94asemvgJJulG4/muh1d80iD87f41N2YYR61RYyE2222hAmba
bxhbarHfk/mVvi+GWSqEjGNS0uOhhUTvJB0dw4ZdlkpTEL8yVupzqqrFInU5NbcmVoHtPWM2rQ/J
18ah3MJDXHv8tBZm9ylg10TfMiB9HIXgm/YOH+3/vl0DrBgHly5lOppxTKpn8BB3qLuj/o0KvZcm
AWcyScqW2qyfvxBfawbJSvDIzDU9n6ehs+C16bgOHW8Opf4M4UPfFeh33YekGKYjZuudJ18PMslO
bsQ4zYzKUUW0SO56cRX6wwUH8p7RNd80oDCkGE9ESuZCJXuEPdH1jVY6Komz4OaUMglJ7GAF8r0v
DJuXQ5z89i/0091itu7hJUFWIfcEkhXSWKEhGYH1gkoIiFXJ11OZgsZ3hMU3yP/lK1UUe6h5J1LX
h8SYVM0/fwxIbgjuvg2WIA5GBCyuH2PtVgAGcgJ16sw/N6LYdtuRHxGRIzIUl2PMho8TZqikGaQ3
DAW548DzH5S8JHNDgrkKjAsladTgt0+obzP7IVUif6Wm7aqbm84G1lLnOY4mucm6saKwnntLt4Oa
VgK4gD4OV/K8NREo5yQNW2E+tfQmDKE1eGsvgSGZlw/NJ1sQupmnY1QeNfAj8XgEkNATGvAH2RPc
be7iqu6DhGpajl54lCtaGV6+rAsClAvIvLfx7i8eblbIgDv6FIdrUcwq49mVxAGSZPcECPwt89yL
R/CvDVSXDcsXHcFAXFYRtjpMnpyldKirJBvdAN58+8QdA6vfzZ7iNFzRVh8c7wwQCFg3x5d2dEFW
lqlosFs7cW2V5IqGAlkJt7ztViblqG3c6OI9TALCkrfKUSkBDC2hGreBKfkfNGYt2Sl1FLbg7C8L
/OpFnwrRUZSbj2pGimlo/0sLeSiYYitFAAz/eKTDqgGUc3KyiIgCsqKScdbtgzkG0pfw+V+sZS7e
n8OQu3SDrTxK5XjQOiOq8bp2VfJ572J4slw0Q1vak7Dm75oeXB5b1skFy2W7P1Crkc1VJezpc2+u
PfkjlbFgORRSYYbYV5w2dWLTFgeNqm3FwYU+7+zHfTlCi60xW9RPhnTOS+KC5wuHyUUfaPlKZE+j
eZvYOJp9edeGAFlxH+Ht2eJnXZMud2n3/pOw1EBk+cO7E0FFXR+6WF3lQ07f9w1WZJ7xAAGeEtyl
CzEotW2JOhazmzejZEGv1UHaoSO7D3dtUmDEth084+JD8WR4FjzvwpSHk1QSNZBySfmMrxMUmguV
4XVq4vvc8AaHu6SwZt+rzDP8Ubuw+vOGofw/9BvD+KN+jZgursNcu0gmnI8DWzgKZTfLbR8nZusg
8UE/BPFtjFKVi+OprcaX56/ObE61mkWm7FyrDhGzPqsZUOOSKbsDvQx2DWax7FR5NDxsLJKnvnmC
weca3TGMss2CpzwBVTKu2OZXWh/De5XQuN3dg0eVk9b+31eVqQ4QnvivXwinFR1AfFosudKqyflK
GOknHNRLUyHwPxnn/XZOz1ji0yzYcYKNmG4GeamDTyJIyvgjS4Jp0ZGQNkVvtAwR7KdUPs+uZHtw
tktSKsDXEYjuQ8iG5P62DgjT1qCB8fezefIkx85iYQZ/+fnAKgzrrQU3DVg3RL8aPB3BLxb0AIcN
CFYhzrK0HPoAFHaOKpf0F+97h1nd8hKsApm7N6SlvKxyRgjLy3E8oustrNOeV3ZJ/yn/q3mKJjmS
iPpfaV6P0aOEFkZizCpcONZTSb9Air7E8LUkQVtLhGa/4UCnYJV4IHIo9f5hraDEGnIu98QaRuxG
lMhJN/7Xdu+hNRb0dVQ0RQ5Q2GgzoOFqHNy8UNEkjdOIp21IXwdyK0wFuVN+XgF4uQRTYYLV/IuJ
hsAw9mCmLjVTYxgFHKizKiEI/zP3I7yD5HdI3jXCLGmaHuEGGpLjOWZqvsia/G4sirCSufe44fzq
k+XXcuHEKN9oByYQtL7bWnVtlrqvozycDAPjpdi5X/NynZnb8hobhl5V8NhrrS3qGRCC85RA7ADT
1LhG1YcVC+q0Qca1GJg4GEEJqpa0n2dOi8FQXYT1afhvCIT6aqjpQVGxNgFAuZGF01reLqNZSTRt
zpZv1mWFLrLVQAVRiZ+YdIO6M2kuDpSnzcb4Rk9mQn3ftox0zzAtcdrpeEqWPmgVPQ+pILCM4W09
Vx+dF7sKvIgltGL/tutQOD9Ox0YNbtwzJsAomjM2qb9tqLc9heuIPAXzaC3oMvWelIpot6W/SAqs
7ltjHI8mD/PWskWemx8731DA1Ts02dHmHI2hz25d69+AbeRi1vYjrLUkng7h1gYU6SKirejOZMpV
NZNA0GeRrx0Ip+ex0TAkVgK08aTvp/bjhhM3DyQNdXuFZjjmx4N9qc5umsIXoqZncu5coXhMBqne
oAXbwSupl/GM2Kzx3cIBJDmHsTSWnq36IRjY/9tvqYPxIVrrdqXGbgUCvtmEPvSJe2YPSitBJvtF
vyVss4cjrfadyO78qjHrczV9LiY5eMAd39MociLB6IdmFwfVbrlz9RABnl6ksYcztJsjWE2ITvHf
zyc/zVg9YUqq3OPtkA4luWoZzODPRk8XDUvKAe86tO9OgH2m5UgkqeI7MSumhopnfeXtKICu6mD9
7EGuJlQvY2FbSkzOl3MxcDN64psdpzCGDjaBWduCPvW/AiuIx8cgLMw/EmxJvf3T4/4yOkLTH1Jy
TX6D21EYuQK59WkmTZ4n8kzksQitMsQKh726Vbnb6SdvBLjvKqTmDmeahh8xAQa57teCA35sYVgR
mMqlosg0I4QZSHeUBQ/xbJrbJuz9WqI1aIWK8GFM09SA1du3X6dIQ/hpJhX1a98fsq/Y6tW2robd
epZnMBFBD92vo/j1hnDDOVA+hyqaYdKj2KsRsXdRcZBvqJ3ofz7EhqCzftAq5wcEPZdf9o/wZeVO
OUnyN9MSGVKLQoc4+tFBc/lBt8+vZRTFiZy31GzWu7vYwc023pWksBflHO24xQZWKAVeJGA9Vsp/
4AJzEzL7oa/iKV00UCtLNpa0hnpxgWA26zkKo3GQsgZpsclE0qPCfG4jMRrwWebEPUdn67Q+FFNW
kZtIq5V+54X6itgzcgk6UWt2ptVYS0/rGFdUv3kkbKCstPEIrYcP6XRjTjRf5RIZwkCAw72wCB+p
J8AzZIKZFN4C4lYpEFCtUQFKz29W8c9kttPTZDomhI66aQYI7lz2kCCVlGn9lSC6xdIIBb2G7ql0
7+6GVUl2KjeaB5qpbEqnvjYu7WUuW0XEuPeR8ObOB1XZEwlo8g5gcDdQ0v3asQjfwpBa+NsJVnMN
AmOcLdMwK4NJuUqNZGeAlww5blyMlC9e+gXNZOMNGHO8CY32Cf6rrQLhv22Lr0T/3x0PRiBMK7NC
+s1MH3WLHZBZKwUk+0ubhdS0ZpVrThgh9vJqH54270tfjjweqQEnp5MPffmlpHbbWmzVHZDwugGu
fFVIr4b/pkt5hVl86Pei1n46G64u2WavgE4xInzaDwY2svK0PvzjTAZrO8KXYUrAnFvOfmrl0Xl0
FtLEmuJaQv6HpqnZQ9/TReux3/BPqSWSqyzhP+1aVoPaI7SnbbeDwEC1MzKcDLykQSczXjWFYvS2
G8eVlziz/DZex6oCP2IaMwVItDaprerqYCOZ3kisjaqvCzO5w7FrQ0zVFH+mQ35zBjhlF3RB94nE
HHq2ustO7hKCeZcov3D/YEdYuRs2HBugXfumVggFwZsLUqL2twnhW6T7Kdg80gKf7bWN/F0sAwQn
MQIfedoCFOUKdZHxkAC5QxUEOjK5n5PlBVaf7VBbJQ0YPcS3nX5orpXv77rr3IbH1jJSxnHAdIA5
eWyNxTiA0Kj+S6Umug8qbc05jhEOjppKhfEnTge2Bwz0d8A8tMHicnEijsuPKmXi2AN2dbZEPb4j
n2D1bfXqPPH1m8D1et3DqPa0ZdI3cN4QRPYJza6PfiRapqJdwtB+tId794iXZtN5Tz1eDRfCiGe0
MZcnQkUb8WpQK8zArui1eWSbYo9rR2xzj7aRWLhUkc+G8N5QrAyuEVwHTnCFjScsVxxkxYz/Bv3K
M6yZiOk22by32L0hR1D3uytrq99nGkhuiZQsjZiPyZNIrpfcgQPEOS3np1bLFwGPoTBPsRw+kn1h
Pd2U6Wyc8iEjYEQdsQJU58LF0afRAj6Z4oPNtigyScXiMgvbmCeZ4qGXWfN1AdgoAzMp3gU6zaPT
G2XzOZH6s/T+KtvR5/ktF7YEXlgCPQgQtYKjugAqu2ZRfY4DwjBnSANKxqBbyO7GjQEf7h8EsqaA
aKWcknMinLMDEziYQeLXxdJuMVPsIssKu8Ao3DlntK7gUiIdHX8anjQiUDS0K80B/Srf3yWXx/Oo
IUp0ayskl9sYmSDU1unitFbDN9CtDJ3OCHuwEc9++u+1a7groqmGojFCY9ZeTB/d+yInL380L4ZT
MEQJNchwe5EJpR/d6sibKYMsnVDiaKQBWdkbnTGTKZnPhE7fITfNGx0goXtwhB8vFdz/87qc32uS
uHBNcVs2AjhCfcJA/V+rln2bPMu/hDXrQyfa+f7SFzTBXwI/UvqikIr8GRjFIRY4bZhp2RZ2lg4V
pi67XOOVyoclnq/zgK8FEmiBCAXrk/JC/2FfH/znLQ2g9uQOXh82P8/ugetN7oVX15sieAcbqC+8
vluiBin357ice+pgSZjZ08Q5BROv8ZsWUu1uk4aEPZpCiVlfOgH35kae5loM8F+GD7ec0zACg81U
+y181yYrytvVAX3kH2rYQ1TLbwvK80jnEwNbTOrd8CA7IB6hoe9XMfRyhwQgNN7hU0wn225P8Y9u
NoNkgWS6nPdqw2uM8ImjZ1Hk7tibi0CEq/hiptgKa4zoktYs4kQp1U9ruM6i57yZGCXq62kTschB
Ehdyt837GJnSertbrquNdCV4LCGOEFkJjsFW0PAf2YHjKaQ5NXnwFqHjnTvCu5LgNQyAl5jVYRIu
g5U2u55wEXJCrdwZN/5RqG8cefso0d9DHP3cKSLC1qnwdWlbiY7fdRI+PR1j2wjkumP38vtbizEe
2tiDiOx7WTG76khax0CeZ662J0MIap0yO2dmi7BUtfr/yg2pAvSO2uM2fb0z/Bs9mVb3ETrG2Egm
GjejXef/0UVY8pqLCEAweiJoWvQIBh1BCh2onOke4lppKQ7I2HlqtmgYHRoMzxOB2Axu7ofppzZv
nr8EPeGawuqr9ssl3eL29+x7bZPNSfA+lG/mJR9D444c3E1UdYJyKTwAPBlSEyK33i+6cFDzl8/y
cmU6/S3V079GXa8VxTIn2r3aPB62RlhjBg4AE5OcV9CMp8U1GVkzga5Q3/gJaIFyCL45aVxuQwr+
bA2oyq84/MB0L0QswI74f1+JhrWEBegwuDGX4IPcRZYQvG/YNghyfu2v0d/hw/27NZku5w7mh96n
1oNRMRGyi15dSUuzrugEV7Mo6g94LFNQvu7WNjgki4jU4cvxyeLocgWBgsuE98u0I+9FFKOEYCw3
+L5Z3zbj8g3sfuzf/NDmoJx9XisevMybWhpZ908QyN32DbP1huiRZMw9mlAUnc0YxQ8nHMB6O4ds
Qg0I2Y34gdYZctsH2AoFr5J8SLhI/B7BON35smiVGTxLdGJfzV/Yd5yhS7obaEwBUMp2tG5mvlfk
TheA7/2m70/wyCSQ8Hmc34D1/7hKvLWyxMC4873vGl5+DmHM1AfYfggAoXVgfycfXLOskv2GIpf/
G7/ZQw8SffGj3s1cOubFZBetyYRGd4UivNqiwCQSWXJ8Blj6xGc5+5pUkd36Uk8Li/NVS96FhEMM
Xb7dMptHpfzvUh572Fc2Cd11ERfnunjt8mIbFHYUvOZSIwHkn84DGil480ZfpXLJyhIxjZigwhU5
lqTkLxFjsC3DPuuh3VOCgxG/EWzHOAxkUo7V0u3PsE++pILnQJpmYFdiHcbvOmn3+FnZZGC+wONO
gFTAo/GO+57aRj4zyzb72W1JFwXu9NQP+TQ+XTWuTVD8XhteH8au52CCqI3VPXiQcggWlVgg6XNd
2cZ/Vz9/umYrWt7DtWsKggBC0T/nbyg7qj1kWp9uBUDqunbcQ2xTl+RwTvlbpNJ7U0dvbFOLl/4/
BFwbUNwAqeV9bVUoEKxetJ3bxmDhElxqZVayLMbBGCYULfqdaM+m11TXGX2dOrvlylkZ/Rzwce6M
02FI09iZFUYhqSzpH73L0wveiujZbgHNX6lXkiYTHqiH3f/m9+QP4U0V32wf25QoKrA9e24Jfxd+
9BVzXml8qJd/c6M0iHZ7duu8KNsTjudzB3cCL+XwLXnPw+lkFIHD/V6wD/Muma3SEVcKEPMzfp2z
GYQZFYq1RzbxGzlTC2IoI7zGKP0+5vZozuIcKX+LfKBQJGUPiDczikBh0xZ6QmIOGYrdV0bcm1WD
8WRBbdIQT3tRM5QD+bxdx/niIrerkcGKlZSilZ9GOnu8HVubmazi3e8Vp2Gd1ppVTHhW32oCYkL4
WU9M/s3gW5xMbQPKXvjPztsoYKMLOLwgc3HcPo2IvwHYCy0XQ6ZV5nzCyzIT4lcwiuEClhVu0VZ8
jdz8fnOjL/S3ZY0PjiG/+HlAuuRBPTbH3W53e3ymZwW5SWpFqCkeP8vjvrYWSnJUQErXbGJy2fT9
fNPhcfKSpNvvlnA5xSOMa8aj1pPzBFGAkzwv4D69tnabV30umQtfMHQjm4mjCbSsVbL3b2+4REnc
MHL56vB1p41j99ELKxbUB9umw6Kv/UqqEzvUeifloqRknSDnb0MbGK/YHsPop7nXLOBRzI/xei5d
8jBZvWhTE8s4jrBJg0txX/3ok9z88J14mWaxmVb77jdwAKph5ygbT8Nh+ss66Gkj7OoIDb+rAvP8
rzbkkgOY/I98sLILkOf93m4NrolQj3qPsstAV3psiaF5CH3v8Eyuzc36eK/uDf1mYlby/Emiwfkk
GSxARfbJzk2QrmRW7iESnRYwNZLumc3dvmLHzKFUxAm6quEHpTenoRJFBthvokfsYP22I1dq5Mwu
o9xeP+A7PZpI7ybqlWmkMmTc0eiaupOZqQKvt2GhCH748VhlzCOn25vtAwnp4uwNqlrH59ZvM0p5
+40kOZOrFlMp03asd/+lcfs5m9+t1NoqLCmekFtZhArJ2zq+jr4duTdQzvP1Ez/F/pr1Y5NRKTxB
eSISSO2qwAtHZMjshNEWx72MCyNDiLYQOXvRMkOu3UPeTuwq/Rd0vJxnlNPc7o9yQlwDf1I/HC9w
kru8qcjgAQZnR5cMdifoEZlgXrGFcHrU3OrkgyikkoA0Pl0UX9exs8bEuPxCG8SYEILECrbdd//u
obON3lqxJztvwhYiqXo6lpQVujzrJvvkB0sGQXXLAbde/uUdJtjltud8TUfBEarfTxLJQQzZ20bZ
pOk6maJgThq/VGzjEvOQo05Xr7IM7cVP5XM69e5EFWw1MLnxEhF8u3R7v1OabOdLV4VYATli0Yq4
kfBs/7D0KYZL8F5Bl6DCi+YHCaeP1DBxKQZrgF5ZfAr/ajAbkZcphjy/RzXdUeOYamcC2tbhylJo
UCW8hRoOzBJo2BkhTEBvNyFW06Ef/G0tWSmZ+AtTSE+2V43R7UF0b/NDKo4F2jZNycODwmEO0DUP
2xtFppK1T8V/9o19vKR6do2B0JToM/Y49nhYB8iZknvXgfG0/RabACqkjMzd/s0IJVDMxAoto62E
LtrwPx2S/UyGVwNOrwMcpfwrHz5HJBHwMAwXWWstXBcysAixTLKO1Nj5AM7vDzHOZuGVbzT9J/EH
xv08S8EVDhUIkTk+RFY2tVbAd2hOdi7/M0NT8rLcmXBZxcSRqlro7jmbUF1nefIN7DhVsUfAK6rS
FSR0vb2O6oBf6yQVPtn6S97gE7a9VTP2cm01b3yXeBhaa+PdZqmAaLFI3us9xb+dBq8KacLJis6a
nx0CUL618ZGUozoCnrmnQAvgNJ0HOhoa6THZDTulcJ3uZ4vRuB4+fp8ErwisOoW+g5GGol3ad1VL
8lyrZmVbEcj/s6EI8H3XrdtIqKch/r4cRzfZseG4khtIOwei4n0Ic/8Yp95LIFyH1D+0d1Fh+PrH
WATEz0wOWQ89GuiW2s28CkXXpyDKrcEr/L8/Qf5POEyQ8kiPBYT+cNtby/ljCjLCklT2n1JAcCl+
pUZjATF++HaVH1W7OylinRa1S6n9myJMsYmUVV4eNyVE2oBChNQrPiHuXfQQS0KWosvPGaZn+ovv
mzEnI+y8KD8dRWHL66zrftg/CTqM70FPuWYViYTUH0+cxvcyNeljp3+b1hiChO8a6VWoxb5OUXtx
nnJiLx7cUsyhZ/zw9ecUeldUGqmMDKTvcwmOuPJHQBYzw1PoGwNKyJRhquNiuRtGvVg69Oaz1Grs
uPLKVgPlyTS+B+nP8Gk0YQhVzz07dRwArEJGQCbee5xGGacKbRYMxUQbhiELXxl5TwNBByB8Q/db
i6Yd8BL00ZAh2o8Rt8zx1Sl9DBF4jpvEnr8t+vJ1L4mnwFJL5GQCDj20F4Rx4jRbYUzxYi3UzSVn
yt/uTzFgG4KCdsrbAu6YcOUbpbMUuoLTUFf/RUVDIIbJLXBVJb8DSvclZ1mcDXrkzd6hkwSPPezw
kvwf79xiQykCjf5D9E71pHKrYAgsVoSFO1i544OhRuqdFxWt51SxiNzBdZuOVZsoJR/QPGVBBn5w
po3//2D2Mt13ackgQi6bZFNHFr+57oDGyV7lUS5n357BBMVXMoRJExIg8gOdjs7S11FhC27hB5K3
N0VBkHxXnd9Da5nDEzDSUskngtJ8bpSz0kYvfJiDjXzzRaevAHsQLt5yTc1tdVzB0N36NaSJ7Vg4
MMyCUYOfdL46S7eegTn8TcMyqjUiXRs6K9SteqaZRnel9zztfAGicyB7katunCE0mBZ4Gu8oOyBi
dqTVzG4dk0MQ1xUL34bJBr5rSna+LSJ8xwWC5kH6mv0BftlvQOlbNlAzJ2Wcf8pww2nSm0PEUDQu
ehQD47mljA6j0lKx+5KpL3zXdNM4bRGfaF3SPxWK8DvQmEU7E+Jf5V5xLkMjH/71T3evhpP1eodw
0AyUdFnzhhupIMHvjlAu1/n5L94CDLDOci7oH9AdulZZ8K3Jnc1PASKwNJXbQfXRHZnaiRKE16zE
EmGAqTUjlcDpTMZwVk3OrJvvjOvpdZOkCwDYQTNt2w4bSYRyv4NgsKlHdfpEk9nIp9fX0laupqmE
aD60Na9QcS0ss/3AkVedDDMUu+/dws4RzT5MOoJ/NCfXLoKzelqPIMGx/xDG8BEu/3QwF4h3IZda
v0U1h1LDkJpN1tVexZcOqlBvXWRpqFUz4WvWSviEcIHjOnnoi/Th8gsYQ2lOGV0+xiQv1efLOgBp
sPs/qAwrvSQlXSYt8wScMFYX+cwG/FEnJrI12HR7qc7JgGCbu2KnHinVOWZDcQ8YZqCjmcy2zJeo
c+2UEm3YRvbcOShLG4oJaAAA44GaPRUad9FLIDlb1F4LX289GHdq5HFz+n2qdOt9/0HKlozM7oLZ
PdoMNY4tJ7F8Z+fqlj3bn753og4PwVPl+M80M/JWC6RPBche2BvQ7EKjIAKrwqlUT8Iox0XZ9v+7
e9GtGny+0bRkJFVfP5+wwQsprVRQUF6pXqThoso8Z6R4ZPVSEoj/FIMdIi2ZljFVzXJtwCAz4lHk
EyLC2ILEVgMzruYQvLVD/bZm8BuDcP+iggDeH85l6ePNIjzBtCb+f5UPlG66utcbIQ/YaTwWFOpf
1+urY7k37x5zDCVnoTXfPgal8lJLgW+qTW/6LvaVFt7GuXqpQEYKqtXYUmsx5uWNk3sOblzWWC71
lEPqgS7KCaUTrm3FSo0mQUFoG5Fn84ah+9kQpVnSe3fSdNeSLw8vX4U1ssOjFp+Cti4owxzX1P04
W9DeCpE/1MSs+S0cOsFBYvkpDWh3yoLCw43qfLhsnrCQWnWPezh4j1fduf3oGFxcqtdqb06Q2tZ9
Gj5popkQHp4o5vTywpj7p8uSCyaoY7cBNUbLdgiqWYxZblu+8WNdQ4+wg3jH9LDCVD6TKB6cPIHq
f1FeY+4Z2qIC0V1fynNgd8sq7dIib8pfo2ZZKvOr53yte6yD002qXyt54QQZ0tGiLX03Ne8GGaI2
9/SGPUe114Eb1sNUYF5Ekm/Hek03T55WhNZDaEHmAx/YfQozo/Y2r4e543IFWh+5SkzbUgdamkIS
1+i/B1TygpJuM5iAzn1VYs29EQ7Yww+Oq290OKRpDaDPXHXIM87jmTKeTeOQJH0uimkRNVAvr40A
ipAW67SAj7OgB7ZoP/Kg/9b5YrU0X5E8Sey6t+SV4OI+yzI7i3Xdf2aKDAoniieURkOqkOs6yYK1
U8Hd1nFC9x1bYWYPs3I1FZQNUh/AS4aiihjMVK0CzvGCpznDec5AeY1rbSkTCEkPBxw4rVydLpWU
lzHUS9sV8nVcSP87Bvc2uS1I2BxwkGmSnZUNawQC52+TEfS//0GrTNXp8w/uCwuhwt7TJVSZUsoH
NCGrQKxA+zHMZd92DgRg+AItK0qnNQAVkJhTOdgnffN0cLifxrYEGVnxtV4A9PSFacYKgXv8bpxv
1hYvTCWHGB7JiI8Wj/2lQJC6QJD3pJOFNZCTw3PEbgP5CU9CMidlu46/VtOoLZitDaHVV0ABObt/
mM5FKhUBQ9ddFS7yYPR8smCy0IxtHG/4RQsNgyFsdqXIs+mhDrcrxX4WosGBSDurRbQ/DWlyhkFl
N0uj/HirvLwP1+JP5+Y4F8RqMBetojfDMrpSlB4YItkXm5MwCwra0WK6F61K8SJ3qWb4iI19tCUp
7ckdTnJ7VPTfhdMM9AM9zksLZGW917QcaIX91a7IP48cYfa1jXJe9OFRbFmoZJjkhFOfW+oAmVpz
ycPBq/q1tU9C26Uu+7kA/hzQPJflJGAr+EldXpaEjgsEDXlnRA9h2Y7im326peO4w+pvSN6+cnRv
ane643E+xgLlDnfy5KvPWS+LAjSZw2jEs5EjgFtJSnEyHza4UlVFqQpCtkI6CrMs8Ds05lYXjNZI
2G0dkxZtuctdeRKSw0X06bvvW1jiaeJLRhQt3s6wYXBtxsJfMmCyT9rvtmT1UVk0THZmpxPa+SzA
4aPDDrpAwp3ohI7XllKK99PNaSSDnyF4rSlf7ntd4n4nlWQzZq/o8PlHK0kYCA9N1/zpgt2uWu31
M5t0IIPhAK1sNbw5gZjgptZs0EOGxF2id+Iqk+7eGmTRTOv7eoNjsDLu8r3M2nayIaYUUcXRCMg3
KBxBgUMJe+CRtIZ/HLs4YBOrUgJqsm06WYeryynoIW4ALwBhvRzck5ddx0DiEbeyVObRL4m2jk2v
AEM4PAPgneFel+maHCByfZBqQUp1BqCTCPA9BeoKDk//jRGYCCEGEOfb3/FoTmZ7IjyOpn4AScJR
ztbFgN9T528QKJux2AcdwJKLB4TD2bHOjhokowc6m6N43RtxXIYcCai1lkXN8ePiYcprmZHJ/FSw
CCLxumQX1vNlpsDXdmEIU/Br4POQE30o/zaBt9FXdB3oO23kxtQTISSOCjPe6DIUbMLBDTakjfKr
77EjIFZ9lmPlcse+zOWda8rK85GVWqpj9coDRNdmE4N97kuCvZenccyPkkzkmT0g06eZ8RfzOR2g
tpa4wIH867j8HVLLI/3R/D7Zi4Uj/fQgavHf2mz3v0k1M9eU+ooGPm44s+GRhkZD5Mc2jB2Ufo1T
L9EGLiA3ZmHjv866LzyivTwDCMDp2czkZuxfdKu2uVE1yVPTzWvKjpg/VTyqoOVvmMx0D7GL8L60
ADs/8Fb32q4kPOSILiOo0Ge1Rg2LoPW0Uiqp6pTdlFgRJan7ifKxyhZiTL99fe6qIMQonJoHVOO9
D8WeiG70FUNO5qGGSHp/+8zD7WnpzdUwBEXZl5IwjrkivIjnKwCVmKhG1WQXpf7GcNeYnqb3x3bZ
70oQN8aQVlsp1fRR+QyzCDjC/XHYoV2Fy4Alph4GFK7FjdgJG+tSVEgoCVU0zQ6JsQGBE0FRQr3e
0UyBPoptdzWoojWIih7EEbYSJ3o+FYOVmXgLk9MR7aTBJKFRU+CUNNKoEVsOlbaNsZPgdiSkEW6C
4w9pFetLIQ/u74n0mKZ1YjU41FoB40SJ/RVWny8XcBkmf8aF6/s4BSDrjZ0a4NOdAXO2zkATWKFv
dr1PCDK42rDbQ4ePJOFW47Lr8J28rP2T2oZ2xmIk2Wx6fUS0fPUuA0ibCbH2yKF6LVznZMPVZYOR
ylBdsi3BaJKDabnvUKM0gGfV7Ka5hzWOjba2T5yGxGRnyO0rHAy8XqgJVmZ2uUkm7mzZ4v4SgrDf
K25IzQtD3gp7go8rCv+RYV/1C0s7acd2F3xM0J/PlM7hFeBMbBaj814XRX9j0dAN9vKn/kO9Lzef
P+hTWRjSXWIfCfSePQjz0HXDXXedr4b/3TGLjeUw9WEwG+ksZjOqbgSELUyceqR/UmOcJagBnub5
MuAanEqTVDn8GMrXDvr3bnzi/WfIjUXG7S3KnzvDc0irb+xuWJsLtWVOxihXIAyB0xFPz5A8SR7Z
NZX3JHRgTXYC+v4yNqr9ThW8KeSR0bWX+03aCceqIcGOMdUalJPKjghpBsZuI/6O4msn63x+Ji9t
xNk05xMA8zBi9Z/dB783dNM0Z5YE93Xqk5+GIjWStGR0djbA+SxdQ2RhOLGzcKLvja84rzjkJRMm
ICXSVKjjfjVHd6BL3OP1drIkwM2jQ74pKnAmH5h07KhIiLFvHbXTycYWs4hRhB4AHMLL5dSafErB
sZom8w42+WAJH6yRB7v8Q2uN7Fm+wAjq2zmbKefc5S8gZr7sSwrXR2dCep0DSkigtVduOzCdH3Zo
ox+5flAw7hsd0Vyx6kUDyuPcOYjTff0Jj41jQTKMI8tWZcgtWnIx6pvoJGwRaGLE2rsQVxsN/YSr
qj+0HdlpP2LmTmcdYWglORwWq9kRTBwfADeSjdGUMrnjf+O1z++DXsxQIVZoCmaTf0p5NDI9Sw92
B3XnTpZf8SZvoe+90vInpHnKs2+AEm58WNxSsWNpRMob9knE/rVwxKRfZ0nII1sKZ0La0AC0pfJW
fikzZ8BdNbeocmxA1Jyd4QmDSd7GHsvupwqGqmAy0KN6mt7TDimBbvDUoEcxAy7jqvue7wj+GWJz
34Lcesjcu/RIDF84I1dl1qF5UlWRcLe1cq9dz9MfS7pzSqikzLWv1A5JBdIg/+o1O7P1181hnRGo
bJk19fhqoYl0jt/eKKXs3aoJrKP9IMNbKOdRp/9UKVQCtVAsDL3leQiCpApBbaCynjTA7qRH7E4K
QF0VQZxYS5bki8iqt7VVSfP3fVnBd+MAYeUSQWx7RRaOL89ryYy8Le2i0P0x3y5AFeuolP3VTEFA
yG6BPEGLdY22si7gfjcpYxN3Hel7rKij8T+MvgLTlvwhnuBnRK/MdxLPW0rtfw73Z+L8YOo3yiwL
hpJUgjH9tJPGbziuIPFkMmhWk4Q7F7N5KoWWgzZqU+KgWYnaIoOXpsV0AioyfK3FFGtomXt5/QjJ
+wH1pqxJjOuJf9yywhrw6ClNSW5b/V33R5cOynSV85uLIvcpNI+mJfB385ySQGAv3s1Cx3CIALei
KdtMHBSXNhlVXspZsHNewrt7EI8G9F3krAdAsVBkkuvh+p0WDjl+hEi4MT5D4BNaJUEGDtF2PKzl
hpUTkEd9CWkyswaE7bPdx3+c6XMwydCaEHfwSPUAw/kuno3jL/EdBhC/mNRXJU6cmhXz1eSYo6Rc
iWcfLYkkW8BOpZhjCS14RyZUIMCqWq6r6kXL0XGV3PdRBS1TRs6JiKu47UIpOcJONeBkQ2nAmlCq
8v+b8+TMPgPl/14Ryq5QNHLiV4O4phdX675iklCNKnmk66KsmCYgYkivEZn5YSv0zZnhpFZz7XAv
d4QQ+SQgSSLGsIHZskJ8JKd8V7JRbvU+JH23MZ96uHZWhnDQP/S33IaKAdiN9a12UhyybydE5Oa+
5gIKjQoeoqTnLYGGNnkhcJJPYBC6BEahRzCk9tNspYQzdi5B5ZECy7JiqaYZkS/ntqIBbxYVP+8G
Wuw79pIZrevtt3OXtAABxQ/ZTXlf3sGmsh9UAIS/i//5IllimprH+nN64bizfJH47fmqR07S6GXI
KAx11SPiOgTw0Bo4e8uKxby9mkJFDBf8a1v+tlC9nbGg6nWJ9x5Js4aL6zwbtZaMDq/vLDKq0VDI
QWhgpVql0428JfjRU7mkoi1prWhjeSR0F625um0HSzRkaUDZZ0r5q/BmBVY4nGoYwr5wEE9Wni5s
wXZlJ/lM3CfSgEPMzU1qEC4QMM9I0G3gFof6a0tN6XmgtFi/z44VDzEoKHnU1hxRuofZ3mr8UxKZ
bx9EwPRM9HMku9rlmO7A5Yo2hC+uBE5Wf7vIWQbU5LNjkKCu/A1Jej+MUYH0hl28iQ7dPGah5oxK
i7BR9jTlCIAk90IzEsD9Ztq2wE0eXgEUMQva1rb+C6XZSMU8fx+uxGPkM8rrf6TjcgXLwgTqPDzE
nBToU5ftF9wEWmslSJVy29DagANt8UqqrqSf5VxZ36WRZqUJynZta+JIUYDfPTdj8utn2xxe2Sfv
+v8s76lx5DfGuZO5bE53n1PVFu7PQrCLg7/JmnUEtBIvb/gGvPIPA+6rOpAPCKok0IHdtXcfIvRG
5W/5nFC2OcfMqNOqOZPcJ6nRnDk6jtTD15L9EnbZeGwRgU4g8BpA6aigfxxsL9EL/jj7H1wcPmBa
ut0j1xXTeoBc+uPed670XeU75bm9l6BpkfahOene6WjFx3urCrYmA4ApQkmQOanbFXXMLJxfuxFi
2gg4UtbYrHSVpEq5HIc/ThJaq9gFxsVsOTiynB2Q/CZUloEKHoA9cRO7hhllaFjw7IhQiuc8RKm9
SjycEilQi7FlOQp/mQ0tzCeUbXID34lrAhLfOpwntoh5jrJgdekA7XcA5Oq5D6qFx/+cO6rzTxx2
/fErvlb3iEeQQeycAAtXELGaIJucMlG9GyZ1apaqsUesCBxWahH86/FONhUIQ8WRfGV/3NjKKweM
8YYtbb+THUSJUvZbv9DjaN3U6fY1GBgqqUdTzcYq/gkh4xI7vcv8q8zf5ONevjFbA4x2UAKtGNmZ
sE46A+EK6m4mlQw1KQvTJL5vAy1Blc2VLINP13Se4WLZPDDVLR2FdZE9p+LZfSC7r6Wei8uEzxfE
TX5VL93rr+lYsXdjTaPuKuijHPyL2WqUvWJCTihaDfddeY444/+wFIF7q4Qzkii60AifA6WXmjPI
9hghp+VacGVxx75Lrp920LRYeh/wfO9tkYYNjLqlNLNUD/5mfn8P5wYtHIqyA7XM5F6RALq1jqXN
4ZqoHtaO7VwZE+i/oyCiPMAYWcWVVBhfZ6sAxf5csIdWOHTeXZuJHSJHsbvs6mCkUywnpkuvK/3J
vGeVONzaE1uPTGxrxWaHUD8sby8ERw40OF37dms3MT0I82oVf45B5yAFEBEluj4IJpWYRJgZLxAX
UJIsJWKDITH0QDBMzN4rd/ffVXnzO1W4sl97R5kZ2fFbDs/DBsKeg/keS6zeGWVwhkUvfcGO4ZJW
jD62cdCHGrP1CjyUN+TPkzdXVPp90jdbvAuqi0GOza/oSgCty9vpzvB6n/O2dVDxXZlPjLlXHyAo
AZuDCwDWiA/PJ8FuWvWeZWbJYEO03W9J8G3SchbGRTr5t2dvltFngDjKyPfjvK1YZ6iQ6fTJagmj
abfv+IAZh3qqLgtXmuQjb2/pzTYIAcOw21ihSsanS+FXGoqaLMDMOdGjJeRwYXdX91jSGgofDQgh
LMnPdvXj/b8z3IvsQ7ilglJ2b/t+u0KAp83DkoV0bpQFpNL5Mauyh9sTrOaYMHZ9HQAay9z/H3ec
/yQ87sMIXl3MQEm2FztzzKJzCzwqwKzUlpUUzeo/Sr36TgT91aeN8xXK0z+Hi8A6l0FQFXS5l1mY
DvR8gdn8gBVa/IvgRpyd9hD6hoheRhhidZCdnyJHK10/Ev2BujOexpCPX3RIIkkIsXy6l+XtXG47
2IEYKqG6gs7P6FGmdl021npvBsHHwc+RAOO4QrkZe49xi++L5QnIKLo5MpfwcH36QC1hR9J1aiq3
ZWddE3AowtYHxrSnqoaNWRN0CbqXr49BOvc7mXIPNWziKg+bE3lWziWdqzwhbZ5TPJXpb/TM8137
qukrmwbbF/twhgx2YKA1BfWFxRSVEjLFdG9onuXMFFz7KMTi1OcO0ro6HwWqhQWIkX9m4fHXC4YG
NrCi/muO+LxWoFHg9Y4wOepcStzwyXMoqceeklEctOD3VQzgqHF6wSjpSUYbFgfCQJEm4tMkmGs6
UFYyepv9jDTeDOULIQkF9yMastYqpHik3wrMZoPzymPZbAUIovshB6Wm1ZovWMZauqKTIyVIu7//
JfOyps0htCOcNmSenQVyUy8k0KiGnezf7wg0IOoteZKC9dE2+p3DhIEzQ49eRgdNk0F1xYV5bryt
cGKcSkRwFxUIydelD73Q9SACNewTGQvgaB6L9em9IsSof8e4/W1+Dz0d9Ji8GuS6/GHeaPqCvFAc
+YsfPTfks4+G79bKUUXwhBsRFOcywHfFIq3MhuImGDHLBSDsj6DwYOeEngjjr9RB9mRpHZrzj9UJ
xl8bAgAcwAbnXzaA/XlBGHIpzX+NexdnPuyX0VeiThVsIjPZ9DOOo09eRahJaW1wrMnsdVwLfQUE
CCqygdO9DMwqC0zgcD26Oa1I/FTQTN/TuxkaOcIE/oHGjWI1PC/sKWQXaFTztObIP9wu0gs6s1xJ
Blb61lo927pamWIOKUjnLqoevrBVYHLEt1yhRmRTUTppgYQaAtETla4cgt5PNeTEmgOfEXTs+/IK
bD5Li8XMDODypWH+lLPbHpXPw3E87fC1z51MdUH6sZTUl2uN1Sk00MwhX7l81VPJA8NLw0nnF9aT
umdXdaiX6UMQE5uBd9o32ZnRUdzVXS+TeEOEhxLXKettzwdb3uOe+1YmQeNk7NprWo8eTBYKsWk8
aAUhr3KIsVjALfTNcsd0NVqWzhpIYrfY36kUcYsrxShQ8ndDiFooP0rWRoCPjbQRwKWr5Jj2Lq8B
iu36FXMwY/EbF5hoXQK5yvyKqzdH+KL2mnkVJgNyRJUUsC9ygaI5A1rezWowv3qRk9lLiHLcNbiK
u5+gCNDmqE9mRh1sIe7dUYViViXX7nr3t5r47ALiL/yo8cyQPJ9qwuKzC0/E+QRWmS4pXt/VmeE7
LRrrMB1j18xYwbFZ8xV4LCP/qhIvi8s+ADfKEs74r5I9iSDxiowSHUNUgTVvXv3MAwEKFY6F1D1c
jpwbRKuWRm7MbJUJwsLiIjPvm0r5EcQNtBrsJ3wqtH9XCNEcdZ2HA5W8eDhZ4CwHFCzjUhLOZOsw
BgqIkGVwjk8YTbMpGVVte1XBpFcC0B8CD50Iyx34KhdbTF1QGbtmpimPL6S86DV6/nhI4Yiq77lw
UL/y6TBePBsGV6R5DAv9wRzVfychDGZe5HDPY6KQtvcuZ2adI5I0thV7Vyatwrfiifo5MEu3L7Ow
f7LPJqALE+sSqOF+OtORPgPkb5kk0gChd8OEFEF4iWfOyOWOmeONsbYRFJv/SdfxP1nX2g/2P/9x
7ymIPReyFJmMmgOKwnTcOwY9Z1ZiIA1TeNaW07nNW0Gv7ubi53KX8usCXjh6mCWj67IO4Xro1//N
pCiiND2Q49dnxo1aoCPphf4wE5IH+3Zbczy39dBjR3MGonetrIdcAroaMhs25l7qjdMJO6ZRO9xB
8w8t/FaBc/ww4TUzSk66vGjwLUJu0ORY2FSqMpG0GA6/osUH8/QmWpIiUwcEjjzeF3X3VWDwg4XE
hZlV/08FGwu2R2reZgqK90+qrhQjvJVw6MJVhFNYUMLfC2ZwfLrnITcczNkieU2tKmYBtKfvddDq
WHaUB1hSu/kSXdiNcJ2zmcnI4GHP+xZwRjtYsAUMydacAxm5cZx+aWIEUewJhRkan93AAkGgbuYu
E6mVakrJNf5/12CCkGZHKdAIYI8ix88Dp0m7QHQOe+eyTchehFkwgcQ6Oxvj3nS72U3FDlXwHfaY
8+QhiKHVKBRfMJTqGlvpRBAO+0DHgAO8bIyHVOx2yQJMsd9/hxTUo1L44ap2KIL76CI1/oz5BcT1
12ewmZ5k88GLPa767XK6gu2lj/fvXW/zuVbxW8hn56eXd6/VSmkRWc/nA7l2khkxoEVyc7RQerie
3UiBAiq0TRvv3SDnSot0O/eVsEEvBqwTfp/pi9p/rlOFyr2gX9z6yiJmFjzlgqZ18EeGbIF8qYTr
fcaotJVyOZl+2ZHpKWefECbKn7NUO9Euyfrq+qh5rHDd/GM2sQwI4Jti7E7XejhsBLQp1E+QXXeX
1TIRY8xP7S/pCCb85/CAfzTIkd1Zn604f+UOwjpATaJW1kwU3F/LH+BFO/rzabe9ptXoz7X610Gi
WZsoadSkO2VWaw6e2TG83HWZYpFTjcVIiiqzvbnt9MYMkITJWoC0eeQJpEMYKuo7jnPJScFjoWjl
lqyCtT+t3ZzKxadtN+I/NLCVz8Yvu8n7rMznKirUocuo+Q9cEdKNR0VpNMCeSFo8irXWi7OFrr9F
kzpKQgTJlG3L0wL6cbTywjEL2Qg7/o7G90aMkL8bShYMThBgEtFzSdfGSdQBfPQyNzyYMqGC/HOZ
twzcbg7Wr0okPg6Mtn3mZ0o17kydDg+SU7/c3eQt0cHE0XXABmwu8REmdEMvf4cbU4Z3WiOFFFTP
APfETjCxk9Nj2siUBmgaJz6y9ttLv+YfMBZKC8Mj397/dLlfzI1cEW+1YueLz2EtlTDX1CS72W3I
omjKWaQCEJES7+/0JbTdyfzSyLRB7dRu55RRaFh+z7enZ7OJnQnHjYcl8F6Bkw5wNphFwihsWYbV
mEggLmh+NF5m+xxoCL0jrHcp5YBRx6lVKBq1jjgwVxu7SSm1xy+vhiT26sVZsXlcTjSGtS3hHWI0
NAYYYOH32JeBGp9LXcAzXyWmwtAP7G5TQIAFZMsIquXPQyAEYrlQaAkJuxUe9BGFhO3z+xhJtnS/
uA+YLAJX7tGmSVRMuJ9rzB0Kgv9xFvpnjSagXCdPFyLQgolOXCvlkFkw+2K0a2yOMHaTyCJZcKLC
DtcKqMfd2oL7NRhH+vRHgv8zqbB8GUcW5YKt29B1qYxi7sqqUATeiMSwYl+SbZ/u8nJ6n5PfKw8W
c98dQtwjcSwjgqyr7p8jLnAXAsGZtRQBHvIbgyO3fuFEpg86HeW5lYELeJI0Z4P8noS2Ml/O5mdI
/0OyG001PYeOIRaSpakgu+KtsKbelav9h3PA0szSWdJBwgzUifpK0bTCQAmXHgv9+rJcWFz1T4Wz
B1iYwKmtyHesU1OSjAJCq3B+xvvpUhP95V46AtXUWnjJz/u8Wzcvv3/rZig1TmFp2em2gXKxL0Hi
i0CQTTbcCp9j5D8Mm8krjHZPibuxMP2h+qJ6WQ+rLW+Id95OdMBgzBn0fE+fTF72ywrOmCmzHBG+
O7HvzSW3TbJ5SUtXvdYdJ1r0qKYXRIf0H2SyMRzAh9n9T6RKD8yIUXctfoXEq0/3mkb0Dh3OoCsh
gpVW5GJMD/jfTthO9EIxmRRaU+4WIglTylEmU/Xm1f9af2ylCqQ4bGERxobKIZP8Nlr37e9a2HcQ
ztEaQkcN3B2XNLq/iuyYLs3KMPjH9E/oCU6/x2oM/Y78EnbLGEZGGCIrjzWGKsgQJcf0ive3NpL0
J0lMLs1v1+6g+kuQ8oLNrl6Wgau0a/0IPusM8YvTp8GkFRFKupdMC0pLz09+oXJDDgcgLDLfRjsJ
JCv+MgVwtNW026Up/CchyKSbERRPQ/nwWRHNvxQYQ0j9a8QhT9bn/MSLsNiNWuXoXRdkapts6l0G
u17mCfS7q9tB3FblV06kG3RS3+MPGud06x+u5Hhv1R8llbrs2oxbNrbUtJpO55/sRGtr+HcjRHDO
tpUvWkeEq/2cVmQn3FC4StFmpfc3HkBK5+SpD06MLJK2tVfoJxPDTCEWGc5taVXDbItpWpkchYjD
4dz/DCoOnmDhgBpg5eDYR66vB18O6eiFBnrwcheSByRX0SyYXioneoswoW85myjGlej7QZ8C0nxa
bJFHmb4SqVqVIlbC6WnBBNJh+AAht+7PqmSqBuqAgnJ6icPt665HFB6OLta7r3lzlcVas2Ql/dhX
3QzxZ2ZyI9H2PXRQq4zwErr11j1CinDTuMq7WwR0UPiLq2L1FX3stTqJRfg1QJihTQ3wKGVmyIfH
JAIesxdrQ/NaMv4n4hOVrqMPbHiU++gWgWjQogHb4qyEYzrQcQaH+/+xtYRjqa3vyioREz39LX3o
injzhtuF5lRRUep83D4T8jBkcGK36G9X3xSM6nafJF5+XZMV/J6YrKx04Knuv4yQF7PPBz/pGap1
HPwlXCRqg1gfDGLQ/2x9RsAR4fhHznFrvpyLagrgy6JGJqfY7N60tgF1FNamAq3YuvhRhUSJrnzA
NKm3Z91DR1O+9635FVU9FA+BaNfCmSXuvBlfSD/t1ZD2ATMevbZXZc1zcoFmtLhMXPwrKtjF/LjV
C5HEvo9bXGKGZ454yI5nd8UzCYNvCR5+36xLx665RR2Dv1q6UEClNKPnBwu9B2WezVUi70ulQcd9
5gx8t6cyccZnfpMrKVlxpQ+IpHxpjdk98ZvzuENPRoP+UIYiSi6DQFXVidaa12LN4kql3xJeC0qn
Rgv/kDWUHFzzYDExzA8QzhcOoI7vp5YWrI5l6AI0no1y8a/iKIr0GAn26Cw6qSQt7q9e2SIxYLrL
dm1o0qdC5sai3HrQk07hqYxjhzgossvdK+z8uLsNSj7ImIRGcpZhZt4VSb1PNNTwJ6yZuuxs3viZ
ni8Bb+QVN4pc8IdWLUXMDwQ4rpevkm0xqSoHvXsFWKByaK/7S2J+SzCgSDU/NKzhACcNNb/Vvlau
05RH+XBG//9wPO0lAIH6x2P2dQuhhbCBppiWTFjFILNeN3b8wJZ4U80lC5b3m+eyz5IJvGE3As43
fy9LHXZ06v4DvMI34uidV2HylumMaRMtKuSLQ/LDgGszys5tmrfxL+96AHntnmqZgUzTbV5/V9Op
M72uydG+9IqlD0GqIHA0MBbBy7b5F6k7W8eJ04SXZzFn+HQvOP6HVwqceLfqcIFSEWU+CcB2nTuW
JSgesw5CxRC1ZhfEu3GV3lPzp5+QOEsjAvUo8auBhcR0A7f6JDKPi9h4hx/yRO+FQZ5ubBWvclqi
FmyKj0mJwmL7GMmCS6aojEQ/ov57I/TAXsqEdR/F16SNVj46q0lNvrZuuTOD1v1M9Pe7whKpPLA7
DSXH6Uu88kcLnPBaJcwASs5OxINakRF+pUjL8hXcoEvTtAlsZInx43ayPdzIkbl29/HJJxDtz0wV
Kq9e1SrBEL4uA0tvAS+u6++6nOjUSwcGvYJn99LVxzR4lnhs9nn3cYeIUiP1vJP0uSdkzbej5SOP
vZaZT0srpnsLqAWXEIIUB9Mlp3BhGh6rBHs+mX0X26vxMlKKDRqbBrCtIasS0z3suNXTalGgWrpY
xXj7Nx3rkTIkAThRiDAGGPg04c7IZvKHOdOEQm9ei2oNJZUAEDmTanDsI9buvmR+VPVfjkoK14pb
OkIyFDAd3yaDmjtmxRCaChss8jQmx3J8FP5tp3eWXp2vOg5BpXKeYP3nFqjV7qpP+48dgmHJopFb
9OVHHyVYJ7cCoIEOXAbNhNpR3VyNxVEvMoDMFUqrYD01pt28QbVU5+Z/tabumgU5T9adiR8fnZdW
O48I5Ds/NHXLJ8cOHPG/iZa6m0lpHPTicT8Zp0A2K0GZM8tIow581dXfZVy76XrHk5Pa+xY6NF2I
6LVrS32C+u0+2oJnVD0+70mPfxSBlKb/ZxSgJfIis4vUbTzH+69D8+zO7+TUn1hJiGu/70B2akST
dWc10Tupesll7tho42WylfaNuaxnx0gBhhrH1C0LEcsKrkdVPgFjKHlZk6Uuwvjf7VFPzp8vPRDl
LI8qh57U/CH7MkGgAr0CB3vcDHPSpg68IgBdJS8BOfclDv66oY8g8ZzSIZDGdMPMN/4HfuI8W+0W
8rmKttFkeMQ5oS9QskBVNAvqVlnlorWpjt5oyhQ8OT6DtITYOgI6Eb3Np+pfuZnrdcJDCO8IIHS8
mGWZ22oUVVRKS2Anui2XRvz00q49R6G1dcck9P4RKxjc3j9ZjgRHjxirxOD7+sq9oNNmqKocEa6P
OaPD5Ce7RyZi3bDQMEBYYNZduFxTkfPgJa5Wy4f4SNYHmPVLDSpM2LREOn7QVN821YG0WOCB3A9G
ND85pbk8QAs0efk2jmVsn3NzNhQVYl83K2U5HvOumTBpm1aIFJxQ5G2w813ozRJSqVjWKPERnqqF
tE00ukSgXydAu32tRnhgWdk8CD/jlcxg0xIYgNVZuxY72llRRLuhNSbrdnuSRkTZu5DpT42x+897
cb4Q+hPpvD/eLG6xHTKr6AUPzGH7tsdgukes9wxmr8/BCxLYZkZwrwtaUIq+XqxouMdCOo5svwT2
r0ooUoXVbhi3dmXNO3RWfO2/rQCkXxPJauzpXaizwKnBB7nMckH0os6VHTqiyhcMGUzF92NeAjSK
+1yn7qNXVCiI/N0nqE84ETyHqjDAtSgsMWlZIFDC6udMfv/MXOzh+tDsXag3CPTZsWJttYW/t1Z/
x2D/IBji9x2vjZmmWMvOINKX8o64r6fwX2dxlmr4aIV4NTyuVabmJgA4fWielRMIkWs0ANyJtfym
IhEWJ70WuSUIVMDfWgV40eK1qrbWle4Sg9NtylRLiDPX3OVx2RUdeaRIQSvAL1b5ZlJtopVJAU1b
wT8fJexxizn4HP6ozE6bQCV8dzXSltwVIyLrB3futyrBnfHioD94IXc5HtnXmPvNuKVP+yIoPdbJ
TQaHsl+v17Ue/ouBuKOUTSFxgrFgF5cmNqUP618IoKJ/J0euge0J3gbfX2xHdTjgnol5dzq0Hfn5
0y2i7y/HqvnovmthiM/zTsdqH39olPk0v31CTr7cjCVHAc4XKiPqY/rKnmRBcYCubnoK9noEDL8W
Qf387NLseTL0GY5H/BvFOyimWFHFVwJ1m/MkI/n4/fFEbNL9cbKpk86nE7grj+GSnccGG8GkGobM
2hp47VGVJ13UEVQsNzwS0SjhdVh8gWnPL87geDD3cGwrOJD+2zOP4344yGaeqHbAyPBTGFzJ+5Oe
ut3e3APPZ+9UqGJEep7jGeOsBfbygwIaq/ZtwdCCv3HL2d/ewCnkauHNntxnE4uj2oILNAT2xr/j
NRZJDQ3Odns5jCEh4fNV2SGV9SqsIVvXOw8WOit5rRMNvDqoRcgUqDJoDLhjslVUi2ttoQ9TVLuw
d+PODOattVPZzGjLASb95OckX5vvcnBj+oH7FtNXYkrZkYOVJtpMCcO4AnBziOrNDulFAyL/8QO4
H7qGVtB39l0QJh8zX2ALxGa0fM/mtctYuGuwkMxuhzUlOVb/7f6pBd5reqThqLI8CyvvJNRHd36u
S7SZMnp2xEPqb2Ok8ONtC0nGZ5CC+TA+pVHrCNzPKVVWM6Dt79OVpHyOM2ZPfMBee253iM+gHGFW
/tSt6Vqq9+LU6I2HbjOWffmacN9t3oOU51ltm3J/Sz6RVbFMielwui31/UwEsZHAGlNHkYrgE00V
DvNSk+mtI4Sjq6QL0rGhsgDlP57W+QOPn2srjhMqcU954CeUyy7d7rBxMkDYo1ha0enbIS9ifFnd
J0VvGaGHed1cmTF8huUlBl5w5nZTu6IwPn898JF0JCIhB+X7K5j3j7wdL9oqxDegwr6gt6T+tUxh
Sb54yaovTM0LI0Do8ToD0QmQd7rgu3VyKiVECx0oWWAyat9JsS7r1TYJD9wEIHrV4tmh4JzTSwSg
5rjOZ5S607lsi35PwhvhV408HlSYmILWZg3Nw4Ks0xsy096WytkkiArsJk9v2iI0Oeb8C/d6U0oT
GWWyUm37LKI9a5g5Gz0RW40l944kjCEb2nRVnwVvamZ/ig6h0CWw7qrsJcUykBK6cuTxQRGhiKvd
Uxe1+N1XpZ7aVN/3qQHpP86ddF8xVYflazTIBsh0o1h8Iz1BAL7IWVpYUbt2Xi8hkbx6sSizC1LE
xTCHvkvV/t+7sXfUurH4N/py4pqkpW9zeABeZjS4cO+5eTZSil8as4WIqIGAyKXMk5RuHHjmMxqm
z2Ky1weQxHEQ4bei++uiBSXdFn06LtCYbHc/sWc1yj+xTIDX1bUVaqzHJoicOZMIQf1d+841D5GW
QOZldbo8O2ntnfDagWFGw2HjT0paCn1EXoM3XEMe6devj8FSvTPuk34Plrq0ZqftlbADhqwpRK/5
c2B4b1V+wjTizvfrMsluGVKzLQZSLWlEE/RquU73NybE7FGLwSF5fTdM1EzK09bAxZWv5XHVx1CZ
OBG0/KReDXkFs+Ua//WpzGzhsdoLd99HuK6zuDE4FwGvgO2v4GZ26kVyxz1wV0S+LbkQgF7a5dt2
Eh8lz7DsUJ3J4MtWgZ3t3YZ5DPTx9mDxDaebkyGWupvj6rAhfGMiS4mot85Jkr9F5YIAgi9ybvD+
CxA5Pq1HyvWBp4pcZHcusviSOQ3VvCsFQ4JooOeYPCmAwggl1yJ5ly0J7gGZHDqJkSSjtIkHB0QB
qffgKYQ9adY4e8vPLKbq5yStMhZDeytoBWgVAi/B1Vh/+Lb0vI6WZb1ucPnHNdM5+A0IXX1+I95+
zUZ05z4omy8u8IB2iEtgarx6HzkxYOTCskeYULXRrbfQOFF8dNH6RveUVyMFdFL3rTvgO1YY2oEP
ZLt2N5hvAz34P7j94mfr90/qLWO0sMy3rVm5f2Kv4S80kj4U1OVFQFDx1e1F4+xJulHTZIN6o8nS
YCXmlAqiW5QgIvKo1vXab32RA5sF4R6dtX6Oilku/Gy7yyZPPByPFUmyp/UismtVnOIY282gwUPH
Z7oBXuYWsrF3Tjm5hR1aW/0JtKXnbs0ZkBUJr2ST/ISbEZbUfMunHd+ibCa4XpO3K46iy4agiyHg
WEhxDILa9uiGGp/rYiH6NV8/khZHOaX4GPjtqLI776ZFDYbLVGMOWqACpNJwMByISBS34+7Ug+H1
4TZPgCXHTqh1nxhPqOGCM1F6GeDcUVc2GnODEStGB6IQmU82EzxYAm6hfJQ/U0OJ5rogAlTLCIsY
tFk8hb3NpCUXYHD0vNxtDZgbU8EpiGhozi9sFhZbXUjNe6xMh7DlUUN5uT+60CdPkdWT0AkI0+JS
vVujLzwx74NEU3jIfuEudVvVYTmq/POTs1CnfFMp+RYrcXhkvU3GWmBNsAQWoxeV9BdowyTFOYzq
l2lD2kJtiTULkYMFLBdh3cL5oIcCC0em5QC6PaQt7WwTsvk/j+of6PEnUj4rssa2FkQoc2lxSs+f
RPgCfU9hJsD6sck66jCqXnxTri63DqSZRv6zObLK74iDBszA2HzOdIjfZu0wmXF9abZjqPftK4pc
ASC2z+HMvLtK1SXaiXGJesghdeISbJT9J0xrvN9d31eac9tOBNKlCMK+rd3f//pwep2JuVtHg1wt
smgGpWsgFi4o15H4IYIj2kuHYgMBlwRU83wkcnzSJTE/3yhzKvZoVsj35vU20HZxUyj0vHCGYNV7
mklc5seGnv2B4TtLrNiinUB80HpM1R7DTOD0AMrZkZmCkMWEsw08wBkSjOyalf8oUUhgOHgapjA2
zTZS/ABME+HIzb0n8W5CWMLaNbl7DvELNKalVEQAKGLrz1ikZO+rdnB5C9rnJikK9ITPWNiIPxy4
JUeDwsYk9wIFdmPFHvaVHNf3Ln5GNy6+wHnVzw1HWOStha5NA9S3BlgJ7h3kKJlPjowJlqBPypHA
+FF+2Fy4XH86yWgEkQAVVXP5QI8AyZImXOXQW+kCSE3QdlF1mLRMlxXdWDFChQx6xy4PKfA8pPej
VJS2/wH8012L1W3QwjBrQh68xLby529iGj8tO3t+qVX3MTUXuTgx4MAcR4Y30lqOG4/IeWTSJOaz
R/DIQ0e4YG/xCzQDBi1vT0wGXXd/bE2cQTM89KAXuYGA/HcxdK0GadKKHnA/fS0DOvBj3PhWVhDV
QnksMXM7LT/1NBy4J3kSK9bgUGRO/Sy/oG/r60TxgAa48S0+HizJ5vexorRcHGP4/eAoNUaR2svo
indpJWo8OYII5B3BE24XEwDXhuEEELMQa/X4lh1wkU6t5s+enck0Yr+jNHcKMrPYBDzQDmrDuWwc
6EsUtXXflkB2fFeMZnx+OPMI2724RRI4RqjE1EsJhp52J2KwS05bUrMiirbinnIIwrhcc71Rb00p
lHhSKQNV0UwfXu3wZDTMzGG69oKNx+/hMbToL1V2Krb9QYyACJxjlKfRjJIS3MGHQeOZEc88L04z
6Ti0Fnaz3KlW0GoERlXIJLhX0ASCYOAWytE3LU9/dRh4GRUnHSvkoJ0+/YTMqSaTCJB6sUClaI/5
Xo8O1+M+m4hWu9/BFzXTMRzaDTSCm/tsdZ6V2AchU0OuvmWtZ2iP2eiTb43dVdIlh+n6Cy5fKPX7
GT9Er/ylYxRV3NM2wzICc+fSOHw2Yf9Ig1nrCAP+QJ9wNV2EQUf6bvJQ1Q6jJAFpxokJUpm/b29N
nX9LlSVTDlH9Q9vHFOt32uX3cnEGt38DBnA0mgRd87BxYBqmKhgucCl0fUjd/glDR/r42bc6Y9BH
7YJ8KXjccSKl98tLCpp72URecucCPAoYgSPmVN+SCpVJAx2nbuKdSsLVyDkeXIVRWRcaFb6bBH2f
mNOEVKq2LIIuVccUdazvYgbJJwEZuWZoJeYQLPV4fNGWVAFpdTK7YOeQ6q3rAJUeX9rw9jov/Qjf
iG0ScyKlll0mWLR6aQ3AtZR5goMGIzErMXjvHz8SI/ZMXjY7Wbq6+ozd+LXAB+CbjufwsrtERszn
BL01q70mQqh3xN+4b66f/TTt+U6XPv2D4osC2KT/kn0pxYUEx6bGpiv1wj4c2FVEzP7loBMI1RQC
/SSmym+MNbl6+I7HYDHu2x7AF0WhDwm1keTTFWSJML0i1OC1Mo1SNAQAgQCR4+Xd7FhrnpWj1cJv
u84r0qAmlGfrCqcSUa7BJAXMoOaaULDOtuUI1BbcBW5ptDtfde/Q7Dp8mVcAjczyquDJKHqPWmW7
lArbOKJoItZsRp7tvDPEmlcn79Mkqqmme+oBrG8TtQwt6OhOpMgK+U7ATN5YOz2NF/X6r0yI57Ik
OBHC9ryU22d6mkTNk/wUOyVKdVL6ATH3AmuMe3xm+DHRNWMn0rJXFbZRMwYn+eaH97urcvE09Os2
K/KhNz5IOI0BqdwWvqzX7DmM6vaBQTO+d5FoZCgMwFZKfjQtaFLJ+QjU9LexaM55lF9T35Uu636m
0Q4FWpf5DSG6aQcECM4h9OuALVo8yVmKkLCGOfxNvXnB9+kGAMYf1enWlWKILx0hD2XugBNZU/jp
gHcBhN+aJ+lkpPwwR9NKnUE3IkkZZctUfALxETF9eNRlV5fsGu0sMBmYsJ97qjS2cfIh3j205s1h
kRJuPeH8ttRMhRLzLqEc+fiPvVUs78pA3bp5FTFwEZyGD92uuWa+hgcA+78Jt/H+HrqrleeKZVoH
VVSBzXRpWiy59bkBvsuLLhdg/TJ7IYPm9QMMen8S+YU+GtM4mQSHtD+HJz5REo1BNUryyIjWiDoy
3tMDiX83gyKwXx3cY1MjUrA2kwIT1sdhiJblZ6ZRMKh1zmM3p9TQ+4HPFmwzg2eTXRaaeX5IMqzp
M4V/zeFmkKegkuIg0LT/4yxpGSTv/Yxr1Hd1WKd33oLrWOrnoEI0Gm9gT/fwyVouyZ7sVl7RsUWf
ciBFxcuTks607Gy3gpMYydCr9yliL3Ru++AHosUESGBxI55KieF8NeJ/U9R6S2T9kEU1RMeAMz1s
33WjVxpCKfhUKKq+Csx6nnkVNzbDzUNJHzwj8S+Isq69XiepCVAWiGKsCMZwN5pxF1CLCWIWGRHa
JyQhbBQJeakxrWOUqKQM6Vubccuxrc4h7vpr9W/gXSCYhhtNx2CtATujLk8/H+b0XapFROZtD7LY
qq/wsCf0A4tNQFroIQ6SrvGXvCKAqv0iO9HZBEsResJPkPtCz1DtgwMfi5wzDyTDCj9BVPfAaZmx
U7IoZyYWGNT/vSuLzvlHq0OAEs+nUCFHBGRCBWTYHs7YEe9gX+3dbGUk7nZg6+bru4Ad0/FDAzcV
MAD0ne1pAasVutx5Nln3IOvsly76B6uXGgtseMyptbyh7sAI6JOMjzXgZ/tOmvrRs4swN0b0kKdL
jxvIKQqdFpJpokm1uBaPvQ7e+pT87N6YRozeclsB4Ua0/EAzYxkC8t/r3KJf76YCt4z0eAxUk/6i
pCBxS40S6z8DuwZ56jBpHIKEjTgyocFFk2Y5cVls1hlng8Yia5t5ERGEgFaZ/NbXH5ndsC6MJDiZ
otSiMoV2ocBvwC8I2VKF82QTJ0Rfr0q8yU4RwvuFVOnLCs0vvWQZiaTrfvX2Cy5cPnbYfdFQd81b
BfC5AY5d2oURlPWBjxHxuKAc9Mm9iF5jnSlf7z23RoQdOXt8LbOkGjn+naCU0A4SJlZZ7CAeyP6B
EAg3xUimp+0u5VYgXqHPiKHrprWjstCFNp2jT7FoxpflrXndLCVq2kcAOrP4dLEwyD5mpDrQrCff
X3I29gteDcvRgH7M+qG4OEubh3nlQYGGrEBjpIgZ1JVE0/EhsjfPvMzoMbpO+UEc47Ke/irxN0bC
zdPz1VQbHFwpt0OxnZR8KG4nRwCg3i9yQSZBiaNaCsdzqWNAepBAwQyYokBHTTAolP4SdbFHXUhw
pxLCd7ZATsHF0TJgQNby3bi6pCgX+ibMP2bHjEllL4UmG/xWSXC6AVw1a2rH9G0cGvpNK0myEwCm
GoBU/Nl5Kn3CJQWyw1cC1a5CPxnRNo+zkjNbZZJEab/0mrGrI8fZCLIHd6evaoUrolPp8hQMJIPH
GOwONX2VNVAWoA/6ufSpUtEBqmE6l9Wb3Q12Weeq3jwU70jczbQHs6b8x4huPzy5QocDFcBtKW7i
ChhyL+PserUuaN60V0htu811T8OZhEI1l8o7FaGg0CggnNR7pnrU3gggjQdX9aH6X3GvzZ0JVeO0
VMQ3OAhLSWQBWmlzw5Wu7N4zrpWTH+dG5E97cGQsv49c/CvfOGYP7hs7P29WTforXuQq7S8H3GJY
7w73DfO831/8v1cr+/AbNjgFTwwzPu96G5WLrojKem8DL0Tc+GcEAqZKuufz/t/SOyeNBF4mKSLm
TSCP4ToQP6cHMQDWdLLkPiLMNhwPVgqlijl7p4ckVKJ30o6m+UfTc7X+AQcUwQx5BVIFKDxl0jTx
Fh4fML+37HpG1mX9+qc+mqtEdYNWNqq3zdxxh+87Yk+IxU4CVkACJvNEuDAHRYiqzNAmcVGelXfO
peD5sVk/w9CE4Q03ExfN5Ni5QYd4AnkJ/jdRABi5oA5wg+2mpuscV1e3sgdnGfxHZ/yNrbkHpHAc
GdcFqxUvbNR/PJPEkWcAEeatTdHmUYTbmBTltoIwLtV6ptSSBokPXyh3oCOan9WeiiKSHGPZjg3d
N0EQo0s5AkxssitiKx4vogB+vWzhVZLTmIykEa2ZMUhT6bU7BNdkHQMYzZU/DHkrwnC9dkXJrUYo
XyCWc0XDCFWKnmxu5+Uu5t9cjmFPURyJWtdzvF+xC8c5pLxFo1P5/Gg/vcVgXYp0ntY4R9tQGYrO
2zvRdHBkumYFU7OblyhBa4xRLXcNACaVW3gT9KuVD+EobS6Gp4dAlsKngyTral0aS7tG9jIaEBfi
IerOL/oG33PhaTP0QjS3chhTeGLln/0qoux/XMd8KhK6p87BVa7oFj1PsAlBQit1CsgdQGiapuyD
eUHfkLQv1sdTmIjrX/BiqvmBnF4gNdSz+6KwrteHRP4hKNvbMjonX92QEoGRxXqd3si9YkgOqIFv
j8ppRM1h3099ULpWJtShM2I3aMvIoXqIEy72SqbM9JSweIYLP0OO+b8IiUda0V+jQOkNPKi+KSJ3
EEcm5Zwhqv10wcfat80h64/9bzRoqF4tEyFrqP3Ps/kw0PIBBOLrvQgy3qqhy/q5gvpnybvnrxI5
kRajgWv342vqiQDcxaSAdShewnjF+I4H06SAFrNDORDtGn2XY0PRM2JPcZ5XSGTRcbggONUHNi1P
LjYHklMSuAAYgMUAX/qTtSlF9LNAV3HvPKQ5HCccVde8GAWULnssmv0XbQfUXZxZxBdRo/o/kK0R
vf0nRBkCB7Z1KMrzwp45Q/jy581zz7//CpxRFc7g1qokc01TEBcn/Kj69Ylli+hXgiXM86dfogVG
iuMv0GiGzIW8zqoIVk4ACZSBt5SGMUeNRzI+VN22esDcrzESSTQ0mYHwWSNIf8kOUYH0Lbn2UuQ2
jcs3SqZT/NGe1/l9MI1Oa0f1ECDofh/fmsFJoGzMTNfJ+lpx8qO4m6w9xDn4GbyEAuGDagzKtpps
6U7hR5wLRDzjdYpbW1hGitkV9OckZ2OAcs1xQjHt/0M7DqsnffTPRDtA8k1o9VJmvFQV8rTHJuvH
Gc2Mb4WIjo9vVFKfoUVXR10/R/WW7ZTQ/RJ602sGZfz5MiB+TjB4soyqNWc48QxX155eT/99xaxG
/4vvwOufD9MKpq7unCiexs0TFIJj3ZQmVXlESw5Gjse8RcMQME1XRmBFTRqgRRDHTpTN2x3gnpWA
C+6UbVdi0aTMkCyCJ1w8LYwkjRnLFLcgMRPDHkwIoopGHjgFZ0oojb8UZ+eCp8POjSRxRUXhGtHb
rRq2qU2/dEdoRKw96xsevROEQEFT4/IQM8vlXHMmBYkpG0U9taYSlGdaCqe+ixSmTy3ViBslU6Xm
NsFdHKDVRDjWSeOH+bFbdns+op0XxdpEuBkwRsUfHP6870e8weHrUHgDx9tm63iFtWLEoMNaLn1Y
/fMtBWGA/jKN2Yc3eIbkbo28CaWzHjYCSqK38SO11G//FZtAT2M4U77/+vfy7ZFlzlEt0PqGLk+3
/3BIzDsdfahwetgxWH8pRJ1ReJkll8JbFrHY/eBGer0T2YifV7MYCkhYIFpsktTPAMopipRoE1Rg
Skl+rsOMiRP2dX3KKVm5KfloEr4tX4wqg4d8PhCXlcNysiVbl4lBaeVgebXKpVMsAEGCqfIAaEdv
2GCaM6FkEPLD5i3dpW9pl7HxOFx1gNPjH4ZBfpMSDz8rpVwhsCu7ePUpOXwPcdVfttAgqkScfk1P
bOK/gGdz5y1VptwwWu7ndSkym4EuSdWu9vvAFrxQ1NaAxFLHBIXD95UilgY7CrlaJ67lpdjdnRUe
IDUhwaKrNV3HBdfWo/MvG7QbuNdkzplKJfWwdBs46TTEtozDp3Byat4ueywuCzniv9hHCFt6378W
BT+hApEpYNnjcbDUnnfc7HtUkdKMsGoRqcH0R5U0tTgjx5K26At1zkQyuCNSrIgjQPLuwplHAcLJ
0ynCdDiVCZWTW+Q76v86r7ti2VRm7ig2UNnJZ0sMhArKFgUdPZrdr3JMBB8Qf1rnRvMb89aOpj3L
I5Huso4cn/+ycgafAMp0lZF3pw2JXiSh+AyuRBe2oZ8h96d2e9Zc5p25UKCHbJRAFcVQpvHmRZLp
tq8uNyIrXLpWQqEK9f4D7PuKcalk6DZ8J+N82kUyPv1nP30HHxHGuNd7gB4f6a9ablqCV8mvs5pM
FhzmG3j+eHvGRHA43MxLdo8IUn3YQ/X2jvd75kT6gqWE0mPuPpU5VaJ6bx1ougzaI+e2aYYhUo41
wpg3sy+7MIm5S72kCG3Uleo15rsNLYjTzAg62gvbPbRQkVMKw51+6d6F10mKNrnBov1DZ0G/mKip
lUZIQ0r6yDPCPURixWAZNHWTNdfWC01qvP6K642/HasieFUOWLyA2ajPfr36sBTjf7815K8LuTkn
KuvVe+Lv+HfimGKR+BS3Db6/O/irb6DTJ5Go1RBcW2LHr78C7+07HIwyWda/Rk1dS+LVnMq7obAo
JD7NZYIqrnqnqsTZpdpAWwR9CyfohmQ9XfFj9oObh2xEl7I/W5Kl6z2L8eVzAMoU676QSkpMU2Xa
UtdMl0zprFo18lMDJ491S/gzoJRhrySuJVIXR4GIlH2d2G9ZbcGRXG8B9zg0R2gNQQEC6/XsLc2e
8W9pRXgn1zZnFr9GKbPIhFTlg5K3zxUgZMZKRY7+Ue8i027Q7e7rewjagemEwc9ieQJl2OgLoFS4
AWpkdPGy3rXa+9q0FaxdAnTNj7PRH+wr/K8GA1mmU0OUmdGUDENOx7v9VnOvvhdS+CHTIqVRl3pX
04tC2mEFfY214yJjtCUIi16JrZnAAUvNWz99a8djlkw6C0MGebofJfWzkjKzJUqlFYI+bNcK/ym5
McXlTNOLPWlYU/WuLeErK/nvovUpPbmbOfBcVxNDfmOCyY901YZRW5dUpAfsAFtH2DRoIMAqskP7
r2Q+UAJGqxWtdIBXiVoa+Yc9D8Bva9ku42FW+6sD7PWYCNhg6v7Bgo6jCAcJZCsXDMU9OxiRH8iT
ZQ0IanHzckxXRRNjoaSejJsRWsV96t/WbkezIPq7p+JUx239X4hvWAd1ScprkEVbvOLKjaDtGfad
wOJ8HwiQwRzHmDgg5IdEf+W+TAaJl/hMzuSs2Gc3dA7uBLRiIMDB4BVl+Z7lPJtoXwMij3g/GsO/
9R3PpQccPeAvNhegoNbrkIF81mzHoqSbe+7V+/QxcVnAMGrZikMNlkQQ+/NpKgc1GRS+nL8abgHD
SnvS2S8gHCuoHaM0+HcENjI6b7mA/VeobfZOKcV+Zz8zb8GcctB3FIB/6YS5/EyrVxt97eq9JA2V
RhoMyaMlH7C6OYH//KlljRdRBrdZbyCD+QSoMWbo793znKxovfufcMHnrdkygwl1HJBrFsvV8P50
r09+iCtOt93e0UilBxdfg1h5qFGWO33VHyIbT1Rk/9NG2m9hSgB7QmM+QfEbsU1Mo7hfG9AfOVbf
r/nPlU9+vGrFVJvBfj5LcOb+hNzWWMccFOhHll0q9Oq3WM5ps4J0v4DK7ZXJJ+xNfFHXdHn0hOQi
D8LARK8xarH3g4pIrBb5hY48SssbS/M+gsgF/QRX3ukE8F8ru3krH2SRA1g/d7KrZtlgkdu3Q0SM
DFHDI1yYOxI+Ihl2NXmv4uY+F4/ad1tEiPDq9FVJr6YaRXpRiXmZfWE7j14vOEwPI1So/jqsExQ3
6WgrriCMR5Z6/8keHATg5CIDM01FaV7P6YQjpNV4erJImmV5j3xcHJvcUuWmV7xns0jkRVvRD9Wi
QZ2rsKc1ZiH6Ibt4Cur88ZwzuEcW3dVRKWifVbei+CR3PGK4VJ1Ffe4Sfgn5cri+fF84Y565RNqG
vZuruTb4kVOG6EzL6VGgXSJZnzKis5QqC+d4Deyib+MGgRvJpTRhH3AKXVb/y4cV96YU4JYHaMhj
ya/5PtR5qsBFye1yyRPYTbzGc3kyOD8VQjdOfvY/4Xypqkpizk/+iWZzICp4zHgOypZdoe6yHJH4
bx+QvcRxUf4wm9boUFVYSb5HTjAg7Yb6w43szCWJXZqoMW75OHReTEm+d6N/pHji2dukGR7Snrc1
ZI1iBscVysIljTQiEq5A242ev+spW9Ur1higQSsMjXlbelB+gKE7X5AgtwVA4rT87Grk25cQ56mD
fJnZj54Oc/LCnl51SvQkuWkjIophKrK+WEmugl13jfFMOX/v9/OFibkZB32zMBigYYoww2Lot2gk
b2XMxbR36lzlR98cZWFdkcHVdwA7VPrlIZeW0Eo4yB+GnmY8NLZ6KXzLrAeMVXwcDqINJzKOeBqe
J7vgA7Cp8cxVQiGJ+Ao4LQqQ7zpcQdbHykmXGzhImLPgdI+AgE8kC+baKwC1DIZyRuAK/sVBw63S
SRZeO4no9VSW+hr/Nz7zGhMMmdaYIjNG2ELfBCcSORiFA2QCKqpbvlblveSTdKNBNFT7718IX/UK
rIdUCiGYCMXYvUfVK05R2aNn8Cg6bG3NUc1NZ9q5KB4ze7ny8MX6vW118qhsFNzC84mwF23x8AY9
kimEoiXGdFRN8/crB+ZUdNWCswy7WnRXdqDRMtBM0KLFpFaoiQ7Kvm3pDJwczaXgsvj0R5k1cKAi
rf581b4RckZZDDtdhsu7JVemDJVYVYcrW+MMxLxybNdZWL1yv26CdvAPnmM48/qUqZZBwS1Gr0CN
PWZD45p2nwPC6ARLXoc+ahpa22+1NnzeMP1Vt/UfrhqvIebtUs7Xg/hPcKGxYXuXJxTssf/J6svX
Bwmf4PL+JWO9k5CLswTgWK4DbZaGkaB6igWZbAzaIrWfu4SWGeVNgOjg/Ur6xt3K17KrRdz2QgfY
+qO2pOmPkf1cMQMvjoqpT3SahHWgCKubLE3cZRSNoalKgb+stQ3Ilm3JkcBACfGieJmBFu1MDdEv
llXI18c3+eP0vnaN6LGsf3pFTDq5yA80FeI90Kkw3W/Hafw/awGcnEibt8Kc9MD8FtfEYbgVu9wF
n4xbtjLrMHAoKRvcZl0IWq84zBFy1quQgPPQ72Fk+DHMgqh3Z4Ja54qmhCh7ZAU29EQ0/DZFg8GC
zbb0gVx6lkbzsGrU/lNZQ53s6Pdo2gru32WSRwLQbXSi7Y7daE1ovuv0GXGtJ9bS+WTfXnApaJB6
ln3mRiuoERPUMdVB0tD7onueLiz6b72OOl2C+acBbgDgH80OeZAOtFh0MiQVVa/QlDLbd429oJGN
vcmxrWm3SgJiQERQN1CF2AsP0nOq5I6ET3zL2pDAsSgfwdXIGI2u6yrj1WSIklwRgv/PIM547saC
ptksablCM7dIdgKnKp3/79AN86rp6+6thQTGdWPuS8PD9dO3q/+knbHjoUvjDvtLU2b4OAdg00/6
Wsx2XSYGkLURtR1RRS9aJnXvMHEl0NykgxvClI+x7QlSswA2MfT06HjObW7ZAEXFTe2MfV6gFyRp
jqGou2GPbmoKTQY/r24cjlMSeuOQbIOyseSbq7/2JEPdrAiKjUMeDDTyHx0opU5IMcW2n4ancOsm
EjvZmgSC9LqnJP3gFWOmoaHkqx7dt3kzk9vZiV/8dR+zL/t+DV/LuM40UMgYx1DYl2rVVZDvQGJA
RrnZwxASqA06LIHrW1FnLTg9E0hT+jMMejx9TAucaOApxKXxiFAtLcpyv+kWAIpbyzV2zIe2TA2l
sJ/Ai8vJwSouAx02P9q5t60zL1Bx8WJnx466wYv6UhwL0XHXQpd/J9thLaVgd7o5KnHF2sChfHqJ
Ziz7pmu4a771l2RXvTdrZfU0xNpZo5ERiJmK2mdsr86AawgP9g6VM1QyZZK6bCkcOOMdRVjWUNuQ
qtyM7wwU+WI83/EI/2CNuFBWQ7Q03WY0MAWgej3c/C9OGplun8eEf9bCT7OgkyzEf22Ji90Bommr
/jEzcVpFwLj6xB1UJHzZkjuY7Qi96rHlj1s4CSSa8Lkd+xE1o89BwmNR8vNVh0iF2k8i31gGVjlM
SDzB+58E30tVhIgaGazljhCpo2uF5lrL+CQ7wrF8AloVtfZkWWJo44slGgwoA5Kg5jV/ohHwfWXP
aKMKD2RgB06nGD4vcAzBVIdmq7eezj3WegbJ7Mnp+runwXcapGFj7k13p6XjuUWxsQhoBKjnVSny
T+t1+Dya3W/T2r36+lzoMTjxHVdXQDPB64Ck/UVgMjIA+Ks+iRJ6GTqFpYEWPzZ4OdYUXUtTp3pY
u+9QHnVV31lN64eJFt3VgjmopJ+Ij/cHGRVkcqI+T+7iQHQvkmoXZGUDcM0Nh8U4ptwHCGWA6fa/
GeihX0xseByTW+mTka1Hw6a1J3h9LR5duhrOXBY0sCeMi44NWziyGOSJxZvWXD2qpHhGz6PiOc4r
m/wr7Dy7Amalzy0Or85wU2ulF1IClt5Rv1r0XxmQRJcmYIZ1SwYQf2Uab26yolKy8efDwoGj2IZQ
BSMPBmIniZ7UWShRPh8XfLS1cQBy0+BboVgB6FITZnoP0ZkVAibqOH8HOVZj6W3l0hdcVPPlFasK
dQMF65aGmwp9GnjCzon2Mu0ftKykNPDRAcAbANub3HfOS/DFpfx1mfbfk18xE+MqpwS5gSNI/jmG
fjt4haPntW7MNCmoarZN5BnShBbSnBE3nJWLH4KNt5HPuwAM5X9AYEITsu2H3pX3fMPMuh8rD806
8l0NbAUWpkM8NZhfrcSVZLZe6eR6pfaUVHGXHA6jrRXvaSMSxh12WR/jyQYxjWuHz16rqPiMN9Iy
NSW5ogol1J9+jmcrn7b1cSB82RLgJ6k4+iUHV1UMPqM5HSS/TKbl24FeDwMBzLNnVu6V6B7q+UBQ
jfYYKF8H8kTURffXEaJqqD1SvYlktRUcxX+AcixrVy6q7rkHo5F8fDT3xJjl2f2lks/CggZFP+l9
kCpCpC2H8KK4w8BBTvgGVM24nE5ut1lDVNG/chRLtoW//kd4jz+/ARffXid3ayHXl/ETMAprPsKc
iytHpjbgkkauuNwDb4VnBAU7nLGPrZHUFV7x4YHZRZQ0h216b6gTzUJOe99+CtouVFQRijNEB6Vo
nEMKi9AcjnY9rOvFjvNkGO4W78TzG01CjpKa1yi7XMJGXm39vCmpOZzlw9Ub2j+5lK5pZRczc/Mb
k1MAqMRwIxyknTYrJ9dlUfuI1nQw6AYgRltTqfni3z3ZKMP32ZzYBE074cxt5cJpCm+uTippUk+3
nJDuHvU2zYokFaK4OHdkYnXnzfG+gAaFBXTiHZRm/pR5fk3TxiAPrnKm6C2LexzXfpr6x+g6+8xR
kRrSE2ykOJzpZEQbQEhuE9zk1CRTE9WYpsO67nGBXn9ATx1x6JqyRLWXmt8h/L03nlbjdAfdKCtj
yXQtzMvtWvgAkIZsQ7NFgfC3uRTxcLb92rD5X/2JiHpHlWBpcTonS6jG4QtnE5j8ByivnXKUS4kV
GPRy9WCV5Cd6kSlt1L8vulEvcleLtqKgVbwNCp4dS9SbZQIhqAPFNZx3amiR5oWoD3OJDcnctNLv
bBF4SbkfK9Sl5VWAkBTIyzJ2oT3jM4Nk8WQbhnTUANWZrEH70UKpLLhR8nReu9nirD229fiCtxUo
z9eQCgJ1A9Ium3tOEqlhEsHy73mkXWoIZwtOnTiEvxF9TzYejkgoRY4uSrfSvTEBgAwIjLlQ+vyE
a8bW1nLdAv8ImIQ8ym1cf8lcimDg/Yhs9I+nllRPhxXs+qUr441vVqqzTRhoXdUTlaUjrFR1CrD+
k8+Y/HNG+sffml48/Kk+7BqGpnDbhAN21IN4YmYtEMpWBgZ3clMV+ODQ0CIOegWKEb7k/b1zRHbA
Q+FHgQDC44itbd3JPalbYAGV0ioni2ny4eaM2Ffd8xmUxioj6DdiH7zpIpuF8WGWc3EoAHVoFUuM
ryl0X+dEpp9B2kMEOaRpyfDumOE3bKCED/sVptBqE2bC08LLLNW4oFCOHKWk7zYiUXthWubZ2ulO
Gk3QIk4g8sQgGVGwL3vBVf1L7BPm/2OS3ivG88raUPOXr0duYy1+hu/NUQT3rDNYb+CHxKpYhwWn
d3Bv9fwlJIg3eyb5py4FR58zJaAiq/sU3iC0CgTis83+YXDH/la8KgzIvLWuaNQL/fXJT7HyP3YX
xJTIMOXZBNR9GhQHp8bwNm7me0dqrUMBW9Ll3yIcMSGHS7DkA2OiN4L0E1CPC4m8c0zFpTDNrOWC
Hb3+Nbf4YqS3GuBIEv/8zPQaoYnaNOMc0ot1CIOeCcqgiscwz6IXTZyAWX/BPoiIch9y4dyATZhr
VsZqqO0Ubt8iUUnInXnhez9QiKPtsW3NaUrfGG83V/NXzyaAWsagP8hG7maJqbLA96ZGexwRzjBz
k1lTg3o2O3ULvvwW3fGJBYk6dh9T6E7M4j6RrmCULFz6XS24ouo4zHd3zlv5k1aC/lN+H1d4clNq
6wiKM8RGu4RvV6K4jOBFmtAtgjigW6zfSNntSS53vhVTMLQ3sYpI/1ejY+xI8rpzXwQRnsx0p/z/
c8R7UXt9QWByO5aHkyEItFHRoO6f3uCI+HtKUGCaj4Vlb9vdMqCqEF3a3IyvjypfEVs39CtEHPw6
V4hJzOvnCqzKD80cJI1syhtpQYiVU3pKMtUpGsr7pvUiEwMgszq9WcAIGZt+VqLj5T+nX23c1Z9Q
mOakCuH1eJNN3FXzBPwgdgVGqGRxKg/8pHRdw/jhocNZ7KBQNY/+2/ByhvnXYGBKqXBfyGr7E+S1
dZJlYnhJ47styDsL4DkJ4YiieWq0M97SDGe86BiPP0gBQMh8+UdqCaq0ck/GH8s0Z5sUd8+2O1Ji
7GtXio0NNIlS1/Cnrrn7lbX89HkgUqWYvYFFRSq6o11BnvOxEcI9alM95j/dkWtl9Qtc7YtDNxLK
ndTRcUGrzjMB0FgTKscU7NeMtBDjuodl//sGCjFGk49fTUkIqCpkEOouEG2kJ1w30PCJWabW8f8L
Nc61NSqBLcvtX/7d0saEhb4949q2QcCkWntJuHVomleh0GcucKQjJ1zdjEedFKIxMA8yQp1/+BMX
GmX0szi3m/zbTBOE7LQj/RfV1UwMm01vXacxItIaJhD3H79PAIbNp2getii82PiDM9hxi/LdO5z3
IamT+zm81gyuoavb6d0K5GmRNwbCD+TFPTK6z7SpsMSfXrjmG9mbSXGyOEEPhg5DUVVuiy7jh+bV
sExmXkRyrZyYbuTRQ3PHYUKVr/yI/OxfCZS7jHNPZ2iJ94PxBYbE8DP2JNszPZZC2Ldybk+Jfv5w
W4QFsxoLd3htvAbFsMud7WWMCu+btSVDKqM58OxeyAHqEQVmohI4FXP19x/cUhtdXl/cFVeD5575
KMCI81JIonV0DQ6BwHf9YN8X5+QdCuolWVC9ZCCMd0vj91E3otZLQiaZgUAfCoP6/XYfS88lPDeC
xL+aRJNS+S0Ml/rI3CY5Zrmn2x+oMqHbV1+ehCu88nd/TXIebIWjT0hybHDjn17qjXllF/9hDu+1
AAEnRmwNhB9CHu1n+qjSZMusprI18A1Zr6c00SX2NhILeYIuMYwNot0inTmi60iyaAqnT/kD5A6G
0J69t8TJhwB3H/9zwfnveuFWB9kotCLCw9hFAKcdR1JqHcHJpISSYYoliR53LhnYp2KyFjvwkZLY
isAAUhPAqm0P4Econ5OmHL3TB88VDNImNHaDDy/NSUU2hvt9TQY4LcY4ufQhSF9IT0oKzHGT/c1N
5KAA9hOkTOsQctwvSZhy9Qg4UBqpDYzFQxWOGmZ3jBmCJ2bIZuSx/FqyGgu75itGAZN3EfOzwu8P
aquYzukUR57MxwIl3pPi8fimOgi4unv3ac7ryxsApZ8iBpZ3KdQdjYhuE0PfkCzxr6Fj1P/EL2Ht
td9+BMh86HDiHkOWK2zMf3+n7lLM/3ddfDdneMbYFLBmQbqVguATq/Df7Hf2ejDnLYYjlN6JOrHG
pMIIesGqEVOohyiCd+ewopGBF3eVIEv3vdIpoJ3T2Dx+WSKcQBapiEtLJ/jaosm/fjb6ezWZz3CX
dGSB6h1ytKCfAj9n+I4oNK5/RKLXzYcehaVRvLo4KjPCvzXTrG2SAI7bXmrZEPkeM3xbjcWyo7+7
6093RlAjNWHXTgwNug4je/vF8X0pjd4YAuVz+vOMblvgzkesETDx4FTgw5ElMlmqQb96NFPbLWrc
WOpU/ZZTVNdtN0W/aEEEGLxpapyZ+aYHEFe/4Eo3ZuWa7b5wkxzHZP1J3qVQ/s1G5LanSRLfCuYU
s6m0wyMYuuFfZTsDFC1pq1jdxM5oe/1qKaH7KbGZFqqTlPT1aHZoG6XbfagZjMDAetX1pBGNny+o
SRHtYhxJ4L9vpka77t9+iI5NN2F+L7MuZkXZ24jFaOwiH3Pomkd3mWZc/Yh9RI2wBGNN9r+X2rHg
BnDubF+/Qxx7ekykR/1q5ygnDRXU0vxaJAkz/y/K3BWUwTUYm/3aBeIuguQGlOKbAV9YDn2lfE9Y
fDa1OYt7zqwPq7BgPU2aJrMwel0oSGWx8UgGUzMx0ccJ6Jen6pupYo4OoTdPrF+LIrPhNvOQ4Ypz
I5lLctZ5vFx0zZmzfCX84okZBBgNIGc4WBwrOCqYrG+vQ23Vmn5YrpEasDne6yGraJgKtiKLAdoC
SfBFvs6wJU1jJGYBwK4Lwlrnvb2BXCcdYlKvogyuND6P3aLoZzmpHEAWtHD/juA51GtoMpc0BUN+
y2juF6sQIjGu5cvEw6VrwOe4hUwCRzuMjhGMZgARw4DZo1oooKHud/WJGkxVA9RPtdeeUKfexEor
ltwc1SK8AlmrZoDbbY6/hTw9wgwl9vJMxnfT/32nTSDkMMlgQXKlQQx9w/JgGStKXXt8BaBKJU7A
xY65QAU8L+qbfA1PkWZmg824mWgrz0vI2vnaRnxmqA7f+H/XcsmhxASAIBPziebReUq0deyxZNp6
OHPaV4YTDFmx6fQyprPG+GypJlkJChZk+H6FuWtGxyx7Cvugq2eLW5DHko4Gq0XUPrsO0fsVrAFw
dHbUc9kWE4qqgRtpFkXO4a+zS1PutCBEumVkrSvJFguLq7f3HRyaiDgzHm0VaTmk5plfWXDqIgbZ
c8Kk4sIH0r+LwCDjGOfPmEHQi+/KxtNNoiNLdm6pWpPCWkgHbDClXCRUP+o2Zx8aQ5ly/RoYGVCw
bthjGw2Fumt3UQvgcuunYYpicIt68aBhAST8Dj4TPJaRYAmS4UoiWLSf9cZ0kGdTl0OKSjStbBwh
AfYl3fYJpIRe0ROMhFR54zVx/9u8zraMU1aw0iPq6aZrbNNQPC2DITZBNRR1L6pNbmp5/EErgCmS
iCHxmre5/ShdcT0xzatmC33usAMxgat0wiIBxFnCNTg74bzG+/3NATUn71k3v3wFYs0xVBBulYQ9
CWP3ZmJqn1TwlJnJnkSGkzBEYCwNq3mJmIXL+DGWgXfKmeFyCnbKVf3fsAjekVCn4ZMms6398cgh
tj8C9NQd0gEybWkDyCoMWvixZt9IfT5wx+YhjnPKztn0MLYKj4B1ghZpKUeOvSJAF2Li7TQtXuC4
/9c88+7fzuxkOR8wXmQB6kHbUvDWntSuFYSjE83viZeNrbi0alOKlD0fm/pfss16hN+99ZRKdlWe
hrYh97/0qyHdEi6hoNmuclNeZSA8TzNB0rQI6baHahVZY07tWjDEFQFbq0yRpAk7eZJiMl71cDFR
+5qe9aRF1aAbz0Vg0s3t3CiWcQ6C5hB3HxWMFf0b/GWQ5WifWjhp8Kja79UVglNyZ/EPUh4nQXL1
1Mdv4nUSKhiWjkdzWBPNfDUwe1Y2Ib93ub9vc9B/B6o6IqmgCP8t2g3URXMLxN8ysTFRSBZBBS8a
hPW5kC2Le0rA+obEH98O27FuRH1V3XJmxvO5FSiZk5Q0qIOKvyvJKsWGtGqo8Q+z4/+DaurKwmq6
+fh6GG0Q1POfai4bze57fAy79+/PW1Q+QfrkrK61yCr/c1Bv6uxllkHEzqg/D/TVPBrYgTkOXo2o
/rviWRdCYy1Uqx1KdUDfXGjGH7FCUFDFKxtQfXEyJX7Q5F5USi689G7yi9Ovq7If37144Db54kei
ahBtehll986+eVG/lwvFxjhJlnhxKx5D5OLiMKAEHI3LqQfzpPDf+zQw45m+p0Zw8YxObIgwNev0
MAA0VbJ8/7OpxlOFNlnf7ld268AL7Bb6lvYcRZBygO8bcQM3RW7DyGoxPE0JaEyT3muLdzv6/BNV
m8eQDM9/e+O/cBUiMoucOVLARsSRLxmOAXOBHzxA78rCeKMWZaq9jtvp0foCMligNvCT66fC4AEK
tnsY6CS/ja0TudKvkll3OTWkjwK0hTxXy+2zM9XF2HuiU0mlguMdUs89ixtWPn5Lz/L8klvxWHHT
nVvFt1KwpaYEk3vgb2WvWW/mXwcuKgp7xNNbr8hFrpXcKS8n/KWRcVzGcWx0MJkHsNSnj6oCRI+j
2V26F/SjXiJhnkF/zeHLu8FfcjS+cd0WkZ6s5pvyCoHpq/gX1D4iDg9AOLhZE1KRda2xmn5rgjEs
kVvSK0YCbVp41LZ5HCkM/1XeHaUMIw/prXwZ4y2CniQTj5NIMVvd85yHp4OmKkxImzCHSVsiciON
cCZXUCpJ8qmvj7DpZ/da8vvDlxK89OfUHDjOaJEsgmGYaqRhPcxmIWEDQS/Es+XJzhxaubL4enfi
pLdNzEXmq2rK8YY8u7Tp7clOaUTfLMTZ/o/a6AQmYSSnuvFrKV9d4mPXav/mBBlkCVTc6IKaMBe+
8ZZcAdio/xxeVfE4zvocwo6zv6IaY89pzj5vHh5H0cI76K2pkJ3fCki2YxZC3+aOLkUhCclz2Ki5
9ENlKwJ82ujFedjVQyqKKnRuxr6Hku/yQmlEcjvZocQVqDwOYHsJ3j5MaTyvNzkb+yDc1wkRX+6I
p/H1M5B8eHdJ0DFc0Fqyq1ZeR4NCk4SmjDU4MSGflHPc/m6GiYA/smtE/4txrFAeFH+Y3Wx1kvRK
NOK2OMLkaCShFBR6dsyqT/7iuwoS60ugD9NcEzITvnpgZXY5hekOYgfkVke5PKwGz0NWSK1J0isb
vHFcyamtB7t7w3Q/YrhFBQlT3T29ZgTiuIQQKdkZh9J9wIbpDwi8HsGNBAxlnqXay8wSwQ0y/XHq
0HhirQAfleJS2r0HDWb+pmj+sG0VmJcopAaaDPWPezL0vNOsrjF0apmK8LjxqqhmS2FyamDVYl0A
5vLRHFfy0RlLw57uGRldvc/j7kfrg+QEKtIppHRF2UvqGlRZu9UcmuhkWgv0iOeddmAnr7W6yrAr
aXNrLjoPXh5zTtBbfw4p4VpQtEKdpehcBT5a21EhWr/oMrF2n+ds2RGbXiAly2NhFnpsBe8LrTts
jUjEWANJaTtr7V/wb6ZWz3iHmJ0vzeeu2IJ7jsby4i+hursq8+VtsJ0za+7dauI6cSO474zRZryl
dbR9/TjFLtQJu80O7ln/+DenAzcI8vftdaWXCXefl96e94jUJMyzSh3PKsH2of/J/ZWdKRudI7rJ
7/gYpDVUW01XUsF/mpc6cOR93vf05NK/tlohhyMPootyKDzE40VPhcoaxUUgDWro3o1WrQhbOJus
DgcCxolhNIy2E5IwJDJsiftzyTipb1PCNex/baUhycgoIkSNXP35OhwEFy/Rmo3fQHdE7F49Dvnc
Do/JVDMxN6/ZHp4fEnYwbjF6tDmhlwxcUlbxI3+yWGd1Yh8mK4VGiBbyI1TaY4TEn6JkXK03Pwbf
OQyA7Iw7/YP14gdJrnD2H0fpX7T2scqt2Sf2vfvHjcv/mYfHlw7gUei03Ok5682iDUw6OhfNpZSj
FEBzJ7TPKQDEXqRNxVYN5kEclG9YVlRBGHm8TgwEBJ2KjxEAZNSkChbnXpHhx5wQuha//hVvDA2H
79EiFoG8npYl/0OnhZKby8N4mDomeSIupE2OhYqQD842q0t1Q+rLoi/w+xGUWrlFktSpkwFAZJ4a
cB/xekog2UJS+0xGKX/UPF0RV90kl484pElHBelWuZtsp4FJPngCEWlmS5iDcvHdy2p5x2+lum1G
Bv1yKH3b2AK0g15lIeZjiXS4lmv279CJASWVStSKg2pAUkt7eZqgYcr+8uipvcBGguUUIP3MkwRS
8kb4J8wENT5Jo/CkoOLQIcTH290SsE5gE/4FjHSilWqHLXeY5pIOaQQOzyCBj9Z8v0B9zN6giTvZ
MnAngd4gOGDKBiKN24TIE0DnUZcw+iTGXpVBAVe0+PSVtDU2t6/voZ6NIuiqyJ6u98wGWjovbGWw
+6FXmPThI4I1CJ7gGjA6412qLjvUweinKVScTUzY6WUtTFvTT1GhKHxI+b+Wxmfd6erbAuuL52cu
b7o/Cn26m4Ro1e82GVv8k6B0wBgnxGDNfpY5yUyc9GcAR8wvq9h2/eaMZwhBlpKXDUPDVDyOaI1u
NXk9ZO6g6M8wGQIOwwRZwpcp+/igUuCJR7I+j++eDRPGL+587oS0rII6W3V3VimDzGRVSm6dVlLx
7tbO6dq91XS2LbzSFomWk1+g/816BQ9UjXvyZwlzRcWA2Sh4Dq23IofGz5xJGMHcwYxna4uGrQ3B
oj6qfvPvDM8fTimDJyzzuFFr2loiz8AaeYP573GnwEqEHIoxYaGXbLIhnL47gw+GEpRFSSf8iBBm
PfIOnVbyFRymTKLNdTl7SNbBCC9aRgk7vptWxpoUjt1aAVtGxkFbi8ES2fhoLQA66zC9IDA9yhxB
dTAV4jN8UXP8/9tivXqFkWeGXfUjPFeq2+njPcfcOGV5BEc+etMR/EYHE3Y353I9uozf8ctCflme
PRxgap7RlaR4Ka+u+J4PTg6XyUOmAa0oPfAOrdnYd9n1iutvHbb6FPaE8kqx1op3cWwk0HD147Gq
ve7cDBU2oaFjlhjrJkXoNDMP6wlKHvk4fPUDBRJtSI+HqamnurNtBjxbRXq+lbJSU/49aWShxPh9
OPQizH8n9vZRoyog0U9NpW3fJ6NvjrhtBuhGMnIDJ/uWY6sJvNZuLdr7tUQOc0yqKhn1+FUfTSbN
NV4RAkPWDUEYdZU/ulOI1B50B00PuToNR9jAkSUcn+rt11ktshcEafW0+dSTSmIW915eAh4PltVV
8VNyzBEW0hPJtNWVriPbFWwJ9eCykXfKBOhtubm9cBGWkMnCitOLTdTKnCTsquVhGqjO0L7T/not
esFKNHb8eFBeFbjiV5ryJwqJlEUYeNQ4w0MBN3sF6EfGCCZ1Fcu92Blhy2Nr7XpU7qqnMhmz5mCP
JOkVBqZAol9bXa317I5woZyZdf2M3krLdnzQ+CMLmDPT0q/awCNUjOs9QYkM/rxXLiTTuDpTmw7z
0DGlMyDpiYkCeAQmnFUCdkmH4nsDNhqhiK8DsKqK+LOcbloKzb2m/BIZP9z+OPIh9sKfdhg+H6U6
UyKs/0nxhs2oWD/PRBShxVaY7v+95v/Opgk9MsqB0S5XIgEjTj0MX9Wj7xS/EsnkeyZvY8+6JjEA
+ktRNQaUyPFapIv1C65kOYe/n3t71zJda4d1JqrQ2xLrtBDt2dPARcdVbMlz97f9AemQiliqN9M7
AwSGZbCQTgvaOHM6WQSDTpf9MsBzdfWJwILuwVL0ONSlTjBWc9pAD2jtvADV3L/ZsQwA3XnCFLp7
rUThYuemwf8RINxd+VLVUUNIzE540Vd6X6HfBymBaGV0LzIIFO8byTqv/XrAjxzxoiW2Xy/5/BrX
vkydF5l56c1g5pnd9ZGWRL21ocqSgt67aCphlMI/84ZLRwxpZkx48RNhG0ZgfoG18fa2XqO7QhyW
wcXphUyXjBGbSGjyKM06XRwC+iLeDz/sH6OLMCi6FiE21jkklpvMt2Mcu403FBpX2kan2apUYqAU
j4b/8D3CPQtw/EbEQG8PxGubFIT39sHoyx2L9t92TAMOWfSfH/6WAr1vCYeJpDtyV+v218H+xCjm
xxnWbKeJjxfVV9KUAVn1jhXD3BHkCQG8gdnfB9FWQaFR3OTB4s0AOhq41F925aK4d7pJPycDFNnF
GyoSo3XiM7HpDlqzLLV9CBDZaYq16YlCW8d7nMP+qG010WKe5ZHvQpjf9ovqgyvtQt1DqRCLvKx1
34BEAV0NgRfG6fddJxz5KkWqQtue/r7vF9TU1Mt0EX6YxK/u0KsaLxmecwBFK3IB3HczHZ5oPa2o
TrpUkv4184KrH6yEn1ys8ICRyNAbQE8yNyjPqqSE0mgMNMlQPICG3K/GeGsdKUfCGbdGGeamqIgs
6LJ00n+XRAlDCv0eohWSy8qnohEDvbOgdmmm6dUtFaUln7o1AvO3Bvqmb1n4O8JQ4rY20X3A5Iti
zDqB2B8nDk/Dx7SgpnZ5jjj2/QxvKqksFrWdECKRy/SOvwDb980+PPIOibU8HIzODtm/eEv/LiRL
rT6YguKjUqbJSUY6hsA1BKVdaGInY9ZUlfjV3l3Z3fKP10ToShTXFHgQnh8eIT1Z6p1NzUQjn6cA
ulC4jG8TV8gNL79wT5W5TNmVjfPQ+NK1F9fyRRNjaU+tI9p1AheB1vfYPbqrNlSrKp3Z8RRq9FNc
LfTgYirHw5Lu4VDoGFc6O6G/6PdHdCJUOQkkh1KbLTdDAXV5GOYP3cU9Wfvgn+iWErKBxK1790bO
8O1xfU1CgHait9t9/OGzxYSthi1g1n91cKJxYDs3tJaYyv2HORh30OIZCGcjQdz5I1R+/z53wlwr
7vYZcBteHp9JI0/yp6/f9GhVxbB1gySe/juy76uaU629yr5Q7jNs3itmqTAZQXKig3sv0SwTfuK4
Ux96Vniw5ByAaU549ZfPF74MREYFQbQkNGmZ50fQygcXQh2kJAuxB2rQhdka91ajEZg65m95zUTw
gcsVLOn5foAhow4nHb+iQPwoN9BDgNWbtn21ccv0LVX/swZ63EXCDQAvMMGtAlae87QbXfasCW6h
3mn+bRpoPtC9GShy/VpVRB588D46xI96iuUnzADtvprlnFzPNHfXApZiiFKjcrl+Q6vyBv4TwdZb
lHig8j+/NqM4cYy9tOr9xU9fI2Gxm8GdalA16QAUlOVglZ8/HC+H7hbxXlZ0pUakfwsztLBHsQey
BAsslF3Qxy7y9qdiKp3+dwNnN6CIRbuxKxMSuOG03oKtCXmAZLGLpVGWLQ/5ZxPAn1F4jzdsdxxb
v7pCw74P+qOHX3oQFAx22WzSZuRbaORgVTN3+3LddA4YyJN5RL10iFz9AFwLKq2Y5xCN+TRiYh5/
sNTUgX3YhBoBwyK7+RjA8yORphS6fQGD+b4pZrB2NiJheosqUmOqplY/JEMMbpHkEPGZs+YXr4mJ
660+otlxPnCoIA7Gyj2RmmzsQ5b/Mo8uqJN2MldhaMnGofxO5wvuxZIAZcIbHPScvFkdUqanuF/8
AevuOBuxTUOXkcN/pU9y44FTzGaNm14sLJoY71YFQ3b3rCw+O48+cBgfth5+yEXd/ytQRWpNiZ/O
H+84eSh9IcGMRtoGNkQZzA0Dnei6DVX0n725MImoXxxOu/uGyulhX4OgeCi1YxilbS+1zB5f4i9H
KFhawLOmTjSsKNtgsPjwJW+VGu/LEI/TCxhcqprShHg8nqwO8Zhy1z6ljmvrFEr+G6/7C6WJC11s
hmMY6HweRk9IApkKtBxbdnLFMm+x+K9OudfMEDV0SI1yettXAZRE3azUpif7LTOFIeZxA0SPJI7Y
5Gsv8pqfbpOV0GOPyDwqfBEoY7CZtUfj/27DOSkM+rw8aLjvD7K0zbLZALztFwD+bROBDxMvAYuG
fQmsZtoTLELW9xcADexXd8OflyGh8aapLeehT8NYayPzGgRG2YpjsfL4XJ+2Iihpp006cLwnnFff
N4Q4khXAX2Sg3xhDAvK0y01Klw5YZ2trZDVT0Qx5+Muj/QFhRABtav0RNBRKEK2VyqR76A3VGfMS
VmuF3vo2PVSu1LNJsYMtKkHwZcMaMGsJaU1KD8wbBMdhl4WsFo2T2MAeVpovplkwXe/JqqMLulq+
vmkv0P8KZLY8pfGfeQp6fjBJ5jbgWBK9dDe3oHTCk01NBVRLrVf08eNj7YtRsRJ92I8zOckyq75a
482IDnZrEgRTNbE7EENwWN1eT8nPns5avlln9aNVqvIcZn4dlqGhQyIXDCScXjSqXxJ9skEkJCcG
hVf1dY/S/kRUQQyDRtImLbVNmiCKSWCgEUPzCvBVisuf1/oX6aXPsiGkDelNsTaUkrgLjlW4MRea
DFRx1+syfm6sq0RrTbUK2EjZ8flTjafzXY8nIHLxPBuqJVIeiInQE3TSJi+1RtklF1y+Po63E7Rl
qVwKDiSWW7aY0h4KoDduKiwyFW+kj5av2QtkjWVhhqe77RpUzB2a4sjss0Hi4gBoJ/+5++7aRSy0
1DKBHXcC+HeYF8Bzpp+JCBUWxy2v53R7OwG9ulug7iUpg6le8RnCP/hFiu+/zEF9FwfJQtiTAkbR
0m9hbnDJA2ny2ivPy5BhoNbpHwwqcFonWoNSrwcTZF8j92TqvRbXxfO0yFMhy0qcJpTwDKxBuqAk
28doyJ5GpHq0jAW3I5uuoEmLEtwyBBYf/ppAoEmi0E+Bp2mV1B22QxCPKpmMVrjfY5m0UfJiffF3
oAVLZlHfV9BenIX1Lxh2GwSoUCzq0Eaw26vIEHpIUqIwFAJU4a9zFGRhDWWpjXeP0GKUQTv085gD
5DOSxZdAnn6QaDsoYjwnN0aCPlMrqHh8BtFH15mH5a1EvPIP+ewyOuEwNJW3ZmuHsru+o3eR9RYd
Nwkj9LR7K47najDENzdI2WS5lp7wvM7HOg0QAxqMsB1SsUk4l6o0/8zFJb58x1HpyqAaWaClrnlD
IyPySjgn8hb/lF86Fy6pP76b8drMnbV7gnRiwwPIUF04Ox2H0+KX+/IpL+VXobsrxBfKLncnYaun
jBcaZOW1xG+H7+fJbtNvmcGvxNlhkCQ8gQBGQvYL366idCL3lMtOceMx5dlD/xt+GljhgWh3xn8b
RNvlR/iaUgIz1gmsiPdIVvKp4HPsKA4MCg9xuEVY8Z1ZKEqjLPm1TTVhua/tckcbOHtNaeV1XerR
nEV7FxklPanX6CNbj90WpQ3D4RdIuQgeiTl3kfXQXP5+9AtzL0fT1//SJnKv++FoPzHr2eJR5K2q
Muhgwd+GkvAAutMd2AaUON+kXJIEpELef7wiLARCbHuFloUk+HN8WYEE8VqKuLqWwixCr8d7Dwld
6J55FgVeMs7qPzNKeZyuGGQueUCSPU37lT90P0w27g+05r6Hg2AQEnPK6zTslGDfkAaKtHBl2+vb
gZPOr9iOZS08xrppZr9gV6HDtHHpYzoOmLo7pFj64wEdXZD9oRSWIs0gFRers9vvujXn/21PrM3U
gg+0cXtEn8sT2+T707rphyELudcOXhW+ZY22A4kLZlF0dId5+fMdxYufhMfSMreQxrUkIccfC0sV
EMC6Vi4Bez15oKpGUxAQOQqkC5yWRPfhx4AWtNDs7TT3LKzPplBQdFP3SjDNdIqPa522dFqYDwZe
ffbr22nWAdm9zQQjlq3h6jqJZYjb7lRo22qVaB0d4bFPr4ujXjjsXoJ5Zp81kSfQJLiERfhsvOJH
IE5XP7zpEU3czL/POYuMR/7lMG4sSP+S2ZaLfjE9deYxM743TMveUJZbjPoDtQaT4t2FmY+9STgf
SeLoKFBB+ouzzmnBxv+fc0SpBZ34Y3OiHdDQds/afvTRL4aXSUTpmqEwTpNkI4O8ONy/nDfpc6b3
Q/BUh8ifW/RsbUat0TBjS1sqX4KVp3SMsKhw9CEAbd5qFr46ar+F/KmnrzOwnpPEPJE7+EUBZP//
306LTUkDsLiRM9+bP4R7QZk7vUGOxE3Asng8y6CaUkjNI/LnrrOAqir+4SAuwCEvN5+rKSdQj9XA
bl0iIsK0uTZnZDwPWovzrt+mLudYZh9twE8zVD9X0jWhd7qjetQjsChHuysKFSgvIdncwrIGNGgw
lHomwr2nHBIqJfxbgHmwA4f+Q62TM3mgcRTm7S3nvDtjO80lBTUCaFaq9U/CSN3uczCweZnHm0h/
9PKuRzdi6FvK/+gBJRR1mB2MsrYbGRWGVzovzx94APLVRH/N73fxy7DTD2beeNB2cJ9iLEcT8Efv
tUVIQd2ydYQoVY5xnTrTb80rda7E2rHoGS8iBPGl992SWf3+v4unPniLbDA5hwzCx/f5LI7qJRWg
s79JuDzm68w+//xOJiajWJu2h/H4AgGnowoxOVuWKBgD9GLm+wzKDC7VLcoro3w2PozF5X1R8D70
Ts9yKURpOjPxszHa+W8dUWds1FHHHdk89ji/i3YJPuhxUUZSvELGbVwGcAp/0btAHI6eGL3jlFq5
abacbu1LHIXqdVCLKEkGDkDA+TBn8MW/VAg0pWYNhF6k92GCT39y2jYg6oH6D/ifHSU2H35dyx/M
tV5Mt0L+LofUNX78RALQz/8+IqqkTl1lBhbpoZfbivlwiiuGF5gDT/54jK/WZXOAhwvt7ep3DUIp
sFPiI3bg+vR4RQEeek6YVVTCyjWSiW6vZjuwMyXwfBGBavA29uIc9EeyZ5Dd3kGza/lKOwgC8oKO
3QD8j+l+Okw6Ejj6lnj9x5fW0etM/B1D0kiey7yuHp9+4PHER7qN1xB/FGJQXy+y9NNtq+b5eHPQ
CGUNM2dxxYIz4bw0zop6d0xLWF896L5Ip8+I0MNhRsASRAP3bZaKqMhKpdQhMUJxCA28DS4Dfm22
FRy3t1Hy1X76rRtEYMqIuyGGJRwH64LTZKLLKhEG8RN/u1JkjEnOFG0C79A2L5N9su1c4WDxIkey
tVi5Qg8C5+pA+tJEtEw9DWU1DXf8SSdA5MuIWfAYYlTk/1cnS2DCIpLckCHR2m3bSZ87XihSc5nM
kLfWrpHN5AZQMjhyThEMwRGu+F0pz5V6y99C+SKaT4/31T82erdnAgGxUJMwmvS7onDdIyT0itK9
UESQorOBoB472aQFD+wIyscC0DnT3Lz5/B4P3Cc8gYTaP6G/N2OBDUsRC63INYRuS6uDLNwgVp8c
xnukdOzGdwu0JM7UsjVoSaOhSJAmvXTuw1sJh5Lvb0DkVs+nD3hYLk696mg+cSdj0TvnlzI76fpq
b3mr3RRg/6MI4q/0MrYdI668e/MmWpz41ld38awkoL6dLxR+halH7IF7u8Hzn3CSH4o6f52Fm/YP
K0g5s3C7kUVPk7XTgja1nh/YytTEmJvz+XglBuc9XxZvGXDVJRfOfGEN9wP+3AG102TeRg5l9+zW
zegiZp2BggJKm2gvq92ZpkBgD349WaESTb5EtKIic+SgXzPhlxn4BZjs+z8EmB9RUCx7QXNeo5cb
+09jcSvT5vUx9oSkEMXRMxLnJ3ZroR1tMFW1ohznx++WA8nNS3yrgYUdgtLnIvvguN3ygyfxKrH3
VLT6B5UkBnkm2gywVmUQUv4MVAIiRMVFSGZo89VX295puvdfwcXocfB3HYjrwe5vp4nhZqHBY0BH
XAacZGK3VhTJIadTmRFp7+Xb4jr5OeMzPeeQIWyONehlz08trUWGM22gPqas2oTBMHuKnJUI7aWl
LjTtDSSnL2TDl74vVkB3F66ydXqMpvKl3lu/bvpLKoSj7F4jOzhk5FGQcuoXYp8mVQunRF86hd8m
u2ZA19pvKyLNYaSn4CcrBsmP3Bwbb3zN1b6rOq/4S9nXpfBLKzUqqDdRnsWG4vR8WW9UC+loUBXV
Kl/3s2VyqcrWsNoP8yESOxZ9yT4WF3E440eFgQwpiOZlcQtxrFMn9HehB4LEQ+Ziqaiw3eDQZdrO
2bhGKtLXbDhe1WI+gpaed0aUsHeWZmLLlCVEh2AqXGL6+EaF2t6y3woNACtqLfF1hj21ya+g4bxS
uA8UC8LNyumtiJoaziscZgYvKVyecLDb3Do/b85Hqe6/PlytgbEHySTsSThNwy7n/wxBw9lUPydt
hATUofULcBRXEBED6QLsq4L1lYBHLvDa6i65oeoCM8vRFcIdX9hjnX5vF79b9Ms024DTyXkeJJYd
rj9gXDEhNNqeK4xigwgLf7C0y3rXFvUyHhz9bj08ffFiGqULLG34N3Vi1nfM+Bu0/NLLHOeI+XCf
hBl8w/9vqlumR9vI6iejHUFrISY0hMpv0Qsdcea4w0+EQ7dHWIjaiqjeP4/0KB44lfgMmKz/f/9R
YMEupFPVVJR5z3EEuFHbh0qzS5ccAftU4ZySFVv8FY/TuyBWlSK37hALNrpYYnsJjoXAjrWlF3RB
NPABii9CO4UwHZX85i1C/l0I9w4/9dZ7kWYAETY6oIKPet7ZUMj2eDXN9apT3/rLlpMl8rwCdx1w
+H7dqwd7G6O8WXL9yTREurZpDy/N2gws50keCgpCWPDuzNSMOIKjMmLWLMxKbdYxD0nfJaAN79s5
TZdLoLfKWu0J9CqOEqu6PuF/hYZfW4o/aDGQ+u7v468qhUMeJgR2ATIfmW874jeJvr/CkTTuSs8A
nC7BuFA+vaDbxLh0gvCam/i3VvLj/Qny3mlI8ly0HvD44Q0vMAd/3N6BQ3vaRugqbHshKYAW+ynk
7sfvfYG340MiTtXNJ0xfrjbBv8kcA4f8FM7pq5t+bK2VmSH4MbfttDLJUbzTOP8NQ2imvJp72rcO
dLFnHPhJN5YPfF/q3Dw8CWmuBcpTu6drO7ZpfxT0GDfEqOFVaY6AkGnnT8PBfVe2E8RKiWTQFbtN
zTKJWFIwzo5VtedFhMubHXKBzNC5yjbs9tlxyksEgKwRsABdtx6Zp80eSVD+TsXZ++au1FG0noqa
I6d7Bc8znksfTj5PIK/yCOz3hjPaRori7oz/GP5q2cAc2bhbaBuPUgImwa/W2o+h2aD2VCQvRin8
d+jT3sBwgrSElGsl5WwWYv4692lvyYICOVNkE7H4nPaBiaO5OLTsraY0FBaaRC7EOalRAD6eDmZ3
M/S9Vhe+7Izgv8dsmQvs8hdUhxOwhyD2aLBLNGCu0DhTLkP83QReZdcVE9WRClDwoceMDAFbVtbs
NvpmL64N2noykHnCqJLaHXcbuOB1FzKRnOgxnhk4a+LnZsCw/BqWrkFUDICYMfqPteJwo8CyTTg+
OE96U3Jivt+NkjeQNycqh6KCFQzFOGgkPi5p9ciNV5BOk5hyJFNl4K2tjJISSror5I0issohYAgv
q0cCu2VQV/Z52G6oA/XgzaFlRPRU2Lb7VyeehuI48IGfljHpuV1rRJUej/o+g4OXbOkhVCuhEAdJ
PJ6rPBdUBvvg4gqzv7WkO37lnxugDry2a0N69xOdG6LyNxh5sArWQ0wjC4QEmo50xZqMkKkPHtF/
Za2WAVzxpnYscdb/E96rt1wzJeNqmilH3b0HZ2Esq+Kxyen1JoMP8MxNJxQCkMoC0p7JSd/7PzYG
Dd7kNNSBTdg+guMDf+W0lIyxf8UuizJjQlVQwl00xTEaskW10FrTrhqyuL2zkunJtvLc3FRFOg/v
WMImSpk68ocSBrZe0DDWsz5259HithSOP6ppxR3YQUx2m7AJ+xrkuDo9ynnioNR5w4nTe6Pljb/a
c+g7aJpKyWqTaZt1t/1iAiFn4z/aftW1wO0i8AVcgl05zvS2WFeLg8vjMvxlcukm3rnfsQDijL6f
pKnHihitX7XsGoGB/pAla/vB3h+G8Hh9HVSs0Rv0waROcZjkfRbdbyvRgMj5w/Ekm7fBOpRNISfp
IwUH5STYC5hUDoWjWBqIQ6QiZsXyQHxHNv330smWScVRI4XnawZWrOhJ8IbbLkrdlL7WRon5neWV
r/2KNjPRCs9P7mRmT6hsy54/ZKjocawoDYxJPAMtCEVXt1IZ9LWe6eldy9fsFnJZPuTA1RzL4yTu
S3pcqHZsnG0xFnqL4rrHtZY3OnTiewhTeD6JTfrQNObF6ywBc57SvaWCxh8Immlq1KSSdlWSqIEE
C7zsQXua/bjKF/9k7BqL5wsEVvC1jOG0afAtBca1JBQ8+7Y3iHkoFjaWDXdPCI6yDilWbF0nUvEX
eiu//8D25CC7Fh6LiweY2d4cJgOEjGavlyqrVRXMVjR7DbUcmB7urzrvsR62IWvm77I/OS5Tw+Tq
MSweaDNzfiNClJlXFMLaawqA/tJ1L5x0rT78cp8987ZIj3Hq8GnsPvCfFiO/OZoYsslSLAb6xRrt
4eJ6GUqGO8PmS1NPrHQKqGkZFjpTv81JatOFDBHtCaevboQz/n6iJT86NWl8+ag4PwSWxG2g9Cvi
QfGbgvc3CoP3/7rX3J59oQbcYCDxqSAlaDeDyvwB7SuIK5Gm/LlThwCxm5FyJUwBLevZZxpot6E7
HwJA44RdXFSyzDO4I8WPcPZiJWHk8urlH00/oPFDUW5sxoKLwUwlceKhXs3LTUrmQRo/B1SLhZ5z
wtubXQIkCGPA3PWkjnQPpgZdx8u/v4/504PTV/dk83MhfXDHvZCuIevB4KUZVD3ZC1sSk6IlgQcQ
xCZWlt+zoT5qCsFhsO/uFMEpKVlk/5v56xhzu3eDwGYr//ZvLYJkVehjnNI6VXs2c3Ua8Se9g3zW
U9IopDOzTGgnvjnYzdrGY0s7BIgznUq7sAMl6jnBiuylV7MpxwwuplEIpUb7KuFgPQaUo6MflK93
CuaiNFR/6VZfZB0FKsXnnmiN8OTJe7Mqzp+Ox6JzBAQN+Bwret2lUFW+T7piKwT5L4SLnGXryj96
P3Kk9bBHVTImQGVTg6PFimF7wG9JJ1+lSC7OnUc2YuT8mV6mYggM+KvE508MEmGX92JjTrs7ibC/
rQk7fgg5st22SvIGug1hunSxcUItcDoMX0ADzyCmOXiPni9GPCakHYCXPmSnXGQmo52XIzdztjhS
E89JN1Fg4jR6ktd0e6N2J3JWGqq2KpCIjw2JKD/4X4Txr5aSHXmRH98A0ZW5HsYqVxzuBVsqPOXQ
qiooy57UEG5r5Q4Xb789D84C0WNOWDL4GbpsqKe8/gU72khEDyWRdgkLGNeJas0LN8p2+qch7dwV
hvBppjxo3ip6qCB/ICR2XkwkAk3zlbKediWvAN+pA4JwoWaLsVtX7riRTD650FKH1k+ACkFzMLBL
DwTPDCiZTucoqkWzTkx44WU6F7EDP8Qj9FPUAdXleivIk3YX8GDVvCrvsybB9v0bhMWqTWr9Mo7o
UHwz0YJfxtZeD8aM8/pkaU3oERZZwwvWZzWI2UMW9TEsYQKTeblJLL8Qxup+opGEcMWtcusdtbbI
slmxye4LHhVl4EdTSE3m+/xdWXXUUJXCaSNU6hI2aPc3dUA9EgnIQtX41KfNwgvBnmWQM05HOKKe
gg0iLqu+C5ydfzrqWlGBed1pzHUgvgBg3RraVyunXWXrtEClOmNXqJ4Hlwko4y+xMjBg4Snp5GYw
FmZg40usrR7c/E3qtre6P1xFiv7KTSk6ZrUvofi6wkF3ABtDXLaRo227oHW6+F/HqLfaEd707W6j
AZcQ0lUX7b/Y1CvzZ6q4scq1tTI4rM7aK/w3Bmj8rU7fCevFBmWBKgpX303e19XN+aLByu4ugoz5
U1aj0tsP61oQjl8m6sUnO0DuuV+OweanK2R2u46ih1+I51W4nGsRnpvzzYyfgVMaAafamYBkejn9
g1zSegpRCqiJiz7VIpK7a+2NU5jlzs01Ku32ma4ee9WxbLsRTba/IObaCrjoysxSrp4UdkaPZq+H
jHfEZK/Rh033XIVVC/WdLu9cIOgb3SxI/ablje1W93qp+JV0KzcEt76UBD6FMMXBWqh7Xb6VgaSF
yctyPFfyfj3foayccHFWU/M7ImpM5oGYSNWZYsYE3JmPaXiP6CVxmaLsaaGn+ioAw4m7T5s4a6Bi
1K/7iA+CBW3jaw1vF+7Vn1ELBs5aulWBM3nOpcGsyn7uEIooRXMD0cPfkbyAVph8ZyDUrFInTJaa
EBkYj6uKMaOFCeDUALJmQ/QR/3bTpaS9OahXRYTvVWrTKyk3TfFyIuqE9pKs434XaQoO2ZS0fG5I
R8PxDO2u5h0L/x/Fy/Ke74nhXHChqofpeEXfKEe9+U36PiYORaiRJLUTIiYDim/9iwUbPI0FIhFu
I8Ewu8baXJVpqK+aAccGJ+gjX99ZyquH9ojYeRuWds3XNIwH5R/Ox62/YU5GQv4PApvFHUO+avC+
yq05olAHZyUxEgosanx+wdf5eu5igEoN0D/GqSxM9yqCCsxyUmDTQ8smsKxISwkRO2EPaYvK/PFw
b7RKqJtsnq74BrWWuqU3ogXE+1J8yas6ex82nVloEXdshus/sGfucIpo34eenyMFZbZw86LOvlrG
hkm4k1E/VpA14TyjOR8mrs6KQbLophN3qLAR89DWCE+FwLCvhWjzX+n2pX8HK936/H/20HfJP1gx
jL7ITmKBTjPA17zdyWrtH2uYeXwghlXLQlgzcV08cFcYZB3j9KTeHQcvA2g1ilIJB9LDFXzUnpeZ
aPcSd/hsQ9haXSokAYaxwSA5i5skfXOOyXMNgH+XIdJXZZmceTrU7q9DaDXWgUsW6jNhrhOhU7AV
zSG5t7WhJc/sEmKjxKXZgUoky08MfbJC6wNXUrOkDOQdXcfL6WHIKECrYZpRX+eQHnYhD0JT4U5h
eCl0e2ViwYRtn2M6Gmg1TZhHYqW+tSZWhYtYPm79EjvwOFOWypjZK/tGCWrI4Iu8di0f2U6g6xqP
5mL1FKqcK11ZQuP73PzTTm+1kixyci0h+LprlznZsqGiaWKTCS8amofBygMj6U9nnL+ry40FUcmU
QGDc0+eiPgXBcGEDuJ8pydTsBEP5h/KizWhiAcA8VTCFGlCp3+EYEc6RT6/Ou1Ccsh+q0oRPRSKB
tw96/CefYd3QDLcSyJ9/jmtw88DuyYs7SHEYVeq7c4XDRHPw2hm/Y+rUT8d6LUBDAuqnlwmSlToo
DXugNMAFhUqLCHo1vTT+8TmIBuRQR75vMySVBx8LqYnpuUuKUVkZEH5w19VrliSlVolC1yWmD+Er
aHJqqmd6erbdR+dpV0/7p58ymIOUCu7UzpmSBWt2RFgCOFmX68NHAnKdWG1R//x6lLJG7QyGFePR
3JNZPCsBLrGdOIFsGI8KDDUmCZnACpkzKoY5GozIeSiMZsMvDEAY9tvWpqMb2/mA4kpDFvTeaBjp
lrJTDTxy9LdxvrExEOGmniXBWtuioA8kP0wa3OsMWg4dvQcYxPNKTH/Bhe13qtsQMAW0vk4i/DRI
MXBrriylQdYTLGahS6c1rc/0tJ9W+oqu7wkqCQjQ+/XonzAwL6/uL99wh6GW0q1mMEW2VLh3PlfB
rA/qTqyb6Sl1lCR7f+KERyVV8BtpyYcYuAc64PB8N/jIM492Ixct5sOT92AQ/c1uqz6HOCMF3GZ1
ZK1x80YRQPBtTmz+jvQHa8WcGPsl50U07lOxKSMkTeKGa6n9/JpJMvpAcpePNxYm2AtDE2457oZW
S6jhNiLBVN+ttR0j7cM2h3tOm/W6DjshxvnJULlvvO753S2LDCAoJsxEsKd+iTD3aFof9ldaDhuq
sUe3w6uuENCR/z66PkNITObCEhWK0dB/loH/y7YLkcJ12YLYdbsecJSXXX+ES7mgGsX7B4EeLNVw
aYnwey1PO3T/sCp6HpEqnsuwLL/1+nlU3S+0oHQQ5fV2PmGI8ek1FSoJMrTm0zfEK/IcvjixqumV
RuQFVxTOINBTDT5BkMdES66Y1a1nMeedILPSWuzEKcqvPq1OhR330q9+LG6TfM0GcZNGtK4qJ5ch
4RolTck89SC/1zu/Dv1uK1o2kvb62Ovj5NSz8HH727yM/RlO4HaqCluLKaTr0hsNBZTyH5ShdvgY
slBwKcV43KqQhnrInMA8cWYCrQCzyCrAgRDNK1GEzeMRCxBvXwMo2PGFRUGSVpBFVj8pN2KtFhdC
LzVBMAjaYLJQwtqtH6ey7rbV9XRJ4Yt5qJwnqxuF1zn/0EACy3w39FuqQzXPk61jffKyrCfoSMKA
ffcc5WOsn/kGTG6e9kWIyMHW82zF4KYls6JuCrxZHf1KmWtsgJYLkDDWLWz9nONP7+fgasikoRNR
ytPXtn/LSnlCLdaZIaFGR/v4LIOQNEE3Fww31Aqi1hbdFKY1LrywffGOR3zXF6lFn/JpSSoXCPzr
yvDZxGR5apCWuboulQgbDvrtfVoBraef7iwHnIJxyTKuNSUc6JrmIbYVFwLTUMdT8MXdQi3VIOBM
fjWrxdZYjNF6xTNOly0zuGsvdzoMqZtPwm995WcUqBH81K3z2ao9bawbN/JNKRQVFN0L5zs7rpYT
QRpOnGmZJOivXSNCxZ6j0SSPnGreSTGMpcYc4g5isqKm/VkbajpwhXo6KMM20g+phYx+aT74zeLn
6UfZuBpXxbmKkGg8qVzZ4oVUiYj0XbsXswHWk96/73JE5B8QG0SHaf6DyznNtmRf5p9XqHJBMlfv
ZchozkQtHPGieT6T/XdvzJPOfcJ9fRCEa6MUAsaz4UIIUk7Js7ABFaQuECCgww/ys7OIHE41Ejrm
s3pSQvIyiYjByaeVGG98rh+xT+Qp24cvWl107RMY0NXDffhgmSR8nXQo9Bt0tiY5zgkTtx+yE9J5
Uqvn6fb33CMZk4MfUAH1RmE020oLJiBQibZw+ga2jbKLc8YLHt06eFCvhyvcMBG2/wsWROEg3u0J
Layjj+8SChoUbeSObmI/7/4mpXPtzVZE8YvZT3vI7LrsiULRLirLWUE1u7rBM08/K8jjlKpl02ee
8JojHxj9fiqAGHNRoUSXhUCNpNEPij7eK2ka/C+znxQD+STLkkSJloJ5LeVG2vS5qDWRUEK5hjRg
vRbE4/exWUsMje0bIBSuVqW1fGg+SuSfAs+q8mzgF5W4r46KQDnX9CZgZD2iwvUqWrz2yAJIHKma
zuvXtZttwr3VjkF55ElIhhNBis/abgKFY9p1qoBCvJgoVxzAvXR8qnvxAECOz3oKuxNzF+fSHwVN
eRSSQ2ImmRLnVD3+g0//JGDLKLIIVrGKMg/vIk+HNplG3Vlkj9HD5ggqjIjKSbJmY866MksdCtg+
uNhMJwZJOEy2AMUDbn7wQiO4iuYSc32ro8kWHMtqI3GZBCrGdCH5BQnDxxPvze4kUxt74d4qPFq5
FVr/Gi6QI/xgAyh2tcdb3j6Bya1f4/9H2DX6EzqupQzJ5BUB/CUWFcEXGYCPzMpNUWTgaPkCDL0v
XrTq2Qu77kv8u5z1vjney4bL8uBM/0JsAQrpV30s05tPRApo5OYfgxOd4ch6nZge8iR6CInMfKXI
avda2U1GVQMgR9nZb4ZEisJ8gfPfZlGb/K+HTi2eybloOEgAja8GNG0suLaRUTnuVHsR3cBNIjdT
xp4pOlt+2EuzYV/jU5MYYYqY5KViiCYfYoa2LUQp7dHy7cN4u7TA7E/kGtA6wlNxQYCcpRvH62Hz
vy+3Yp3VhMav4+ytUVrzzVPraIGVgvEMdMiMZlpsuoYUY3A1DJuq7U/0+wOWDUlmogcxw1S1JFIR
GM9iTFP/xp5DvvV/3A3Uz/273X1/qNthLo+JbJ+s/oh8JIjqc9SjMU+Xh+uLQRtUb5C0+kjgGZQZ
/1qHPGJpaOTKoJQccPBjR2TieegpDRGb1qnAOUDV1b+uZZosFPlHoZJEctFY/gDwf1PlNsULT0yJ
sMr9/2VEF5+qEdCzCsNbyD3r3pT24CKoUd8YVyRf8h0PCbuwnwJX9aTyphVmtaU/7/HsVrOTbnmU
nqiUSISKp57BCzgyVbF6KdMvLNHemfJyDd90hTVmFdBP+OfLsnuXvKGse0CtcEceqEAX0Uw2dEw9
9IvFdZDJxEemtbumB7b2JI1EMGmb6yuf4Hq3Wou/CG51Z7oF2N3H5icn9QqnBaWJw40W9hXO1YSx
tP2UQSr0TiHpWH1+lVuofcf/58UuIGS16V9bKu/80OzueHeDTYE54ajAIAWoygr7HNNgLISGaxEJ
WepLpMwECkVSXFypfZH2SPbbl3vdaQPl7bZx3A/me1W7uZFk9tfLqQxAjaeEbZzkOS1wyN81WeoD
kUOXYrqhxetMjL9EXBIcf+0+NJIWu2wWx++ocmJkz6MLSLJ3wdjUgpgPOvjy7dpgA1YNknVoR7FW
0P4/DzSzkrbe0NCuyP3Yx3G51Wn2ceUJ4590VTdZdOOFFuwZHsckzn/K5RUZfsCiCYCtvt1ZhuRG
VwtIuPh0hqw2HyTmfLq9S2Fu89KTc8Y+OII48ceHQ0JA2pceeq8hgLxhQeLDMnq/5CroLipIKWEe
COIwpS2hCGgHgWuVxrrzy5asCVifyEI98nVq/5bV1f6vl0PEQJaohXt0jJFTLt1kKeiYvSarUfH4
o9GUuZ32H1aA7p5gch6Qm5CA/7NGltyE9Vk14hfu2ZKaW8i83P9cls3zn7HoMFo1Z9eGhkWtUrnt
3fPMg+b1awulJ5SfWea1LsEwp8d6LTL+XY+Q4AEAkMFUEOhjJNq5rP4yXAbwXSgcqMm5Xd5tIpYV
fPpPEtALkiB2pDr2x1xF10CMVBcvE4rrf0pUY6Xf79bqC+jwB2H1CBdL/lrrQ++8EGZzgZFU47KL
WcToTL12qWH8FBp6778IIXP+iIUdmf32DzE2H1QDqMWLLpJupqREhRZMBC7gyMXp3UYPt5ZuGJ6/
ov/fQwXBpHP+ihIxMa6oW1MrW32Wiy2/hiqitNOEZHC2iGBan9jxBD5trJDJC4Xpp27X9uSMW4be
Lv9haWJMLQrmp1FYu6wxmF4aSeBiHlCH5v/9ADWa6rNUzzRpkkiIwLYHPVt8zIBHjKBhC4QJHVgL
fk2ZaxYDIvJpqLZfLgFWuaPoIW1W4rBHRZq7c8EoEyBmNEJFwo/iOkJFlSSPACGv846lMpdrRkTm
/RK8TGoT+CBU/iPya1YAo/Z1lPEmRmCpC1FAAsBwxcpb08X7MKmLRW7fjdKTSiadZ29CyrJR9S3s
di2S7IgY9mvL1QUE+m+X97Drfw4UjjCacXMaT2NIpNjcM6Szu4aexEVgdTDPevKXRqFT1Z8kqa/I
Klhv+MRjT313RnRlCSMmNF+FxWgcRl0TNQLjaWPI9ejwRrCUtM+Bv9WYN7X2cpBbY/BG5h5pQxIb
uCbTd5jlUjO0uICHkwziJnHaoIdr77rTuJQgavqUBQq4DW87Y89bzSWBjs3q5t2/f4o9Y8ZCnH3O
akxv75VYdC1sA3v1xB4K1KvMQVa2QoSIOZ95Iir2bqOYWWWvobWI36V1g8qsXZCWQDsxJuC8ZHne
QAVy+3due+1byur/SHIzjHdZ+iHSzzFwbUw1gZYI2S7RWaDM2UjUrYUGmZm2onPPrP4BUZwnN9ZP
vQupci8BexxUaMJfxwia0VLAfZz0h4OjpITVqVROd5KTEVPKYqTqN4VI0w9T8rWyjL5k9+fzKkLV
WJV0Qu/fvK1W8WvVnFZu0KfMJXHbvCD1enxcPeQRaQYgvQem7Vi5WGXQilIRoesRh7d1p9ZxNeDk
VYlW8cJ5gbinPhyeoCf07j0b/jHBQKTL9AlgXsPkcQToiYmQDDYBqes7sZH7CZDgWQnNQviaknXe
oZ3nBB+EYa3ZGDW02hfxOU8YEHfsnuOPOMrYLRMbAHwHl/qnoMeTAToFswmM8kJqr5sWqYRbHkH8
NYV1LYFtCyIUHzMHd/qpLyUrsgEM2utLA1h2iQzzZUDza+sAa/kl4SIrsmSC9qH7WaCVKhE93VCN
maAEyqzSgi34o99algiwWjWxA0aYu5KEUW74ad1+dLYZWkHSiuYy15j16oUnhQXVEc729YmK3UYg
+uBuaEqbb7iBMNYdh6Y2DZXhem3YXV3Rg2U4qnV7EUib+iI5PGVKmeHc8YJGMrKnQpVt9xj+hej8
gNAwvMd5+/jn3Szdcsav1ux0/kzvQbuFgXx0Gw8Psj6aer0ABfRlEwXuI3BtzGDbsKtLn0jvfBYr
DU5j0YH8ljoPkl9xR8JJka6lZvC/5VoTRexCWHSw/MNfkNwmwVPjksciycTUlMiMq+D6wS0RITJc
9ySY5yfHtITpBsj8nK9nY3OinA1X/h0W9fTD8WvD3eum/i0wy/+WgoYsPXr3lJAC79Zhjl0TxPRo
p2Y2W+bzeQELxDsTl/x69EVT/tJcfGkXevidCL0saNGbeSHnbhnzKYsK9gdSR9tFLN7Mqwc1DBCA
yD//GbT5b0Irbj+OybYM/ZA57+fGXCHbos6WY0KnAhzowAylfcD2GmwAMUMNqrVx3oOPz5ri5w84
aoNTDBX7idsZgvSQEHUeCmzWh5iN8x6U+V1u1iFsW+iJ9xUciOd+fvoa8UDjJlqNsHViRwXis3lU
rOhbRgIWetMSxjcIrxkzSPPjVnI7bxvcEgr4JHA16EFJZCeUmLN8XWpmt5+GryQZvOgQQPG3vhPE
N6egvckm8h+j5E/Zf4vv6pbXTSmMOz7XMoYTddVZvrc8sFIcwc87tmPC+ze1xIspM1qHPSrjP9jf
S4Hf84XNfBHTs1fGdXOPdMlPGPf3HLVi6bHacn5KUyB97B6+3h9j4RPkILGNcekl8SVLHO50y8f7
fjw0WL5RgU5U2fBkdYPVUu02OvRLcKxOK7m9zBPhLrL3j72CPe3N7xyAr+K2n8a3W5f3OWIUHjBg
grpq+WSFqVz67j2SK5HcXaJ/E+hMiphvUXZddwga2MbRvhF3hes7JS1Svr6ywv52YvfNPS6b0Y99
0vpQlxr9Dyt6MI6HcOk1ck6G3+i9q06fg2LmWi26NRgjCIC78wFiHEL401djtGuPe6J/n7lAH+hf
5YTZlLbC1VLvgSE1eNsuM4u+AT6UDeBdl3+gOd3+jkDQsHhls+9jVd9U0tk0eWW774SW8PXBU/P+
/DLM0vZ52onziUq5ocGduVR/Rnxo5fbH39jZ3YFmPsZfS9ZMdlrlL+4ez7X2wXqD1xsAkxBId2S+
4S0kAH64W4BAEqfScnq+PzSayCvj+zY7DCBHiN5Q+2SumHULWQnKb3vIP/CfOo8RAJ8O6D7YiLDI
d6+9Wja373Um7YEnD8UueaJ2Oi3TIc2MJZY4TpVCpQc4lHqtC0zsuOe4M+VDsTQBcS80vLbNenfq
29hdmx9DNhHhKLzdlr2GnzEAczRQL/GXO1e/hJhkdItyRp34lFU+FWDqOHc/Oln3c/xSIkNznYpu
iCfyad49l0lqN4yl/dUKljBJOMPzXds0A0smHcG8Z1tBiJY8Kr8ZiJP/AWYN6DxWU+6XQyjy4BOf
MfI7m2u6MPABw8RyF31XnZsoH37Tp02xN1t+ZVQxol5cDUTfOTS3FnY1+hVWj1XjlI+cGnlXqfG1
cmA6TKjvb8EtAEno/iCdDig1/b0Wk966cGM3jalsJZVoiF4Wwd74CJPahY82AErKQXPi25Yr3CXi
yMSylX9MMfzzF4HOdzEGRnwtBbWRRrrTmgWtxQK2kWx4nCnLWZKe12lu+8lhQ3ey34mXPx7N9j0Q
5Lq7BxiB6qrA3O0sR1mwsVplJKv8oyR0ggeWG5NR4E5wx+W1qZlrziq8E2Fsf7Nl+Ix89QJc2VC0
MeOlaCEaEXfms0zP+S96r9M/HkmfmijPTfLMtv40X+VGyG9U3xXx727STINtPr0POMxMU/STOjtc
xNix0jbgdCndU0IrBGttP2Pn37yFy6Y8O4mUSA8KJzeHL0EdMbJpMchCM2XtvvCE/ZfPGD1qcRoP
Vm7jSbNwMPlHfiqhgvu4vnhzdDsh+gKb4itg8OLzzlWY1v4znO0VYJOGINSMnyyZvQAfDQDvBn8K
ONTKuVj1XG9ATNQ1BXe+FA43ZD8YxlM7Xlrqj9cyzgvB0hf8OsItrljPwLHg46uyU4YrphSbsopk
RJ5lgdwlvtEfeYawMWxdwW8C8q/ZtUqLgOnMhKcTk6XpV3gkq6BGSVuYQ6pVmKmOiHqZV7pWVlRc
nRxXM1KFKUmfPugJWaBsRrbOxliZ1G/kReog/wR9UYQzSCBVcmQ7vkM+ZKL7/Zk8221kbA40N5Dz
6PSIu2vdnAK+8Pg2gcKzp4WmUKNj5TfrFokEGAB2hWzdrSdlc79XcRh3eayRnm92Vz91qEmkSNZx
stZ3ZJINDDr6YD1NG1sMljnxXx6+KUQ5AAQyUmVlR82fqatBkx8mmLmZlNqQ5ggUp4LLW5m0smv+
pnfr9IiL4dBuBWy2wRXcMjYTi8DK8nmuz2DdwPnw+pjWD8g635cWYHLZYBXd0tLv9L2W2Sanz8i2
cg2L44wEmXFGTfK+maeg9CL71bciYTaMQMYSAr0EvQxrfXGMZXMCyyxMGyrf4iV61/5+ZuHkkee+
XR4tVa85qXF6qqa4sUoKTH/qtyrlnvnkPihJy9usc2RAdLerGIORmbMm44SCloffmNyJTUHOUIKm
Qm68Yf6ztRQNNDEhZZvdL71WpFi2bbPAb70uCQynyr/MHr5mphF8Q/tvEH/flO9SB4Q1kZhS0Lys
NU7VQyRAlCCTd7sI5LN3U4o28JRdh8lnythcpZRmOYqBf8ewgCA0jqJho4GMzs+VnSzy88m480Fd
o7rBy9ES3nxNbQnKWwDw5xDUDdaoDS1U0mdD9rstF74ywJ/pDjDJjnHBeUii5m8lo4RaPcdWhutF
76wDvNMG6DwR84QUDoBG8142GIFy752fs9VwG/A8Vo9+DUlqHUiL3Mqu1sYOlfbJk0NoSLHCxzIj
2ftC6uYC1SncEU0U9aWgzfys8/R86vkeOvXhC5w7P/LDAiEbBn47jt0cUPtkVRThly6XDaqniE1R
UvPkWWlIzNaNlqmAFrZwGQHawyVBZ6G1yLEc8khhU+EyM/Wth3NfFKMfKJr1pBl/7ENll7TM4Ky5
TxdFtym1Hlu2mx3XUhhJLT4afm6Q0u4BTwNiQU4TM7ZrzzyuFiTD7jh3WByS1ysix4LL5ivKj5nN
ABS9gmgDT/nczpiUNEwtt29mtlfLqWfZIv+x1f36NDVjRbH/C7HuTvkt6fWEMRhtQTGfWCcZkkBz
I+sLoZpGtCwKkmpQTXY3XcJ1fxHFZBE9YPFmrEWW4M/M0rlApf4ywuGyGpZ19c8QMPOIvcRPiWeD
o2U5ytd1Q2diKmoXVFvVFl97MB2Y9s6X3eBoiM0LOpuzujWsytK9fYAZS/vyaP7fLYtrj2/2cf4T
4DclAeqL0YhOWHOezdS3sXjt+SvKTEjGWYMhFk6wKncXH7WbNPwakfjAanE7C95ZjlhJ0DBnlNvE
6NwQd2ltv1udinIHgveix3bsTt3XMo+i12UBxw52kPuHpt+13y48Z1KHQtlLKRdCw5KBRqlRHUPL
nX9l/yQj0A5zEH50YKRnWwxEjj/qhRre+M186QGO/KJG9/FaSEl4M0ZTjm62HYeBrzCu0Z9Q7t71
XIbaWhx2FekEZUVwM4aKNbVqFmlIhhhu9mhLeRPTrWJRGT123etdh6E4vL3uRJ1fNwDVRTZBdydZ
08CvK37vuZoURgBuUyItT14LncadeCKm1Zis8B9a5oaFomQHXysqiPmYZU4QF6Jaa8VP0o3pznlV
H3xc28AM7zW0mOmbmQACq4fa5qNLCTxanKvV1LiS0SrMont8h4jiZG2rU8YKUXmsp8v92SC3gcQw
nZLV+l24wuoEsasIery7QK15e9QkSa+VLbyHgc4zObycUo+qjQT1BGz1tswuBal6R4who3Z6wqDD
w4+c0b3Fp5SZzpXy2FRA3gkhzpHhcw1R/6WSeL5KXJs6nDW1bfhUkzLuJS+zE6aPgfZJVtkJXbgi
oUunPXv8uOgzZQHMd93DgjtBgxITb+jHEq1PKjZmq3fVAYkkb1G4PfHg6NMg2nSiGLDLxLtCRprO
QCIePWzmVmJPgHO3U3lRhk5LS4QaMW8vS02nhqrbJdIgOUoyNZQV2EdKM7A2l9jF9GZzaCCDnLxZ
IIxwxcp31x5itDaxwyUNBhaJq3tRunWws2M0lbh4YXAwIifEdonAMXuBlFcmG380GuVHSYfKmR2w
zF424Um6RjbVFgHIHlyIiNEuUEZHTwu3AY0uKzcMPeK/PzknSCkDuoiYvtCtD3lJl5F4Uej7oLJ9
veqxrudDjXZT2n+pd+GbzndLnLe1O5jhdB/V1KMxgzsFYbRP9jqZPsKlVjdkFhAv13qLnmpvaHeu
ccMuujFB2OwJ0/zUEGeHXoaQCItqp2hPbCK9U2L/QXvLkpFLnkuSOMmMeQQD53iCYzXvS+PV0/Sy
essE1+OW1oQnVfEGg2glPCfuCvESihsDkwN7E1w1IuI0FpL/polJdEgG9unabElnPnqMt1y/1B3+
Kn+gUfZnpq8Gec/eBxOVyylroWImyR+U8bND8ftD8jZHavb+UK90G9uGL5zNTsW9Vhmv8V0o78op
K8lmD71Fn/ixTzP5IBn6ngelfKAUv0UZ39Rr51qxcDmZzB39SCFkQWwU9k/O7kCnP7TigaRMmR1s
DMyarxDTKaH2XFVhZlC8qHDeCSM9uKN5GIDS/wTHickTbjQ9lOc1x37dvmoe/Se9CxB1VCiBO8f1
x/q7SZczT9s6wHtZqlJ9WbXwRdaBXz02SCHt3F7u3JoAH/VnMXm5hR3BacsfPO4lFmuLrk8ZGotx
tkjmZcrxnXSC+72zsfJayCRWFzgdfqj6hCJXC+Yq79HnpeCn7/RgkDNzYRYXassKTgb3iWGWndc4
8pxYQ73fryP90w3y5njWv1fnnVzm9LbAv/3XHZtM+N3XvKoubyNFZ573YIohupx3gjLr4r6BraiJ
cIiZbR10CUA7PTbopRpRChFvYK/1jESGZidZoMmgI24p41zci9wRGfISyp81IcI96dtBLZHXjLYQ
+GLSRKe302CpFN/66qwvVlny//UU029XG10fVXztDqv8qxWrqIm2CNj9MHJ11wSofe3KnlADemnj
l0e8MxFx2ZuB+tcWfZKkI/jkDZ50Mx2AdeBmGb0eKjfUzYP3STaIanSl/8G0Fv78IWZd4nOQjmqS
fgu2SQFyx/+Ot8gY0vYNmVg30ef2hPm/grwI1385CN6BIbDaQKtnb3qe10RdPV65kP/ZL1sQRjXl
gKIR029UGEoomrKwHM7SMUJteUP3gtL/oRnhdQ+3lYp5gL/vB6FM53DaTJ5BnaWb3MTPI42v6fVT
hQcZM9SETBeC1Xt2NAWAMZwb/G9PIyvhDYKdnoSWn8nrdhgLv4crY+eGKU8JKS339HAsop92e+b4
nkSifkeZ5Q++c8Cxo8zsV4e3SFi0trZ8UPbh2H5a+Uu9MSFaB+49jox6Qsn5dIv6CgHO0uIPEXBT
OHnJfGUEPJTRPTOs8W/V5vyn3yjls80bP6qzsAwgPgAKXeqern9hyAVwNyH8WtSy3P2Yqax8IDk/
dzqA76C7PX/rfRKfg5fEqqyaeMAAIvpEg2v/eMPAY8FloxchXtnP9pclDj3HhtqUeCGrWVGle7b5
2JdVWON5cWTXQOvy5xOGbtK1ZGvnRJM2KOSVdR6P4BDT59aNhzXY3pRjVU1EWY83V79VuS5Mp9PY
YabQg+zusbFwEfIcJSp/1/SrwWnTAYjQlWJ3I/KJv3UvhbMU022xAT+o+EIVcWAQa9nWRcjZo0BA
UqHw47TlX6+W3PsfbsUWbE7vfV0lXTF594g39OxmGCR7urvxCo7066vyv5kca0AneM0lcyuFWhdQ
/HmDJW44Fzh/M9nog3jBPAQ1rHipGIb4T+JoIP/4yPjKwwmkqQoXO91Gu9FEoLKKBQDYxqxBO8p4
mJSm10+0et3ckK0kk2osPx6kCV1sd2B1rsI1WKB6RwJvY0x3zAXwNFII+fOowRCUXlraCv0/DkXC
l4PnsDjKkBCQU+FQuesMMOxmFqC439j5ONpsLiHZgJ6Zon+1Rzjw2t9/UmqEuEmLJ7Mcda4COIA9
+MLMkNz2cIRhaPnNFzr3E+kZTd+dviL5ghfcfLCr3TZL3mT8CWVxysxC1gOFMJvnFmCI/4M8JZFT
xnEFqpka8k1eirTfqn9CjF2RvpJ63w3aDDsE7abenTkQFs0qeJ3Tbkd/rz7rE/WHXs9tiT85Z51j
lYWW4H/PRvFnZzvFg1ttt9ynJhoStsahIfZS9jdU05cD/Inz95/IUnPhB6OyjzvmA/4GKqAObxML
c2vtV9BSIcYLNyG9ymy5UCrAIdDMzlnAViNL57UI2MBC77/ftO2YVL+gUlmZSLs3x9ROu5wLxCQf
ghLYZDaexb/OgfQeHO33C0upHtHL42Ntgh0mJ7yCEpKCuDFbnSquWvf7D9Fe+T/894lC6gcDeNvY
nmMS8mqYzgoFEZexvDTDplFopmitkaCF20mKfyOjT3d0AoOfdaLv2CknnFFQibYWnJkX2bCGFHLB
J0gXPztN2oqizxGxYcHeswjL7p5gppHrcvKa3ryqvPtjcX42rUt/xClh4DnBPMSYzAHDw4ljxvOt
mkq69EwaZY4YElmw95xYfUFCoRWp3HHyNJmvp8DBmiImczh/6A9PpOIh9B7Hb2bCBmxqjJ6Fkqn8
lIq4q8LLPokwxlPu2gtpw1iOSSQhpRkJbNunB9a1M5C8OpztazRw3nqBX/ZBSTsL32MmtzTQ3jDd
Qd+HZ5iiMGVTe02qsExBBus+mjI//W9FaYG245+7wylwtv4B8z6t/4nvDP67lC5fQMmliNhvHhNu
viJinXhmEJvPTVgugwQnVxVueRQ3QvoyaK45L1s60CflT1Rjh9FP8LTlJbyWe2431TmMg0BZScHT
OO0k3hPmyqtj++OqlJ9eDls0wyVv0NLVomqo1NDLSAVMze5c7xIqfaObbRjPuoEmHwqolZwOHy1B
eVJX7Aq9qFBmF1r0ydyNGXC4sTILphzHEM0T/13L7h7gV3Lv/hy6CvaLmzI00JI/MWLuIlEO/4B3
NvLATNxWQD8uJ5pcM4hFpif7J/ShOSr2y9/C6jHJ8UUxk4sk6hkUzMXk7yH40o8v/KHo8it+8BvG
i58m/GuN41TFqg3priM/Fgnf/20+xFKuUeZwEAOspxImegRyRfrXEco3JHNzaCJOtNR+F5MpMaFC
M+NQTEDC2D6lAdmFot6l3W8VMydNecRPVoff33W6Tuy9jbYwrLa3RbpKXulhGGIdceS9XelpTccq
xGV72yWCStZbXTWPgJIB9JOYCs13V+2h44Z6I7ADUZs4tgt6bgD9nZswUb5XZbVOiFilTGqOpVhv
3QGhO8BiUHw5HLzdfMMymgmeiai4ewMwk+4yaLcTUebgckW1zGlLfbWqKpxlXhci/xfKBE+XDezp
xCUtyWpvb6xjlrZs363Z6Ny3wj3sBT4Vogxm7QYbrH5GqkQ7JdykOGEjs9+kjVRPxOV5gGPOl0iz
JhIZqcMSBunoQgIQaF7XbisUQD+IIAAc6m/2Rxk/VLEdAXTQfqb5z4Id1U96tROxmA40iJEIuEPW
WYRIDI7C1SwmlxCc0B0+c+SNOlitz39s14lg57IECkrlDNM+X0ofjVB0b7kik6S9UlaV/VHh4/ot
M6/fKvVFFA9BLFJYGSHuo1t1GmOVvOogZZe4Brb69a3b8LtcIByZ/NnxGcOh1SXkSRWZukgIO4D4
WIL/q0ObjgiVzKN2hENf3XF6THolPe3tobRYT/B43i3ejjqw4fSyH+Pfh9m/5aGrKulvWchkNRcc
8IpbACocq6IBXbk+FU04b+blkLiE7crQzEZ2pi+nGDRgE3MT2xab6miWola+Uhq+EwfYsEfD9xQ4
AfW7OQARvbCn2SHRh/zPqFEfoyUmEwY+6ZweNrXIOHuO1e6NeTRjL3umsBVmpzTPM4J9zCwTrdY/
ePPQ3b9sQzf++WfbqDStzrzMk2eaymtnVJQVonzkdQroQQCzUameSE16UKi7UHlkIqQyhsLhOKmz
6N0eRLMpl76Is0Khfz/xjTAls8vYOq/rEV/1Cxsklf/xnQQCsIvdiabdcXUkPk7I+rRW28FzRUBS
R9jzyV2oqRmXJNvVABph82rAIUaB22ii/dmobu3j1bXjFRsHX96gV66n0jT+ZA2D0LNh7mLfAZ6u
dsKCVg/trn7U/fXxv1VE41NaL+0YuS2ZBY4LoRFCXdX2JaexMcx12Mgjg91WYp0RiIIIuPpGb7Lm
NiBXcpPILCPT4QkSkCoGhKUa43eYYZFnNI3I4eM6QdnNZKP+4CFFyRpWT2tgeJ8YYWwnhlfWJjr3
5E+GDXM7rTVfnT0668obYfYGoeR/lUxFAUzT1kcyfUBy6Tc6JjTbQllpqTc2iCP02LWZl2djb/l0
rXNfFhc/PcBp/GT27uXi0iZlYKPxjAntkpIpBykoRP/ibbmm0PG7zBXGmJhXnPztb6DAj3m7+E2T
J3Trikm6KWXmpzOZbov6jxlop59h6PSJ+fW4aKxsxrypqiTnQL0j5BDOdoWJml2DTrktYS9TOTmR
VOAhefs8fChD6+2KhfxspZQt5PpGyXFewc63Z1W9WtRmdEtcPwGRhpsPmCrJtNjpqwQjbV6xyK/2
NFQ+qGElEmpnstIn9jEPg2arLvQBBsLt4GK/W8XMQVA07oRIYtkQcuapb6kOsX92qXlyGNpCfjf4
d4Z8fzZVZTIYeRM8srhj4h4PDT9Rf6yEp2zaFo/fRii3tqy/yUTs0lPrydtKyLhkAgOx3H/ldgGV
hZRiGHrHJXr5k1YfApxi8wSDzdug70d0LPdPvf6VyXpsrJ3Q5lB1nC7RqSY8/9CGbasePJTrOU1z
ZBtoiRux+aZ7EvCEApvckICcdLGLuz4ZN8xEWiNiJsoaX/P1x21iaLftJ8wIayi7JZCpLZ9yNrXs
B/7i07ARWyFgvrXDYk1hvqyn5pgFUcPAsrKFpZmlYzXpWGpBm9JpxGJbixonibKWSuMTsnGCLzSg
q0b6vyJdxTFSrlGcAbo43jUnyHL1IDWjOLGU7Uok4POL3wFmJyv5pIMZgM8X4SAOJLIMSsujhL5U
iwm0+JSkeAwHVU698r8PvujB50SnU5XQ5TyQNi+1NQvSGg4PXTbT9XnpH7ql2j0fo5E9qC0PsMNS
4I13dM5Uag9EjZwJpHgf7+h3JfCm4ZpHP7ds5WdmX206jbmkj1Y1Tjm8KAu0iWOgyWFi+5Zx79yJ
cX5m2Ghn/rjPe9iEZ6592lhX5+94//KH+iwIeZWOWdmzFpnJbK2l6fGYfdBhC77/vLZc+F6/H1qW
DJX8cT9pho0aq4YbUmaULK39ECIP7ethBgNezF2budSICRsy/jFwlfDUTZjwuwkZJRNsffdccccv
G9s7YonG8WcF9HwTxVr3/mre8PowVf4WQ0DDOJOc5Qfg+NW4d6+r2fRWfCGJR2duGNSzOPzYiOmN
zwY7OM4wOndTL/+lVpPveu/p6YlRdjl9M5oCiVH6gnM5XpRarBzPWbBrzc+ra7dC3E5trz4xhng/
gwGFJtkw9TjH9WKxO5902ihq/dd4Q1WC/dC5oIYgXM5wzpBKPyXW64cgP4BgeNOTwIj0kib1h5cH
N1LeDbkxJ+lzfyPVg0m00YfmjtPcDpDZWumqGydufYH82VrM8BSAyR/DCN1FocRneSnTiki0kJNQ
2OUyr5UDpNXVDOvXPOsh7Bn2+J2kpuQ0jao9oGEB411H+bzPJo7W0rtLvH/7l6TIZWTKLzNMjvh7
JQINGgZXTJ049srCv678vXoD8G3JyrqxY/f6pP9FaYmJc/GShABNNADFDoXJ3E+AQqyuJ/f9NULN
kzxtDSmdzCXYY69fxwc4K+qFh/ffd1S03kMAGybIQfImjNrK2Rr2uNTxctuZrfppBTxicl6Vt6m2
K7gykPwZZaRme6w3GGIPA63QodsHLmIKx3Vwh7eRDqPSPkXTEEqx2B4lNCXQFXnaXkZgW0fYaKYm
lMU+RqgGQhrKWqxk42C9xl5JnEhhstJAEGqFZHyl61IqZcIuGYK4rbpcLwAcPs2T3LycYpsvA/zf
ycWIxuyGqvzGJybr3Us9Z4V9OSiq0S/fGPq/5tzOQ71dGVRv7vds9fUWzKq4kz/qIl3+LE8Op3+d
5TH2jRpruu4vcqANdVgI7pbmqoeSB4Tw53SD7iWDbN8Q3dTRbNQiFP3Plu7gpIsjwReGz4WURDMq
tx0ZpmzzVaZrKz8pqSHTIosKmWM3lR5KXEri+BVBheJgUdxvisPGNUdT7++JxN4L3BRAw9p9nv/C
zW3CDviNoBGK4qXzUQLLCDrsTnhJMDKer+W5i26SOzEvMrD6wv0cJrlk7iao2JN2XJndSfkdoFNa
Lr7GRTIvX1gyP1Q0a444rAculE+lSLAHCZYYPMVg4FefTEZyGXfaZEFuK0FCC8qFeYeyFuaucZey
IvQKuGJ2ClM01TZxnN8r1Pri52nX45doO7amchxzI9uie2pzGlVZjiGDdDE/5TkuBPQL1sMsVZEy
pfBQ2vWsD+rZTZyHr0r5edsRsV23Zf2bfPGFD/N+ZdA7wJuJxcZnUrBhWYsrQGTcBaAhpsmK/YhH
YrBBndlfr7DdGBeDzaNVa1tHnwzHjBT+vAABHIKYtnoirn5svbkn1r5w9VV7ekacbcmsaguIlPU6
xfyB+pzdKh/CbHGe/yZAmj1b2QrB98liQ6wjnhUJwEMksrfGc4WYjam5wSEQsLJRCotneklR3VYZ
JWEHtpJSKF537tmVIHIwykpBwfXf3EhvMPBNlE9XO+U9wsOYHfUl2aCg1sBCeQL0+DMsVm/hLXuq
oNv3ldukD+FmKpC0PVgQNfhlRiDUaUFAHBrKRY4hSRaTm3pvG0MTWsiOWOzdCe+DkQRl3QndCnuH
MWoeihGPj/VxX5VQVq/eHEeY8T9pFYnrl+gK4/R5ti4Pqz2xs5y510CKU3oNeMbyenAN1wJknYp4
j3SmI7SfeEu9D475BIhCKgrMSTaywwm3StJtZg2wPEgihluhojx/IzFrhUecdF+5B34guMWtpmZ7
9sfOsIK+gx4jgkvvkBu8laRhl+db4x0mrg0V4jRhgd3icQzRhGegQF8mV3+yKKgxsdl2Z4YAVC1w
FYeYMERemkn/sdHt0HV9uWllKdJ4/OP9tAsZjLXFftXkMjFkGkcvvIYXnIDsXnRzDXEkP6iAalQE
KVKPwNK+bZaKlHmY31XghRWksgFr5QKhHlDGJbCKwaoy1UWF3oc6NbuoigzSCBeiJbs7KZbITPCN
qhhdw1QsxlZ7xLbqk2RXlBILZGR85ctF4CRSXCU3gzuyiU6lS7NfKR0vR4O5QZL8AsmvoXBz1poY
ahNIRJtN6lpxr7RLsd1oXg5k3m/Z6KM+3NJUV6VS1cLgwUyNT7lq3tjgk9dRTwlWNpyoSPbAt4jD
mHWFIFsmtuYnff1ipe8M7PrcAz06NUbthBc88VXRr0qutkIuaYBGKStHolAgiu3Y6DpyjaV7LOro
p/xj0t/D0NFXognb0ceRHxQrX4vqgdjPpZ1kRNdmD7Vei0W1WDdN/mmqVOHIMewu43bun5Qdq92J
P4WNd+whj2EmEJzbEmxCUHiL5Tg8I6rjZJZIaA8ORtifdy/TXd2J+mtdDPOYn3RZAp3EpEJOPjJo
RD39Zk1FKC5MA8aqhZ9BF6f0hJSo7FTWDjtD7zKMwmWbzYChH9AjDQTeFQWLCaNdsRUPgx1u9/eW
lP+8q1eY3PHcXjWYME35bG5Vr7YG0Ebnlh0RRZLJqxuCXoBL5MqeFPkgDgTlqJzf+stTFGNk5RTC
9q0ccmrH03klFx1ViCCccBlu5OAN+I2wecHAV/aTcJ9e1yX1skM7mdJhvGcL1fguhAczE1JceTD1
cGE93uMqXuGSD90QtwSrAgTz+QIpuEyshuy++Ta035KgXs/7ECX/wCAT5PbTTorKjZFMxrqz2vdv
P9AElk9PWH+qP0p3KeQw6gr0Mc4uub3M822VBX/pxBxXe8I0DSIjyehzk0SUdyOpojMDQ8KWFgot
3f69RFfH5Zy1CLtjmakso7OoVXTdYsfZmNFpvOrnL3gjvzGKnN2Y8tLtE8bEJGYMOUI+HihkJdjV
yEl/693l28vpgjfvDCSGtcyrrMNnbCLuU0TV4CoKJpHL9hEfoBrO0830KTePn0xSVFRs4E/WjnQc
KlAsVNi0FseqnadGAAsH4t85Zaz09hbdpZg8Z+ix+dSjLwPrGvMT/AFHO1q/mG0jUPc3L1zEu4Ly
xFwu9m+fH6rbc42z5Zf1zRVmtsatwmnJC732j6wHQkAhVdp2j3wmRGnfEABmhME0g9i1sTuZgC2m
a8ixSkLBkDwFBesw2NVwSQihQrglF+ALWX572I0yRig0EuTno3qImJD8a+ldHU4dYxxmAVzFtU84
1P3tNWJmbtUnnIcfbinFpqGnj19qIxgRAukej41WNwnneZ4yXXSFyY6GRiCt3SVlIyPF/qsz2gOc
Kfq/dhHvEGTZpozw8CLnJMOsaOLqmAnLBxpJKyYZPRdWXlZAWRtcLUxSyJzUD+3Ul++cAb4G3E6p
nfNlMJVppac6rc88qGzOJ8zdDlCgBTJc4PQ8xI+4qWYQs2H7IwdOvDo9hFEXKIuEzEXls1lCu/uR
+g14nMsquYnxMQLV9wfDHq2ytF1damaGDBxnYxkZdF5Qt0BMigszgXC91RIJbS9dsDW1qP839Ug3
jTWDnuD+QqoApJLCWiU/uvz77Xt2krnGBaCi7kfCDTCc1mBxbEMiD25Ok1K6O9ZAE7m2q31clej7
xSoBaBBGVEbHa+boQ8eZcoD3npvWzwAzYfk2HMei77TxoNV/Ghg/l6P5eTGaCJrx55bcQF44byeJ
ad0Oj/gZhm8T/iYNZPhNShxDZzji4qLy7ZukMHmkYoxcYyd8h+WsKE/pvOgP4oJIsMrB4yb9pJfe
AhsCjCCImHkjIlDx9jkxzfjpfKkrDBVMHDI3SOZfDFUfLkC6Js+qQanAl139twoTNoE9Lh97BU3V
f4Rn2JsjqgHCCxqAmxj0QGjHbu/PmdDX/xqhhAOhAdG9/SrfW8+YIPzcPB+qUcpT7YwH4pWr8DeO
XGdYmYY6ZCTQyM8HUOvg34zHkoC4Y7LUMqh/6sdekL3rTGkxg9tFLQQis0S7sfoAIysIMRlEwVjX
qWABtMvh3li1HML72oXoPVBLI5CubOA439KU6WaPkF1mFzOqqsybMGul8Hx0ubm0RquwK4tse25s
dLi6GTTtlBhovAT1wzLIH3hmJjhWHZ0VXzQLlz8Fz2QzIN6tpoSWcN3nHNTYqLd9obNAJZxImAUD
aYwYs9pZ0iVDgLIWddUqWMs7W1s9yR3X4hA8PHEPMI8rq059QlVfnwG1t6FfzafeIBY5AXpvSHTo
uZNcv6xzsgeUSGxpaFNG48K7jfnNz5olbfnSTlPZCvMHkadoCwt6stkSMxxHAnvV5y7dgDTKhNJk
iaDQ6fQ0UnnvkCupQx5WWeOK3vofxD9YbA+K/U3Q8d9RMfQHk6ULng70lWJ5ybzYffaw2RVjkLvz
J0iA626EnM4P7NlUyzx1W6huabMSwWrqrCocYZcVy7CWdiAnTy/LtmuOLfY9r86dEXRPM60Uo6K6
fQ/Q5GK5mbwNz+N4qb/TJ521BylyvfYx0Js5U2kLF+IfT6blpgdNNIG30vIrdhaOitnxbbqfm1te
XLuA/SwUlYBsj+nLYKnUlKuWyiQR6oOjB/NHEec6E2nf0bs95X2t21YSVbJgBDIzxdRHr2zIFaj/
xQ8uKbd805rhqwWOtYGfQiB7eCV/kreyx2Hw0o0SIUYAStCwK57/KtgohcTPVhAZfQU+koxyzNsq
3L37/l4qhcZqftCRX91tFhe3KVaQGQXdZ1tPlNU4Tp8npl85onyeUZfQKvKbbpFAAUoRefKtQtFu
G68SzEu/4YfunSEnA+UxIH0gsIIz+SaBBdattrgHi5XAWCqdEWjfbKqfL1WhSvfv+OUX6Uqv5A9h
/aj8+CdtO5Aql8W1X6L+T/IEui7edC39paiV/fRwkxTV337qCNrRkpEH3l1P7uLNv7AogdZVv0kC
3pLYur+hM8Zw4wrOJ2lg3ZufN8mN4rmYBZAc2VRJ+FSehIpBMHSvuczEov5qb2kwElr4lh1uKUvC
kkl3SB8Iinygwgq+x9BckOBquAnNxrGaA9JHTs8VTZDNRZDL0YYZFmMNmB3L1LWKsnA+dMmjKAZy
BUnVlKPl9AoXYIL4jEEx/sZB7UlGYPojlS92Y6nGA5wAOu0/VsuDmTcugw9toM71O/rBWq1f1EhR
p8wAXAb75IxoTlGSLbrfPwqZrdT1VKa2szz6HFDISZvjAptvYd/KWCJoo1EjVKDUyI0W46EMuobW
KbomAeGLFglvfJIMAiKqYLqAszh2Puq+nsIjrXIuQspbcT2hWPwSdiLhyrFlokwlMoP+LEh46UBA
1KuAhXe+OJfZChvgxhRYLIByabio23d8kVeJzTzgfifrwdv1boQDtc6zIs7MUI8L0tTMJFVhNnFz
JsSb32yZALImRPYT2FBLVZXp0OBQcM+m8/XMk12coQJB31lKSibikIkezV7kuNcfb0T62hW5NA+w
RieuwK3OvVOf7N+WPgD3098kTVWg05kajk3djGG/WS8QcICKCKsbvX1UFhTFdmvTQ/4LSChUv9jW
ymr9JOlUxBhhMia3+2gcjm6pJb0lag0LIbC6BawT8qChnBDvj6+1lAhFsieCrpUDLyTu2KLKZUX4
ZSRC2xbX+wiOm0UzsAvzem59SKYfgMd3Uc6dtfLeh0nHHSqsf/MPjfO7S3tqviHwe6y2HDjdTjjH
3rwnAhCtMDsjKo40ujSiWJ526GK1GIopeKz6tQxC2wQ/U+Z7xhdW1aN1KRQwKyCa0JPIv6A957FD
Y4RdJg/n6g3NJKZ2NNJzXcY6NrF/5tmjY4G2xo3v55QXfxhJFxEpWcUFpo619AOxcAyqmGrG7Fnb
DO8ETsDjRWapwX60ZfBDbiSudJ/soZTYq765THTdog9Vc38ZuBM6nTRCZsB4l+Thu4Rz+JFYJbul
BWI8QErHwXcqq3feV8u0aMG2vWaVRrd/KlVuqfuaCw/yxo8xuzNP18JAe/S6kX2oLF3+U2Y353Pi
my9H8H49FCI/9yl/EY6+BEzgfry53FhbLoWoe6txky/Q8kY+4V5EW+VRzaN2O1scK36yRicCrD7d
dgBky/1mDH/l/ohU3727kM4kqStpt4rP1eK0Q3e1TiB4s8DAztqqOaYcDtuKtWRcK63f+TkWWjEA
HiP4W+ly9DFAx/NWGdWVw3u8PSbR+b+w1OsH+1C+1kfdvQ8GsbKb/eQwuqFRp34J3VqS9bAYvp8D
NBOVbsqGNsN76gz2ENnHx0jG37mAxR52CIYK4AlPKix4jAS1Y7XyXokJDU3rokoL6EkAEP/UZy6a
AIzfw/NDzt8aHIJfCJCBS8I8QaIxBINXeXjRaN0DIT3amb3DQ5/VJnc7s4mdFYI0Hkf1rTZSRMng
REBVDRP/w6eisuCjAaJxyybcJpnnbVFMGGcRg0iet+GRmHCXMjYMUYL4Yb8hdSiyJweIs0hwx1w9
cp9PiJGozn63EJrirS339D0RboJSk1fCE2MiI9r9TrHS2dvdHfnGAlbBqZvOvH6AKHE5rLeWb1QL
51h8XYFDB/cvmV2OhWQiDgPTSudG9g0/Z4AUD6cg1H0mg9agReADXH8PjBDzsT6IpW4d+Ndzpklz
BlYTyJ/d/gozbZVKyzK4nY9K+HRoZjUrJfc7AuP54Cx7nEv5VC4fArxZPg/vf3na09YUpT+/zlXh
Guu4M6m+D+5hyw48sr6DM9RaK+w2jBKSevZcNhxo0Qy96jsYV+gRlczQuU7aF/S7DtSaiD5oL6iH
ip+M7Na7RjrIoQ1g7tWFJXtnYxD7h3UWMKoFlH68ALmHgL9DWnxQwwClkiyZHWrw/Il+BGOqC0rt
OvKuRQtisGMBg/EqioJ7DKVCbFqHL4IYTUzBn5BhGlPfdrkBZNyFP3kQyqz9bp5roTcrfenuW/1M
2rVSlx/S2ZMN03ySh3pfwMBf+3KYXYc/9q/dpXzJ66zENjFvKmHJ4hW5VxGWcRWBf/cRLZ23zcQc
eV99DdBk9Npl70We850O2HnxHUbL5FI37rF0Zbd1J8a7ZwHPzUaysLeBTR3gWrwgbO3igci4Bqzz
9euPCRNCePSwreYq4h+clRJ0/1VlZmFGPqINkuxt7QHgBPpCG9aUGdnZO/MBcMAGFMIh1/gH7+Bm
Itxmp45ilvpTZOl98+W4C9Lo03+hm9bqCiuH7ir2rUDVwQFHrWvDJsWRhKx5p4o9s1R+uP49kaJ8
M2wlAf1YT1Vqkw4FKZLVeaNG5XhlxiSEcxSkWWSRQBCFzQNXV03ca0EaDogGUTYJ+toJffe0zlEI
jK1Isgnow0r0eYA5hW4omvolvB9umL8gG939SffYV0EVuSCeE44t8ayfTOzlj4Xlx9bmwzFhfwRA
D8Ggyx6HOfgT8QXU0MrWX2MqxQQW+JVRFEPwaW6DeNXbaSmtDGQLmU7HuQCwdtiT/yK2d5vAdrjq
XXUZdOkP+FbDfJxKFb0auhnKZ8uzIaZI5yqolEQcIN4S6nvDEfF5oMZHr1JAaStRECC+/Dvov/fj
Df3Dl2cp8VLkJxi+l0sFWl4dCrVJG3WTG4PUaqqc6Vdz6uA4dxRPrjmOQNGQ9sdOKxd+SWK5Mz1i
Z9tofdNrBauqQUAJ3rfBAbF/xnByF+2PGn+yAnolXB8KH2ZaS/FwwdsCAE4gxxe08nuzqOkLiHis
lf3fLUgvgOVEejeolpI2z9ii8aIINVh8a3lSi4cZbNJYh25lsNgJZNpuRc224ASZhVctCXh9yM9K
qPC0KHp78hVjCIwrc5+iR9xKdGrckRuXosAAR7+sue3NJGaDAZXpEvB3j6kl8o3DUbVfR0Jc6ifw
Bo7MpLRKv8dz7RQTm8HywGdpCLIjp6JhvtphugC8mRbrkdOX7kPv6QabBUdLh9RIxjLfoy9xuDTX
v5yfAKUmvL9KPvt9+6N6ZZncaPr6Pg3FgbNHUc1MxgbUOEmWOUiVrjzNJ66uwxeLSgzI457IF5/l
IFRXisXSRrmaghwoA+NZQsMYFl4o63SDMrMyu4iJ4Yin8JJtHgDGVT5hccrDNXyaYn5sUw/eBK4s
LPvIeaQ2MLIbePXFmMw8MM4KB7yBoPNa2T2dnDqQS4ZtegTqn1pnfcVLxkpdR3+hAynP823njj6J
kK2x/QfPDmNRzYfcOY7BPs9UOuGsmBM4Tv3DJpNTZKPOLyPkkxkNf8zKnXdxVI0wBB8Olasrcl1E
kV++OH0NVCpzjsxX4YErA7Nt/jH6nkra9QO18b4EVjx9mDjAyUifC1APE8k7n8sJwQPNpGkEkZqh
WoiFiVeI7Smn4+pHPvKDmXEzeLYktGKHjRKjsvVUzgavSYYdgXd6HWP7nIysXMmTMomgWGBFYuaD
4iOz2mrBDrgAzFX1fE3IDURHQrf33PhNnRcnpUX8xyekMSn4/ywqBn8RyUDpTls5+NpCyfaWVRbg
LgIbLo4PNTNKSuy/A659NSpnPDCVt8P82hEeDdukZs0WflpwsQRRGfvsWitcIHoOXCu8FE2I/IUJ
nGV0OEZWlMhq/qv7mUEdF3mLHZOBvon0AEef5Ze7HBvgw/IGkv96DHPu59MQT/iKcTqK552nsse5
Z+SGLHiT/HLIdfScPFp2Wvdo/suOLHlI48Zkr4NHFTt8lDJti0/PShOu0cai950c9XuQgvIFMTOx
PEoNXo7hT1GfDkPK7a2096/UF5+c+xOacJ1e8I+duOiS3OiQ/gaVAS5fRvFo2jM2iCFquudUPsxf
f1+B/JAWRqYF0EKEw+qBaoVrvUrDm3h1qU5Oh2qelgBSs9mjQIpmBqkjt/nuMREVNqChOa7W51XZ
oJRuPsAo0TTmmKVgtxpliJSUTztr6fBk3yFeePgRUFrAcDPgJ7jDP44L45BcpYrVaC584c/0znq1
4AkuEbRJvVXnHn8bKO/iAgwOMW9veQbNnKCrbkf3mXJhkPkxVbWKyVYwNnlfsJFaw5HD2LDfTbK9
DnfgKbcv/lclZvHivol5T0elsLCjQ2tq8goWST3+EOe4EKkMRLrczXENEq+gFelT1zPyiivwrBWd
ooj9hTAgpi3FcCL+UOgXOj3JB/UmE8aXABEObFXBwDbefxldLRqQeZbvWjTi2M+DsayXTXJvU3HT
ZOZAE9Elz8d1AXBXIavpNxZZA4x37fRlzOFqTd8A490fbBllMSwnM6zhYY5XCVQiurx4ajQGQsSz
e0wftKPagyUx/YLOzdFlk+Dw5RX2T09VGcTvkMt9OZAOe4Eo4t0fTennbEgFaEyGd4QHe2cYPXvI
e6YKCFhkHjmV6x9LpNZNMhIEX4CJaiPi9G+nh6bMGfytxHKxLOFDd9gy6ZbjjGCRPApMFGv1RwD+
TUvGZzQoSKBHt6ZiNCsrKC+d8F9BQ+ynpv4ZMASruXmH0kzOkbdU4I6AQH0ji4L+8rqZYmW+Iszn
xQMoYvyoXlVX5yNsjUZUudTS8iNbhinsfJPOjU1dL8gDTAYcEkSlBfQNgnsJZE9eyEJvJFGHJiIK
Mt7my9Ry4hGw0JwmN3/KdjVxzApJQRTlts+vuyfPt5XGimmNHmeuoV11sXD3rQuHJdv1AoMX6nBI
ZlXurOs8zSpSuZ8eLf3KD73ItdIjzAHXwJ1YPtlbNec1rPyMi7UfQreuS8HagH4U+tZD5FCxwEw0
LNd+WtPwf4cQDP3LCrmbZ6VM07GM9vnTVmuW+nweaADw4etras6AMFWSoo41Dkqxm+fJItxNdwZz
daGwLQDM/8r/jVByXYSbhJ4hgk4d105GLr3sKTOBFj//Hpgw+YelRux6Ak/Ed2bcIzTVkB2q5ZrL
F+3SpIFeyh6zRzpi1UAp0biJ/1OABOTGWNl2l1G/UV8lMbtp5QHLZ4lFndNLJRTO5Rs86R1OiJuO
S9n6ui06AQ089V7Ns08UBRccGAudOOm5NWUlDOm9O1x2pTkE64/sLNjY3n4eDCJ6S4HVX//jwQ7D
ByUdyUXVQ9eax2xxq8I6Kfo9Q7j0JegBO/YkshcU6EKRVxV5d1XxWmZHlsbecP7Os09+RhAWE4S7
h767SXMjoEijgurMtcLjvWOpZE8vdxxoSZlmoJqjvd2SCSpSTo9PNQguvPR8cT6lTjrpD1ZEabvy
vplLGMQEB5rG3/FSwCeZlY4yHuwG82W5/bEPqHO1EGHP6XDnAWlnRofqjdsDF2D1cvsvnooBmyMV
qR/OfJ+g9VkIzO40l04TMa9ttFE/KPCqJI6BHMzThfpFujXtxc7rGgGB+apRKCtcxoe1SGI4oJ7I
/3enJfq6sRqp57egReD9YF3V3oEaOXF/h0rLAZUqJli7Wx6lQCvf7ajACWl1SVJ37joXfC12WsLz
pIZZMMUeYmlIuGxk1Fc1SccC4s4L7NoRRsfK+VoES3oPL+nGcYj9Izkx/ZTdg6N0apqn+jGpDWD1
b5nEPVLLXaWGLfWSuJkC+LHAPxvb1QqhZ4C0E+P2vssZWLN2ftum3RRVScQkT2SVcX9N1qwM4NpM
hW3h72LC8wCHy/cD1kn6oDetg5cfCJr3Napdo5g/xuCRWCbOIB2Ufsds7l3/Zm/4s9dMBhCIqwL4
TFM+o9E7JA/s/yKUUdob4maIAhfoKJrZs9CwuX17EFbBfQfD3M/KzMzBA9d4qYY/4N3aeS3WTj4t
uB4WqBMK7AzLV6PBnxTCIjOn7bgYqlE7DSCu3+fG86UZn/eLBN0oogvdxaAY1PFRTNz7gD+do7du
zADQ/WDCbjOVwT1XmVTIT9U+ssuoAGMSAftUjB8xaCsKoInWtd6iayzjBlHhiTPPbVcqY4kXC7BA
PQzVJkMlYGryoyva1FfkLb9SxqfpHGPd/SQwqWFN8/aCl08PaEUt44jNePYdM+LINIIY3LGdvLYD
keHjEyxL1rDGjclyG1OY0UnKv+UdzI6H+fNWRVkjsvAahm/mJzY6q4atfIulIOPT9lrYOS+mu4h8
iWqdva2PR2YOm1xOHevzF1I/6LDzt3tj44VhHyChsjQKCOBaH5RT7WMV8CHh7Hkt8hyLqA8AMwKr
TJU7brwuIFxC2h4oJss5QdL/rJB9A/pIl9ixxMI67r4x6CLEuwPj4i6VbXzB/P+aOUzL6N1k/fzl
fzC6FqvaxzInpfcC7OPgiyPgFyfGGlRtShAhQiQo07UJ55HPRlR1ovbTmfBQXvsUuBxYGxMU94Xs
yFQAAxGARHdvFNl26T7kyQsWcOurcgaLEGb207Sqdal0/Ci/UgMsrcO6OT+7i9IRqFZ3YHHseQR9
IQBg5y9WB++Ify15YTcNUtmsnLFYUNEKRIlHgcqNqAKYaXqCxlOExU9BqLo+axvviiHOrdCgdgDE
R5IELXOY8CCvqrqMHrvWf3hqco1ah356y6aX5MeA0reoTAYHBmAYMmjaoZp6aovrURTwMRfWXuwS
4XrTzowL89b4wCa78avKJLJdujaAnUwIHfjwhAS4+EpkhyOk5u/eG+RxP9F/dNlGJOMQRABKVgz1
1aC4weCKYhayTx409pihKTdeB3nLPObdWMuLPx0YQtwZaAfcTAD/TRFvlD+adZE+npjA7SuM2ORu
NcCZ4Y80xb8f/AEYb/0PAlSjjjAUhNZxLF6UZHXAwGwVNKj1WDsIZvDP5tiyQgP7cLY4lclMaOCq
7AFK/MdclpLCRYUeTI6mgNYpAqsz7Y78FNzoRXLsTSOO50W2boWBfb+psyCyOr0/1i+yEVHGpv4A
KKJub5nhjw06b4KR28NHykIQlbfVgx/IjkZ/IUXCFycCFGZAfWh8vBDi9OCYisgb54657z0UUirG
3iBsNYiCI3cxIishBqeFlsEFqYy6q1k2e74NOxT8lqNxKOR2+oqKM060rbSqXFdyj2LDx4EJXUip
qSBFZ+ewNlvABVCXt1bqVVMB7Ct0fAUfNlt7GZgwYlyLDuXVibe7xOuoMhW2pqPm7ULaXanTxkBq
7vyWL4DzTqVlvC1NtBcCex/I9GQ+WXW2kS/uW1iBD3eGihznIlG1OtzxwpvPIGIkU8VtmgdPEIPV
H7wTS/j1vx6bzj4ft+7lQ91PBvWguGpcCy8e95tADnaCaCqhcvmEPVwZ2A5Mg47JKWxq8Vsvy2G1
qHwHfbl/sJ/YeNNIGltZILRJna/ZFxXEOrYjOH+i9HL2jABEnhQp1AFJIqeyHchFjBu6MO0qIQge
xmuA2yuFr14V0p2aowCG/dqIT1MyK26IQqV8lXilVHEzEP7v/GnNcMNqlXhoPEmNo3iqw5VzWdjh
c2vyLmmzgcuZyUMGu3T8j6nTd9hPy8bFX20dyuAf4rm611v4FYs1hWMb5DT+3eQJQkaMTLgkpi0d
wnUMj7AKTM+XvwFaE1y4gkvbvaCjHrGuaFEh2jjqS9WRm0l2q2vL6acWsfazev9x6QvesX1j2jGG
gVlZL4FmwAYkrdp78BOVlOyXkOX2xgJWg58m/63+PiOInGNwfc77AtV7WTuQHQNcVaUGOGAd99nf
iHNEdGLH5QQ2TevrjCbqZ75o4fDZStFw/1V61mVXkY4ep1786o20Ej5durDQBh7nyrTP/0N3n57+
3r+Z3OfVLy+PyWLzs6s5cvcSByv4rYXXHjnVfim67Xi+xAamigIbCpQldodPCL+Lor4C7OJV1c68
M6arCfF67swnAIbNfrOoSdvRfxxVgo4DbRCzYVtw2LXKcS1XxtUMlEWVHhWX2Z525lc4VoNUVP1t
W4WAJQqeE336cVJOaCEwJIkk3tUR9wX1hPk4RtXX3mh1RwtstEPv0rt/bgI9G1IeDB7HTP+O6A94
dCTbzBWucH4+bln1FbddrQTORxKKApYLTigY3ioh7ikTfawFm+X6cImwEfz0/HFU4Sn8usChUmM4
VdIKV87QsiMvaUS5geyvya24p6oTBqitwRdfOm5sBH+zBCG8/peDN0Do836sJHmPYAF6zrg7dK5K
kWVViS+sOVgDmRNRi0DgNggk9djGISsqMMRd4gr2pqDgCmOeXbfJOkGsHVI/CO+1rQ/fxGhO1Nf7
/abuqywkC8GubQ5tyUjYhMNVSxZrLA63M/rkGjSj/A2HWWlRcLd+w0v5iKq4nM7lKNSif9SMjhxV
VjMDaJDJLKquFiBifEZziRxufc2GGerr+t2gF7FlF5NBiMKun+eXwP3yb3oXbTx4PDjgzVIoa08a
wkUW9yDpurkMieTp1DQQr4huloYvY6yLRCULjgiI5fR6g8rbT9zv/GRomGItoMETccYOxY1D39hG
TxcQu1aiRrXnPFL+QptZoS8wfUIgGE89cYvE76SV9ahyUbxdhahhqOs9Wijz4eefvGHawRPD1MwE
kruc4zgJpSk/eBziDXs+xz1vYYrNm5UFVe74xgu+cJxc/WpGpop+PYOhZt07T8f2rJ6iR73DhdEU
MBrQAfeyM7BSimfNS0A2ffKChTsLhxfQ6uEaIFD24BNqDlQz8N47fi4qGt8zSMAlIe+qJhSJsTJY
rtPYAwYqpZDQnBJoRVrXg8o5Matuodr5PV0snAVa9P9GEuAg7WbwR+Q5kLmS/MehMHjwNsUHQ0D+
eGrPj56PNJ2BanZk7/aVWoQti/2n5QHDOLpfkaEwuSmuNMTv7d3o/AwdNESMEg0VvB08S5Jk6oJ/
XQMlfU9c2AhdRJR0ITVtkePYaZcFpKpEZwspPzhBECkaFniyoFwETog3TdI94+QfkMpJorNXinHt
ricfWm8DBQavaFcWVg5oUaNJs1eY3lGYZq/WuSpB8Hcz3UORn1nXstK4IcMBtah/Ugr+1tDHzAG6
XT1CtK4uXikj5H76c7C3PvK0jS7wcFq+tE1Cti1GEz0833wWgtV0rb/4tkA9WDXskR4XvniHUsna
mq/1iunl5ei3Gg5QreA8Ze4bSDcGkN747iy4/yGF8vhNqIoaLRUZzO47FsVezPPvwp+9zUNTNqcq
DCGmztJDCbwqYinqI78cWawAn8sM8bYffWuQJpT4ke5GtiXFB7R0etyFH8U4ofN0r8VpfrP4lyhn
Uj/qyVjq0Ar/zOolIGBzOuFP5hp+7q6yovmR982OhT0loqCnWKc1frH7upsrGXN3idN9ZtrK9DkS
NzWHOy+P8dRU01KrlXtI0BCRdx1FRJYv/KiCtL7WKFdHINepJmPC0ImZY2v/iPjTf3gKHD00Dt9L
u2r91z9Xc1WnAZKxQn0B0n8po3okIcbFgpOg82905Q+1wYUsI//tO70Fp4yHJH/vh2B2zsqkFmBx
twTF69xibppnwW5XlQGWNyIAFKACURCFcORBOts2DDGJJExZkTcLb6uPfes4o8FhDN21C9k7JwxB
lKlbLEeCcCvpc6/DSxvkwDxcxF1/KAJxW1VF3mZTO1HsEV6zntFeeObpLO3VTi0u3x4EfIyTbJXQ
v8Us6p3gM5qQiVUGSUYK1NKHzG5XavGGtvoXLJwh/t7HSR25egcWjLQseYAazPqj2rI4Dtcr8zGO
j47Nf7DgQsV9x8a229K82I7LpDHrlLrvuuCM6J9ZkCm5CnsgsOHF+9oCFHzwhEbwxS7MIRwM5xNW
Xt037fB/jm2bLiG0fuRxAY8c0VJ1IsTjIxkrrwQDQh+zpoLVTyeOaDlzTbIt1IQ8bL3Sb31yv0ac
6Jgq+RPqZk3Xcy+pYQrea6JvIuAvXm/+e6eaSt1yv4ogIEHuRxjfRN7gdTXXFGvxdbqcHha9jDhn
HDQ1CUiU+cKB4lznCrngaJ7vgCFAyds4y1ZwO4f3wA+B9bx2tGaBMOGXalXHDZM+SGyGgGoYlbat
4UPUhWfukupNpj7HOoaxO8+NYYKxxplHaIf6W+LxFV4WiAeW4iu+BqD3tZUbOP/yi0o4OUPnqzdR
K2/UXqJ+itarlj4xkpq/DTzAEczjxDQOZQnWMaynKpOrixNOa5PXulYo9L9EO5W4+M4ZGzzeuAGL
g/JyeofOb7/HEY8U7Yb6G6cn8FcMT7U6Cg/kbUgFwsbQv1dJ8q2l1ITIWKnfdNzsJOoOmh4XdBVI
prESrxCXFozBOW6oynBX8UfDtscr8PFvO2RlNCqIRM+3lT2RbNZqJbrkpPwIl0RfOOoOrG9EFXXI
O8VQWh6ndoxU0EJapiwJQJqogKSTyFlJAS65HMorJFez9BcyKBjdZbHjfcT1AevrQEFkvLC8gKZG
aFXjAsqGh4EuGWk4BeI/gLLvGwNpHFOyPImwDP+V83pHnpouN58Gi6PH8YUnq2aipYakVTHOYYfV
NnCbc+6lHfT/JaQqFRGOKvxzADWfETqa5+Z3LgS0N4ALohOtBUQcz3ar8gIsmHEfLMtIPwHSsUtm
XXjKroNJSMZ43DafjvD5ST08f37Ew55T7GDzrcv71DpTW+PgifHn1BRuBj9tD6uzbP3jM47GfcKK
SPJUeSkKMzJQx4V+pTfAKmF8M48hMnnMeF/xmSS/cgpFUx6eupGC1ppS/0JNTG4FBtiAB4O0YG5A
b7eP2osATPnPCgdtHfzMnsDh5yXGw8RGPfwUZZLRMOvNbJk/b2gf9mvdNSp3RBKinSH0kuwxNLtI
/2ahrdMhnRC8TaeZ2EF+pE0HcF/iTv43b5rDvWxmIl2BvmvqN55j9JIcqBNEWJDJEzx7rvGey/2S
LWgXvT7BpD/eK0J6SF7aEkleFfK2BgISiY5e/dg1kVfGH1kGAZ/ie0pl4sOwpqyZAOPK8689FnMB
LAjz/MMAHUuY+lc9DHMzFY3NFmvIaFkVAwIvJ0pI2PzkJvU98XcqbMvXDgvfEJmWxCfrleGFNFi1
j9f3z1s1Gb13etUMBwdnQNYUXXxP+85H2ymzkFcquzMp3uO9yXNR+0RsGbRnUBsHInSamDFz2+FC
lD/aqsXqbwiuJqgJZHx6Z4uCBBYef3jvRQZOAc4Vrn1H3/UcqFMJNAkXT2UhPYe8VsnFNUFnZjsO
CaOLYO5KjCdnc7d4jUwC/DMbpNEUEcyqDjXQKi/mbwUzzX2r8nh20PHrlF9uKErQYVuKnmOj3yDa
usB2u79mh2swmlOxxrbEGc6hR5pkiFwV1UwxFl2eDbg4N4GdgbkCGrFvVFotOmLgEAeCUP6+fWZ5
8nBdZLRBhzUTx+Q1fXeu1DiC6RyPtdEt3+kcl+hsKDQYkf1feFKZANW5MGhWWRNlBv4qytihgUkj
8IVsbpbOpJv9JkqEG3QFj/TygWDxjYeISzPpDOs+P+vxFEmHb/i4EH4I+fh/eNNdVsNdW9rbhWtV
LS6SDSEeAn9P1+bDt7/ajxwNQNxaXqB3XoPJhG8xJ50upe9IcscSAjrmyZApyj+bUXHl/iwIM6Zy
iN3gYO4aKhIAXIobK1V1jpB2Sd9m+cRvJjKFHyp7+MkZcx5M5CXSKUFIpWBDjbuFm62Y6aHBdqF/
YzuA3+v+Otc7ueC1c+6JKCnD8NDKXxumFD0pgYOu5wDkDVIc7K+uap1vbtjKaLQThfVjTbGqx7xJ
e/OwCLyTA3komGKU3XLGGu2GoUHxUD2JnRwJPYefTDWU01izdy+9QLTRwJIFD5IBeHwxyOIaouXy
VrR1OfuWMlKcyokqMrl61HhZagloxTY/zjHnB61eU8aAiKev3IJA9hPkWqluIWFGH1p5B/3t235i
q3N/JriY3OKcVh5Tzdsc1ORW3TsuTcpdR99ijiVpzI2ytdEwSkpUCbnlnGwIgC0wne8YLJTZIwIp
bWzsWeQWeXPy2459hY/2z48ZBm2RY3RpyZhCbOyaayTy7W/dLoDVwI8vZce/lWS0kFI254dhZgez
3yEGmym5iUZNL/fWSYR0TcweViJUydcAQTN4Km9Yhp8wd1WhQfdtu4zk+007k5DiFofG3jcHdqp5
IwRduzZ8B3GMqAPJRe1PWtqM8t+iXyFH92JHSppscr4vINLIh9gb608oRh7nWwF0XUeVDGu1qnNI
JaEAcznAU1Fjgw7AALSPR44jWxvsGXXtmxm4QPkbspAEW6m3PFsff9LSKM5Ogpg+13GUF11+Cjoz
SlVjxM5l5VVaN8C2ZFuafY5VNpSXSuVqcX7zBIgb0bB7kRcW0hL0bKverN6FkwEbPcoqXw0RE/b2
/la6/mgCHxrMN+ZCDGd+KSp/L53J89IZpCKEtVEt2xalrxLxCbIxT6HebOKDGadgpX3UWFQAgv+R
2jIhX+T9IS79utDb7Fn1gDzvbvUUHa3nbDtqiP8u4rqYhdXo2wrMNV4JsnYfPHTJKg/Lpjwo66gc
JvjjXi8u3H5Xt+43FuNHZtyHH881VW23tsZvUk32qrie5ta68an+M3HyNHHPcdOxFx9nPckzSGLi
8cPjtxWAHalEatkwCgk10svhX4Wm8zfmK8JxhhgwDB3X79JBIzw7W9jEzsy0IvM9eJbOo6wibRpY
df1CerekMNqwdHvwtY1WrHBSbFgFVw6ZEYMfhCGxV+5Up/x/oBggZLWld77WdYAhB/sn6un4h7Bb
qf1LfuKA8WD9Py9iyNq5rMgKnTwgCg1ZGZl1UJ2ACRkoQd3i7Y/PTa9Z/gCXxRYrlT2iLyrDXJ4Q
widl45p77ttsKuqlCWpCqjJwxPEpwhUI+eDUg+s1n5bgPsDNrX/6lGHDuFO9FK6bvoS9mqyQxSaz
+m9udtapaM0UAyTLocxSdKYF6o3/TXkc1ZgnH3vdFMKq89vkFPcPiP9ZYy9DpVDEN7pMBlGXNHZ9
Uys3U2Rin4vRtvGgmjxoKIk8lKlvQRmOAnFjyHQuCJzNzaBU4DTP0D3FI/HJghibhajIHEHNIJVX
dN/4HVJ6RdBgFI+KPxx9XLAlRnqlOm1kCg3y4ZApbYSg3yY3DlhOjer6T/Y+mhorCPQWXRXot33n
0USDTEIF+2ey5RIxDiJ3S2wzlYSHEiKCerUsrLkAuulvxlny02lFesZ/l7cp75pHyfh35e41aR6A
3mQfw6NM60egNHfAIjBj7FvMOFpNxEsjlIVYvy8U1ksOZbqL7SLSc89y+gr7s7oq6kDjkCsNmfl1
XZJWMuKOaAFGlBKS+/Mw03Aa+nAxaa3RmBrx42Iugs9RwSW8uNwCl6GMJi7d/+5mppLZAqB8ocWh
WPe0ulK5dDetUPm40AHLMnnumiBQsuLRUePKNQlg3mcpy1vwzW60Yz4tFppnK2cHo+PT8yAQKGN2
8Ymkfavm2BV1j5JACV9hXY5d+lyFCKWeIqxa+lC6/g/RVuodRtZCbh4FOP+MK0sNOo607rEgtDn+
VxBfP/4C3IdM1f7OYmNMFOc49qEXCQmi2mIjqdRRPPGflhOoEim12UHxaIhCKEHhzoXYTSH/aO9Q
9dLJwBxWtLLCzW7C1QtjwJCvco0zYeu4GCjEZuJAMstsMjdAZCDaQvzGiZbQHrbpb0ODV4zQKdze
Gqisi5JgE86o3okJ2Vut5kISNmRMvj4/11XIxo848/dM7dnKiQ3lv+GckyIS9ZR6fQySiwfX3Z0f
XRV52vOils/kuagS8bf7QBnxWQ9ft9XlCEC7wl/OUB6GcAp8ADG4rYi8O28KnWopx0xduTCJtSb2
KHyAIhF2ybUEaLUl5Z6EqbGbMFTxOIOMP9AykYR9qxl76ahlxvmGFqZeLxuT3rbbuMBJuxG0JnpF
jazKQbJRQNL1AeH9pim/1bs5vFER0dnmeBBHSYub4tihxG/40G72TcT/8iRXsQMG5hHWoNbcktbH
jyE66uU8mfnM/s9svL+Dhu+8Ot7J10wtkjtkw97Xrt/nrIRWop/guhAgYm5UhTY6nVh0y0usJ3jL
9WVlJ6cvlZ2o1QhK9N/v/dBV+ffK2dxTOvCEGNUfBjhKIrfDbIS9GaiUsjVGi/xi2OkX1+dnJtH5
bVpjpyhrwp5OXlErtWfGzmi5XJZ/CwoFbEFI8IlrIWKbCFDLoVBifHYZCMZhIBjBtaFSH+1u/9hv
zNXXnqYaOw5R98S5OkIn+uoSEAHpwRjEM3lO4b339MSlqe8oz7hLjCeg1IIKcwD19OSKuDmIMqMp
gD+vlJ/MBrmO2UpUj5jILef5O38hMj4sH5pbVhisOXqEHYgajg9i2XM8iX6wXlaobsDJ+LKxkVNZ
YJJu8Xb6Nx1d4LAl4BK9PPVVVRdRcKd1KfrM+M8nIKGQocMjIuBVnL466wMkc+IkpPzvZ3tIAoFZ
eX7gw1OC0KiH6SNJsIsBXYLJxtMju+i2XRxfKG+h9xxYRKtw0HNBPecs6SDXmWU58ohu4dfzlMbO
SLCGpoyUwAIqrDqtb4znvNJcPt+/rtd+0BmUIp8Art59on9ldduWHMmo6rRB2C7HEZUOvKVW8I3G
78qvbGYnYZrqxLTd9NsUBU4mBTL5h6bnuCJb8mMwCBjN8Ao1F6E8uV/5QN/7mVEQSI7tMAt57j+y
03OVPpt+BKGfDsyqhznZ5hdTeyMO5Ax1+vgF9xfJVzsQrM0pwisEi9Jjz3woSojxnQtONyA8l+5E
uP7fLkp81b4TYEYqYefwge40xq+HJjykM85gvnZ9giA+HAEF+BgcGyJn6L70AfjkaatIvos5bDZ+
Gntt+8XQBeSKC1CWaBmnfxkx6I9O7E6vEZg8cxm/1PnFuP00VKNBHLCp49fsUIMaCshb0X8IKmPG
sizO5s8QMDsKr0XU46/FNh7XNZiRdSBDnL3v+INl+WAzDFTyW7UYGSsOkP7mISs5h+16R8NfAWTs
BIJs2n50Uu4CCvVXGDKTg+6C+qAGd7NDfTGF1v/HZX120t6HCJH3Rti7o8zp/ACOH54h/Ksw5Vht
OCEgyvYER0xdzYBKtzyIzZUW9Asi8aFa1s1lRt+OGlu/USJ/f7uPwL+lHuZTjYwmgSrRhxHs9pij
882q9bAOXMk7yyWBeXNs3rPA/nG4OaKJd/cPeXS5L/tit4CKAmUmo772XRXUOdn7V/opHSnkcH0f
Kx554Plbwa5YpQ1LLEkC4ot25vi/haBVttgsonSe0vxbDyhl0nF1SwSr4KxBYtQ/+kb6OWb4OJBr
q+UPZ+HiWzPIo1ZbhfRGoUHYAvKZx1U1UihW2TRe1NfATDT5Xh7GPOf+/3y8YN6F5nzS0ngq+U2e
RDRnpEDBiWD215hPoxjGBZh1uslWuKhpDhJvjrnt3PQWyyt63IEl8HbOIwbUITWd4UeDHhheZVFv
IyXl3tU7nBVdG50ygvLoou6a0G3B20vPG+brm8FMb319EevDzk9R9lg5n68kUKBGw/PgfH0jbVd5
P9VmM57HWOdXwb1YPeEPUiCG7Hf4z6S5e0qZDnqnchf4eD42MOm6OQBgmv3LBKPDtfbGZppvFd0X
rgqTCFvnjFqqIZG8QxIbViGdnkQeGB1/25FgOYbfVEVUSLKL3S5T4T4Y1ERdK20XRKkpO0IaUrUj
Pwz+kPtM1HsuxmTwF+WMntNSDyyiZ18AgTehZkJQCLIxVSILnYJG6/08zB986qrXKJfbrASfgQ86
FnbgxIWOtRJuC2bQ6AI9sp551HUmR9pPyCeocIQY8v4mUWgO4XlOXelardKS6UStTsRGrnSznk7w
K4jbx8OPpeIiTrsa2qe4WcnBqwSnkxPGkDWweKulBqksNZQ3ibBg25/93tB8ubqo5snsd0UNv+Sl
m5Ur1DQpIs6yL+kZ2+qX/sD5cODoP57L4E8Y8caexfk0y1IgQQUcsj3qfr9FJ4z4lU/AK4KeoREm
YNSll6D5aaWQ0DSPq8FNRUNLmTIR7XYGPjLFv7FOzTw9dEZMxMUJ5Gc3276hQLH6tB6lDmHLie8B
L7jMM4ZaabQnf0K/uzDhcV6CI9I9UZS4+mAZ6sKA4Zgqf42JMVwz4lJ1tZmXWBZbamuyDWgAYwCZ
XZUXdnDAk9UqIRMMNzIlJFrl4GrmdXp8oRr9Fuqto9mR9eBKQNTCwLkG0+ucnSZ2/NIPZaN1Qum0
+bvPIu0/1WiMMaRg/eL8XEHeIgW287ZP06UkrphRU9qbl5ddwidOg5Oe/vgEFdKE7nKPYL/fwvpl
6xIzklMtJFMfd9lrmiNy0/7rI63T57DiGAbc7eiITaCc5Cf0UD/Efu66ay9CTj2Ai5rUiZlppolf
yxQD7QEx7Vgwczq8wPVAyXLAfl4zrvN0632CXSottOCMhv5420kTWOe7+eUp5JIQHfpaaO/y9TCd
0OMQH/YNqXfkcStylrTNgWHcGol3DpLGr/kIXJdwVbsRTTCk23UXyRWFxzsAsNd+pUNDno/DB+9s
BcN6nG0asTY42zkBMysrDnWg9enPkkPBv6DgqVYS+F5ZyLqJBUmoLvne2t9Tv41t1yCS3Z4+/TPS
TokxahlUnCUQjTjjRZ+3W76nh8v2iFmlvxF2yFx6XZP03p1Uef4UIhT1YCHlFUk5/xjNVkgXkwFU
qI13kDt3Btcr/iCrc2zUoqcQdRSRRfiRyqz9Jom8SAKMQ+VwVZx06ucr8tCX/SuJz3oUyPPj1V0b
xlino2BonQntQ9aomAFOVCLvuWx0J+4fc1fqylZx7GaQxchTHc58mUCCHovxv8gPDfCyaiKwPu2f
yywJ44RML5C2+ne90QyHLRM9pe9s3mG+wZtZtGGcVOt5wKkjjwOuTbnZAgshG1ypmX9Uj/x7clil
mbSAzxQzxuJgP+Xu7WEWd/tUtJMxXu8ra+WZEL6Rcp+KptHbpPZdX2mIkAh0R5eDerR3pTfSlahm
/c3j5GAPsd4XvcIBFMpJ9d/ZY+0CUhfYWUycVqQ+76PrGBdAmC9SkHGz7cCuRnXY5dfo5ixKgmSq
6czlc+pkrVFY6Jj2DnqKgSaJE8DwB/XuIcBjUqYolWPCQCx70iocKicHxps48NjKsPVnEiwyku14
wkeZGAHpKwtVvsX+5QmhT/AO88hGaXs9mQKIR2uVg93sw2egT5pJ2YSqKko+MbXzngPiLEK3F90E
Y6dauemjy2+IX/f5EGdYdU9SASawbO34XNoyaAKeknQqdlTGm3CncRVhLX6Elz2F23NJPd3Qed8G
0Ax8xETGzTWAM8ttfyifqVPUfN/wHLA9pLApFhJYsfsNnIBZLCktkcZ1LhrE45+xoAiVU1cusRzR
o1kl+lFgQCOO7toXsf1cxTeRQT+1AWpl42nfV7WWJbryyxuL6+KSB4Rvx9yWwUM4pf1ixNb+c0hR
fV7oZVkrjX6V1JkvlUsKZU2yJhJpKEKrEhsSL3w1l/Q8p66R/Ehou1TM4dTSBnkLOkeP/lYNUk9r
tTn/HG+lq8uCbPdv/bj4sk8CpOW5GkHK29QseK+juHd1F6jhFPIqZwcv0SbJD3lWXlQzzvcwK78u
bb3DbIYUw3K9G7cAwbxeYMb+XniQo8Dyo3ig6XeVPMFGr0nAsscXDeg+ZubEA1yR1j5OX3WZM8ym
tXXM9Uod0xaXMK6aRE6rxcZbuES0BXH4mxwdOOGNzVPPlWIjon4zZUZPiBALevUCmhDj+zF5tPUr
xZSIoOj5vsfNbDs/EGwcwptr+yVrPcqZ0VnhMtdGlS3EzHD/eiql9jnsN5EjQRuiFLrGndrjGQxt
veq50W6hpJempeLDKXHCVGDXuzpyoU6zSADqvprWOeU/bjJ3TYCdR+DkoZu8fhsFgtiiPYV3s/Ri
joiPFybZxqT61Y27FKRLWDFVJkWq11dMMZQE0p4cyFRlD9RS0epDnP2OkCkWIMSTF8dD4Tosd1mu
7pgLOSX+mAARXpKfyQqgEjymZKNCIOmuvWXohelUMpq2ixg500eIJwr7zLJixOJsibTodlv+tE+9
Nv+uF662zROv/HODwZJfnFbEnxb/Zg3Ol4OlaWUKAN/tOT/rax0NdYXb2QfKbVlloGPeqEAy4T0j
qURAoOtbEonexGRnm+5OScfymeLdSb2zaJBFBRjJ1BLN/iOJWf+wauxECzOPhlX0eqdKguGB/JgX
vxKmYbqPIWK9IMDl0min9IJXJB/i7vH2ARq+1psp5RGjDgMNRf/oVcZpthvYrhkGWoDLY1t35Ys6
E+b1b7e2bw1csJ38K5+oUhpp3B6Gxp0r2iAUNgkZrN2H8sOOXaEoANlwrCFocQqKazWogJHQ3TMA
Eag0yGAGc7WPpaP7T1hERay2peZyu7LQR9EDg83/wvkVVICRMIWXwIxszyJ0ykxDYf74X6x+DCUQ
5Q0c0Fgubg+YyX5YqFQ4UGTH8XsTUlmC/qAvLFKwJJeGuNBZMuy5keIoG0n42koforhTXeRf7Ify
CIz6mxlNIgH1AwAemvrUsEX/+VitRaT0n1tbEMGpGbeeIBeaXS1AjBUqDx+VrL5qF53Uh/cytR+J
5UcvZIE3XOo/MssUCru1f1SKXnnKHi0Ag7W52N6yMKBjtdqckwPODwnfp3FvrzaRZuoo20DMgZgr
YWEwENOWrDcg737ZZRNs/U1b0Rw9nlWm5tIyQ7h0ZsH4j/YsHe8zaK/9cYLOCwWEnD1RBvuRCFn5
+xmvfQC53HyiqRH0vtsUtri0i859YVrM7PQdxZUzJEjG5RHmCqGBmherfBiqVhpFaq/SwLfTrBKZ
DVIRzjc4eZBG17h2zKEuKmakVA7suAa/7kX3SleMnhxypzRd2pHH6WGp8BrNqFu+lUjtUhfwfkLF
4E7BDDyCkDuPtLBISX5aASvDOBJgPa7RdxanA1WEBe2A04OAPBhkJJd1AwzmZSg25QW/V/bBkv7t
nyrvPxqWV3cqW/58up/Z1UJckOnsqA6d/7CD2g21431AmXdk6C5FZgL5WrREAy2cr3vE78r+50mq
517YlHRR9fJ6eg0Si9l1LZafVEsW09DNJbm2pAT4C44Wr0hF9No2CChKoz8EFCFFlHbMgkghfzDd
Qoyd4S2mwb+Yw+/A2yb3vSSlewisRbcS6zknNqi3nPlzjOzPLPja+Qcqijbt9Z/ia2A40VGjre0d
YVrJ3EiJLYBrqKRAeAqPlbOp5PEwXgYeWZ9L24ZdU5mbd68eeCTJ85AugaQrpUiEc18Tfd8NxmBx
BhkYhKtZVA9Gd0lczo5v8M84dYoTFrrKqYuqSu/r63EMHC0c8ql0W2tVzt9XZTdsH0qh4d0JlPvE
PB0M4Kq1/A/CbHHfFHKttw3O+DZiOPtflhEEFOwejkTrOENyRqaL5Rux/I0J3x/ZfeBTXUtwkVxE
XjRyNuwf9SUISPtbog0xWyM9yuE7+VU2TWPgaXypcH/6xMpfkAa0Eg9At19l5j2RWpewPt/HA2rH
PxqvrTsKhEctcvul6/Cc59PtlFOA2EV74OlAk+czYlAG67kaMhm8+R5KXwD8NyfuE/MGHAGTPcax
9mXji/bLheW9s6tESYEx0OWAYU+exFCT2xN4uG0s+RXednRMEl3HyKlHTfwY8ut6SauK+/kl+7UW
3zGLkKJkty8iNcB3TP8DberwmvZzHrU/0vtdhj2KBSidT2LeZj7c4ZVtM5FEZftuPuT2QZH/hntm
A6T8rf2ASlSx5ZzPe5X6Xl/+PTVum+xayEz5mO28cG7yVJ6auGZCjtI1G7A297VosBSX9/ZAMsoz
lP6kAdYQIgfhvOQUuVVyTKMgvDbz7y5MYy38op1taAes8f1Iu585RMDl6n1CzCk7hBaNe3VNb3lO
8H8g54g3PLc6dm59ChNvCeSkgyLARQdm77SjER2UDLTETRKVVpghjCV/hu61nGVfEtXadbVJAgRk
p7EJ62TyJo6MZHLr0UoT7LxmHhZd92IW3lwJ+dlLONz8b51AL7alDWL4Zazcj16HA0lCmLYdPOXh
3aEcjaHI6gzo+rvy5BncSmaE8h3ZWrUVfRqGpY1qbp0T5acmZjc0dSlpPQpDIVXp7tPH3PR4ut6+
44YAnBmKckSwrobPaZmdFJWDXufrPa+wKOqLjedS8uHR6Uthkp+JyvSiQoLPj+tejp1mSlbi9U2b
6EDbCrnsNP0OeLYOSwYYtuAIviFh2fQfe0pUZ29ii2SCkXGg+djX7zpICGNbyIWqHojeKFQ1IArG
5FoMmbRfXjWiR6eWZMCPX7wTPV/QQULtyUJI4SQzm/IaV0r/+YXtVO9SIvoJ6/TWDv7sjI1PsD7z
mbLcYBfMssyfBc1IIolLiFONrXD18STvz9+lLHiStovKbab54mTw+B5RcCMD/OT4y7XpQ3MRdmiw
O1nrMJx1K5dQdORt6CZ2zfe4rU4H0khiPA549h9bNyyhWllSW00+uknp2zqkX3IH49jn2ncvgWzW
mBiyzlByQ2+EdvCEUg+Wlu9lhfE3+vJDuED4Up7Wt5c99jiIBdlatEoRrjMpHmpaB0r3JGo6kP9x
S8qErUsnBn9Jn+2jBtikBUji/1zOBMoK5087e4cwQRSgqkS+uuM5jMEZvu+vqkrDK7oT3J1pl2ES
GcpeiL/wR80Wn71jXhuCDevVc9wIvfYY+WJaulvGWP1jEAQDPQkcj9T9j/DoImCXbG6P0JZizWZL
5VSd8H6IyOwYSm0w003CjcNaq8GfrS67skuUTP5sJvP5nXw8u2xkIp85iOlk9h6Dkc0Eg+r96HDb
hFQQmjUnIIBlW0GvAKFQO2/QFjJ2i4Q1oEmwRW4c3dR8of68vZDmC57OtSZbUzLeoSTwgt59HbwB
xzoihqHZOJhJDXZHEKCOhwmF25HoiULHXE5cRKFpsMNl2ftBEM8OHpj9zciKfPuOccMtDJQx7T4o
oqsq7OR/IBcQurdvQ+9B+tB3glw0OXdLfmHrfjWr/7CT3HscwB5xN4kgJvk3q1/qqTezLLtLaGhq
MKOaV/PSVnVlLJw+envCen8nWv5OHYTlrTjU7ZdmxFyzU4wcd2vtS7kMaDBoA8B3Ss6oYM5jwH3F
G7Stz9PNrgS2PwuEAntpKF2DdbM8zbULeU1Lagb9Utv8wdi08qLn0pQ/YJZJOhs4ye08RZ5jeBOY
pZN6Y8/SScM/t45cLucME/mMd06DIIUSed7m67hylwm5W/PEBUMVMLfxxFKXYsB5KgSeufH4O1Jn
I7vMyifCJZQOpPnu8VK42iVFb+uUmrYFsXAfvSdcerNPBmjNVoMhAvNXW6emhxkXB6wnmDI3wqQv
f25h6tRGDP2TJ1oKLOzHP49VrAVE4tE0m9FhTTZuPKOHfmlTv5Xz8xgHwTgEqu2COTqwO6uPbVB7
6hIRpqKieQftHznSmBA+2OOpLozXzf+m6GY9qFwOoC7DNrmFSTr5tr+BtQEnPoX7W8izOKff+zUj
Cgd6eYYY6j9LV41W4ap/KMxqvOyJNw1ePzWulVKvQDnU6SZOoVEpB38WT4TPiSLLSW2UGhJKVby5
y17cNUmfEt9Wn7An3Vn2nWbWCZLO1Zae7QDU52G0KR8CVatVtkjkHUwvkH+fWRZETpdefALjJRRn
9wl4LUS7+FEljj4sqsT+y3yyaJLcnlB/hy4p/4FmGYfbpnaZw34aPHlW1yu6/s3DYjBHESCJ/8B8
LLwuN5SKHx/GDp0p1bFepXUB2TmzRZj0T40IKs5qLzPapz0VSIu7ZFld4EzQQpR/MIN6z4n0gvo8
OVG3X0rCfnjbtPEMGW/gQ5VZibEf53eX8SFVDwVGQWeg9FFlWFP7jos8eFPepQJoOSBoBGL7B5xH
InM+n9KkncIIC7vMB9wU4vqzp786NDIEBBJAjc9+fG6fYpG8XaoNGlazMd9GJClDQ5RyDb1I9M4k
ETj/za3ArOcQTwBB6NUxAqQhJ1slHmpK3JAcvCZKYyTUp3/DBVe4gv2vgd/zSH8EMi6M5u3vlber
PzD6aco1n14d5B68IU6Osme6cGQXV9j9+C7JNxIc32xexHKAJqHLKEnCIKh9EPUhbdV/ipqNzKPq
KI35Y/oYXKBzBrl6u5CQPKdsUp/toYitpnmg5kKPHl3w6xXpUtD7/XkarV5rYYRN8PoImra5LC/w
DbwVDeDdq8EnHSb97n0gzRoghqbW1hpzvzad4HqLSOcDdRc1x2D+vRXrVVQf5Jfrb0hIEctIT2EP
420nnuCcSTdBYgzsSTurSp5q/E3dGAWRf+3iOcI0ZzdSmIXyDXonYOtto6oRT9ORIU2rQVEiQ0n5
/Cf/0ldnZ/OCQw2t0atptdMumf1edlVghNlgeirlBXQpCtfTlskyq+aBs86NLwywz09wUXxgYjoX
7/UoP6nUPrOwzuC77WO9yqp9/G4+ZdTdIivChuqszTHmTTvSARPEeIb0CMxw3QbNLb6SyHlHhZnU
eCmyapN+OcjvJWUVEmE3PsiSV7JKuIyseOy0z0is2AwCcYKy8tkMsWVySmlgeihPRfobpIDnw3hb
sMxHOoQlSWqsWaeuCyq6FtGsX1ZwHGtt7ZeBuAw9EfS0ncCQFdBy9otBaTDo7DzakXSw1HgJXtO1
x8QBhr6ab84notn9FhjdEQR4zpYwZvfm+v4X5cu8/tOwGFqyoAGhVbBFVq7Dvp/4gANl3jhL8mXU
8LZKyL3g7VTXxfbNfEP0Axem9bYZd/7xOF8IGF6ax85OXAoVPTO9qqiYGbSevJbfNhIYrw6gef2K
rbM/zESMnNg4Cgx72Nurr9oYOxEFwTSqt6Wv1KMz6YPSO9U6WVTF67ipEVIjYUJJsi5wIIc1WXCo
kFhazH6mR+5hipOfSPBdyoi3MUbpijPy4VtGGLFqGA1bTC4lH3X76e8pv0f0AgxT7PyM8tcXU1Ij
J6Zwpn3sklrTmB828Rw6bP+qWw9wmf2E+5MKXbXFX3xKYW0tSgUzMpUtqFQ9fkg/YxrM+P33O8Rz
ZiAbyTMiXzxIAnXAjeIduGtgr8qIKwoHO3bN9cYn5gTZMJx4zBGpK4MpFhodXTWx+ufXSlGjsQVH
F+N4z2973jJNzFuAvFP7vnEgFtMROxT1SuhW5bfLIWDXb46NZHM9t78rbp4MlSYb4rcoEyiVplC1
JWGqp6JiltfLxiLaZjmyI56wvfh1mEvq7g6d/DkOZil0ZEhKyzO05uJA7EGXyEtWmUSOvmzkhO16
UUFbtmKUtl2khEcXizs7wk2F0rN/DJF742NacoFliDB1+cjb6lFkys7qspE7u30rd0adq4ZvawL1
waR8c371/wxBNDiuMyfJ4Q6CdIAguj9fj6RnAySQ7k1dPHg8B7kjUzNRwad/OEjC+QikGamjHKow
GDEAbJxUkJpfrISqpvUINM+id2L9KmLxU0T+B0THpHym8jHDslrUwpm995dO8h1hRtn4v+FgEcVf
VKAQDI9I8NrqLhdPjOjWpfRjEfZFXZDc1OhkL9kjF1z2eLR+aq/jRZ/7rw2y/q5WfJCC7+alUA2P
xvoTIhLbQQGTEUAJTHJUYj3e1yKh+WT29f6JJlVyK3dRgwdSGpW1ZXyLKofRE4JcfXDnO007/zsB
QmK+ilO8YJEoR69SNv6CbxwzJ505kocGpx55oXqgPhPcMTe6NJtEcHTfjtJyWBaekNbWMP2C/87y
w1FujaYshc3YliK6lrZedT3dwVWrRwUA4WlJiTIMIz/haUpfJJoFUo8SMmgRpee0Jvvmyi/F5zhE
P48oRGLRH7KXn6irlGaWUz2qArdHY0mBeF1NvheiYDEcj95hFBrIKDj2RvQAyqVX7F1RS3YuWuCm
E19eWUO7GjoJTPpESSD9tAyMBa+I36tL+NwdYpPnDShs0Ut6k/QrSECEsyK1sJT1CDjdQa89/sbl
2n+MjjaYaRXwXFc3owHfGVSE8Gg2+vdY5Zw+tJu/WTdPJ5K1g2c9QuC9vtl7Ay5Ux/S1XHS4lSR5
xgZFkcWHejvKGrpPTUYFqSCJXJYmeVc4tnwKDEeRbpMY/AXFFPjsPtDc0FIspqjHoNPKITzfhguP
USK5wuiZhEhVBREHm1BD0y4QksXOaYxE0h+v1GsfWEyt+taN0rlgvnN6vVAjN/EsYoBF0V0C9QH2
IgbMAZeX0TWIChSefXaWYIYFaj6Z3xcoT1TQg08OvvvkR2rZv8cXwxCugMqkSxJlG9yVBKSNJIyx
oP2POgTjll/cxu9UzfvnLOu8xkGJBTznot5Mh2nPNkUN50aKvZvjwwKSuJ7ecGr4z+JTgQg08fNT
FFlxGW16a398PARNK4+hiQarqhMHMZ72nRgWe5Zqr849k4gk8OBF9FgXyI6SzOUd9Zs+xt1cSHRA
rSqnFOetRF5/9Ql5IObRL59+4FeP9+uFrWochmwF0QL6ko8VMTtksFiZLb5qDDBx5mZKsTzl3Kyr
8UBmNthDT7byp7huQo+HNo3I8cmrJWPE2kfNrpOB03pUBARG5n1KiYd0Lf8Pt0fxNb8cSTiDvGOk
16mg9i1DKL6VXpEFShHbu9oFBZYrMFVoaSyb3n8PA1SZ0Z+25ZIRdL9jLGhhWqGu83sr1c8tqeCn
35Y6F+ow/IkshN/sXJ+QgSFBPJD57WuqmJXp8KQTB2gjZoZ8WP3Wd51Nh7QE0Vgn9gTB0WpViSz0
yHyMsb9mTzK2j48KSybRYzswUjfrYoMiVWS6siuxdF2qjaqaS7sgA6DExyvBQKnSid+Cp1CH8N+a
YU7sVvixHNhxxxAz/HZmLQfXmyBW30p2mqHpUekbT5xhChri0v5a1+kami2a8ZNEBjn7aEBNuxEP
hjbNuJIA+4VQAQkPDT7ToYr9+cERSggBFz7s7ecnqycpitMR2zLsYykPjtLvzeYMppfeNSPfXYI+
gnsg36F/slbU2JDV/ZC5ezTy3GmaBKnPKQfko0j9fmC4BZumjx+iqSln101/Ig9moHnAv8GXeo/8
DEXngfuUSDYF2ibvxfIYLh8TchWkyLrvJ6g7v8CgNLhJs3AQCqA0331nFga6Rly7HdI0I2GzNwcg
qKoZgL18nAlf8vAHO49W5D+VVR29G8bXylhCbjSZkp+FDSqnW5vki09TCDcj0E1fY5a+kmuTQI2a
0uHOwtrHooyXiaDJ0RWcAw6JXg1Cde2gCTlcvRnvWbQ9BIHJxl5Qz9XrbGxZOpVyjfC4k81qsWlX
YS6CczI8Z6URbzoEzKjQmZG9BWy6H0oUwy4dd/vdR3ba6NlCW3JeWopgURYsmERKLIBW/aLv5b+3
QdihicNk9ehtmCS9vnKCsG06A2efBP6N7+qk/gsS4+S1y6QkjcV5lzvu1ec/hSd2QQaPBFOBxP0o
sQlLhb8ZrJkTkPSYIsrUU8C2KA+XlmOub9JXkjKHkFRXQPsONAl+ebBPRgl050TKBfwT0oSFreYM
p2V3DOzvOITLLw/2w6bwAoEHtcPmAZiMMIPwIWgcVz0RD7vqmNAMY5trXNdG20e/qr23HR7DeHg+
NsTgiGjla+JVrDPYUF8iZ02dnQq9GpV655X2pzhSNtD55xh20i4qdGS+SKW6aDuWZ9hsrfcNm4cn
PR+8PEiqS5ngyNyaOnBL0Egtev+0Tn00xEjWu3OWEXHYprNjC0+wMA9D6ITiAb5OeTPaJPes7wWp
PAF5eU4HMP6pAPB4UJT5NWZfZv5lVHWTZ3iFHzrrNjrAQHnW1IJN++6YMxqj8iyX44oCVWngjoGN
q0V45VzXZcdBYpSl8UbM+yX49UyhBSZ+9A4R/qhXuBSID2WkAXOT6zgDAbVOoTXA62PEdDe8DCtl
Rp1QGPaC8TWUeOsVgt8m9qEsLAETuKiIiSTo71Wgo8tukTpwXm7l7xE/IwKAK0zieRurhwH5mRuw
00OctlD7bdaOAhAalUHVw+E5PgHv57vY7dweLrZy5nklAS5Xj/ET57hS+W1pQDKnl3qLaFAwvx8Z
+wOlWD4ykFR0QtnORjEbRnq2z2n/cmGY7rAIk7V02lvhAULerIqt8U82kpMAYMVlXy5gH4zK2Q+R
CC1PDqIrM0T4cJ9+tyPZXt5fs54YseZGXIr0SKcrRWG4efht5CNTQst8am4lbZOEvxrb9Q64bnWp
yIvsU0RYKoeag323XFBeWq8v2sZ8qEVUQQt15zmGlR+3e2vhWpaS+dz2+I4RX8uFxR2vM9MV7mSY
1i9UQGxpB3M8UnpZOIq6qUMLF4gkdoRQ6Rg4cxOXvL2WzYu7IX0n7kiaJieAEamu6t+5I/gVJeaU
el9Fmgt8aJ/C55leX7q9qIhX18r7k8F76rg3H4QFk3rJ1xMJ63l5DE7Y0EXwnJzTZNmXV5/MO8Wf
QjyVHdSFUwz85XgNgeTClx7gRr8qcQZ3KDEMVZNrgWIaE5sjBaenQvbrAJg80nvyix1OPtw2O1cC
RLHTYtrTZgzdWZEBpiYS/8AxiE4zmzeuNhr2xCKV/Wjtk3/Io1kCPfpSYJZ5J0iHLjle7zO8Xw5S
B9qDVuXkHTFdhozASmWCozZtDy5/vex9iOpz6IRjJahMyyGMbRxJkvXkcU2AMgcbOJz+/2Q/AfjM
6w5bqi4EZZV3UPrY3vdb82CfmAP5beP96H+jBcuPh1CJz475k57Bm3Cnuf+zc50eFQ/2z5Y0OBEQ
Xbr3qjhqjvX+Oybg59eHn6UUSbee/KOO05yHbNU0CjSj13+hBcAZEkK5JB7gy2Jqcs0lTSeObfCe
VwXZWvkwd0dC1UC6Awa3foojmBf/vAID3n31dB2Gb8g8Lbxl264q941WEnDxWcs4NuMqfuRdfAbs
wDbEQaZc5dV2AQ4l3J3iSoRdCRBLeHEwm3k/p4l5tqCFUnIYUBSpfnPkMv0m0Appji0GnkGJqphT
Vj13h1COvaINvt0nJN0tguqIbS3PIAGNfaF+z7ZzLCP6rDFtXgREMbOWnmppm+ATykp2harxpX5Y
QEVqnFxQ9CCK1TLz6a2/EEqa8+u4dYcreB0kWm+MLF7SoVaJV3wKvF6Unu1wPowRlCbcPbb6ddlR
XGlP8zDxvMzhRXg/gj2QkjfJe0vkwHitldD/QTb6L3N/rI4Y147BzdEhkmB34/BgqzJkJBz8KwrU
snEX2gWX5rng5T4dXPRtlXA28YOQm2pWbv9gNQza8B6MlTqZ7AygNCUKDsEEwnlxvULO1vtO5T1u
hYbjPiA2CRwQmPCWdGR2qPl4MJCtBg+CC7tMJ8W0Y6Ywh/URgxL0PuEEQh1+OSEX0/PfTCadoxNn
rcFjz188NT7/MUYbFNY1XnIJMtnrax9Lw5PN1Pzga1xP83lR4Xagh1CMdvzG4e431PR1ckA36OOK
KxI0xEuXRO1Jys+zq+dyowlpQiEKglIWsjBwFUMYNtG0edXQCkDIVXKiGTk3/RqzI4/+pb40LCxk
UTbu27wFH437PG+HiV7jHQjniao/IuHK9cItxvOsG+VdPZhKha0gxTy8Bv0eY5TZK0hRjV/oWBsm
Ia7UJcbXn7p02AC13Ga97MxJOHPi7gBCH3sAEoD8+3LlbvoBREuR755DqHd1FRFYapyLnk0K9FFj
i4fuTDeJrWvcnNf8WI61WxT4dyC765V9VswZMaGvfo5VbmCJY2s8cqVNu+0f0P/YBG0XZjL9coZT
eM9IxaymEbGNJkh1/YoUN2Otp+shzpxhwxjDN/P2y2sliJSRpuCubkRdvi7Rs+/Vx4CokULRrGrq
RijUljW5cbZ3Jn5BErKCa6WJyr7lktFVPmyWOKvIpas2BJMX70ev4FT5w4E9QEZIv/fqneHVyA70
7UJE2wiEvBNkmqODlrjjMlOWRvgp4qb5lf/DlSR+hyi1GQfhGzXke2gZXg5os6BsVBxGbCTgOTnx
89NIo/gWSIEDNVah0jWuHPf6wUd3F/pt1pyEPor5UDCEj33faCQzptZx/IeG2pr56JDOroUCHXV6
O99GqSWcp6zduu8IPrAc1dNyLtme7GIhlBJ4uEqZCp1YiIlGMzJmMecAD8evhJ0W4VvvoMqz2o/L
8bFN+63D1UFpBpGXUEye0cdgU79viP7kmEi4MoWZFxDhfVRKfkDX5CbOVDntO+6bczcOOFveVg6A
EChdiYOXqoPrE7dFgADN6Y7eMMRwwgxIGhb1U310lvg4sZWNIAOUaPaQhb2eKU0o78Q6mYoXAfSu
Fp66YOxSYBMPAHMgGHM7q/b7D258aTxeZRRJEs4kcsPLkC+SEVDTC678lA9NSo7PMpYLyaa+phYW
t7iXOND0PpUQ7uni3gNAcZeJ+Dvb/1f4ufVaWqL20AEJzRPwUdkRJCI1JZwgMaF5E8NWXxZhn2ya
yxfybaLebRWGZisRb2U6Ddsmu3TjAZf+6d9Sg0FhEAjIrtuF/2hCoB4imIruM/b2hvbvpPZrXhIq
6MGQUo48VQPrKVpBBnTtoPq65/uudfsVd3KMugfFfe8MsfdmLMs69+1sHoqlx7RjLsxI09OuLS/A
tvS4qBBaa+8lVLlgyUQHtOgcCOsZZLWCw0mzJzSn/aA8vqZVdfx7XXghUJeDYYKejoIOepS/5V+q
uuBMWU9hYwEZi09h/wx7L8jDyHoGFFO1hxgPV1gPj4bGLwn8Slw0l/ynhYi+1YOGHh7J73Md3A1w
eBfhPANgjXk7E0DD6aEr/uG6PXf5/u2uAtLtVvNwTSHvEfmVdln6W1BLShf/a+MTLnlPLr9ISGpH
SnSvJ/NP72+UABp0gApipHR8ZUwPcq813AKiMRPyUh47OG7v5AgFGptvlFMqmZQEp7xM7tlsRFZa
FAY0hZzoDVdEtIhtrT3H3258FJ3o5EimVJ1gSyGfK2JVlADXENFN5nGfyJJ97jr8GbxCGv5iCKYx
zSin/4wTjlqQtnK51sSvcHFE5oAv2jgvJddxST6FegJ3mucr2yuNH8Cq+XHl95lo/R2GPz6cSg5d
X5mM4xX6XeEuhJ3iGp1OObn802YaO3HSsfrteMnBclZAOXVrkdUd9Usb1PvVkKyH3eOKROcysCV8
jG2+3x3qOLgyzibFRM0eiPySwnMnucv66rMfZ9FDdw6TDDGmmo+xIgRdhJXHkL1Mj3a3LHNngzDp
NRRGAvKejFFez8IMGM2xgF61SYgCkrFg3CGYTsC/8PRdzqHcm2PrcjtGvzetRJpPmS5C1CtJtlpY
+PDMHFRiojqTV4t+kzwJM6edT4sqUO/JkltKHA5oaBG+5jbZRcqlBoYKQDYBW878a5J3LozS8gfR
g8PbTkmOMuoJ1JoEizxK8I/j2Rx7mBqVvno8wwe2vgHv+A7PDNifzMRUqKy7pk4N6HeEE7aKtkI1
xWE/I/rqnm9gfMxXnKRf750XJVPNlI6Wn5itCv6Mrh0mBHxElvCQaCTlPu3SUSc7LqGUD5/b9vNQ
O9u8P1jlpTvV/XzbwDpvDEdzzYsH/nM5gruWyx+7cGns6Jev4ZRgg1SH2VabCTRbtqOSxbi4QYnB
eHj45+u0innB+ojZFnV4FcHD/XF3MP0SAu4z/W+67XJLlz8ve8AefssgYzcc/Rlh4yiqU9hu/3Iw
ekYJ3nnwm9WqvGAiK07OsMnzMnWFqP4WPB8v9UgiW4H5thIwGq4doBeulPUEhaYQkU1MJCjwYrgc
YiT9A0A1x5rXeX8AJry2OwiXjIXsrcr+ELpk9JYm7D+/OWQXKCzRyvJQjgf7frLskdwRMii4pXrH
VIcDXYz3KyAL/KBki6Zs6MAE7Xd/5mQOUASEWUYA6z1pX0F9IrDXC4MT/RqiBxUKm1wzp10XfSBA
VLcWmtLE6HPGYNR0BdBlJ2btrxKAkWWYwEkW1OembV9dG8xo/M+6n5YPqWnAg+8UNQfnfTjJDUJu
MYTMkTc1DTJxImXac9s910TQlHdod5hM178PhQV/Qwh2ed+UClk5LG/OPaNoaVjJKUrantvXuw/+
NfxHOj183EglDn98oesGnaOJO8K7upnTlDbuuqBd7SVu7shm3HhwgoUWgkoqGJ/x0PLPQ8clwmvK
iDMnDLfbqqehDetahpe+Gk/N8QWASZ2AWwtdLopZt2YfGnGxPfXqTaTcD3++BUP0WeptHQf9IWSd
Cxb5z9G59oFTM8/EMglS70U791bQgxtRzyQ/DeW9O8WKOekOLQA58tdB7oor/osp4Nsrm0l8nH2p
hE87qto4YdV5azJ+oMJFp6RN3cQ0b9yfvc/HrV8VBn8GbSa44mMf3LJft9I2bSagVF08Dx97DS7S
wc6ec0AcMyZkDWEvTTvUX4ulxHeETNwQc95NEPuwCuVAvYTHFxw5Xe9/ihZRCpTcwPyVG7Y58oRv
qxXLsJvsVIxwMtrTB8M9QD/mgkbgDGBh0bCw+WD5MdgXaaCm67q2W1qZgc/WZ7eJT5k3HppQ8NFI
QVfqlHWLuuC+1lidb5FDfFYr+YKUOnlcegZYlJ1r9t9mDlG3JD0ASYyFcGvD3BE/j/baSy3h0Dpa
jw3EbluaQlQbZ+xxfOOKpJdycPBpzfnOFh/xRKks9U9zYE3GnbOV1bapaYpVOea4Q6nHPS3Qlkz5
QqEF7BSAz62cgcWfwvmp80floj2fXOfMFqSI3iitXy55SWejXzxTHkl06kEgIeiZPoQpyE4Yp+1s
X3Wm8hPua4R68eFhAvDgUitmx/LVRUdMQZ2B0A2NhcQvBh7ZTziYCGJO7P7pJJfcxfsUZZIoMiyX
RAwDTksIU6SP9S6coDWECFZYh6A40NscE4uje+fe58yf63YnGv6Zx1jRJYie5Fep5ec3zzX1E4np
kBEcl5Xt5wWVxXycFE5sxFLZbONJ3ayLfQ/NRW+Gh/0Es4lguJR2YFCOVCYvodgKqXflOG6DSl6H
XuXwd9GVRxB/SEwNJatF0ZgDNkRW6OxLj6sk2uQN+TGiNwOcHx7lKeStOt5HhCyksbHjZ3iFfw+9
N58zqRUVDTn0wTBacRv33RBFJrAqliXmHjDqDNm9U94qLr7WIy9ftrKdjQEI6Lk0i7guKAOpuchJ
vBmdjI39R3uWR58kZobmwZyZCZOMLrXc6zmxmpctrOY/Bx344lQ3wOSsOIRaJu2o7/s8ZzW0MH8G
98ISEwBmESuZzy41d7S1eyN3q5d2t7cZTziEX9Z36Va/i1CQtaRJFNkart/RAQsyIWXRJRZ2U1wN
6f2tSnmIfSi/ACjwPHivIOMwfauB1USQOQ7fBvqlQPF9Mpkkmkbp9zCIVbugxr+qHhmM30ppEiNc
P8Av8M5S2URVNF1OJzVA11tb4aOnhTfQ8AehTS+QXHHm7hTu37LrpVHsZ/6ppjfrOjsofTw7sMWS
1qoHS9Lqmk8P+FiiG2Dlyf80QPxdL9UW6r4Zb5aarcdBEmXrBPHZKf/soXj0UBXc6+m3T47Htpn9
4avqpK/SMQWsmdbHfZqZeIsBCt4ez35SItLohggQIam/xVVWLBbNWecQn+OB2uBe5f5SqunioSrY
XzwsBJSud7aj33douypisPRapPXjyFP/7myac52vzjYqI0yPGsvoF8+w/dRx90Dc+5GhV1Rec8jC
DtCcS2lixrt5Bx3O45xOtX2WFZovSvGRyvAnR/9f5Ji9WQMlRPeLhtWjhviNoAqt/+z84Yl1DukV
7iuZmcxe+pdRpIJC7U7+XHwLrnLA4s7kv/yF8Y9+IrW1ksEPTMVPi1BZSsm+1jvfdL0y/y0c5dju
Le7rFEgBF0Pca+KVmKv/iCJkxpQsDkl08iLXq5xRsD48swb9E5ugovazV90VYYEJa3KxepekYx8l
VAFLT+2QF2igwPHh6DUruDuFwaFSPMpxZ27MpVQnwNLG7r4cy/ISDZQyEt6uUivXt5yXTmdYw2qr
g2Y/LHZw4ytpt26eAVd5/FqVIaIQj814VXCHlkp6kEf3HOkNU72n/iPxlBAYmrYK2NKRC3A8Nd08
9o6TN1ptLjgXG0fXgwSBR4H1yUsonFxPNQms6nV5KFf3Al6hr8zMTKQK09UiLFd1aDU2dk/u41Za
PPbW8zmiAwnGcFlQPTMWbAQUcglI/FAwvOPtlo2Ye2DAfSu0u8qjHnS9KvxqBoXRMTvmYM//Gx7R
bmObtxIJVtGZqXgdSxXzIOfegIZf7ooei/Ysn+/W9sNtkFRHbJzKgYZwfOVw5SKyjWyx+3nYEXCW
OOURPx7oZLyHV3ar266tIkPv58ATh7z2b4f+Un2oFC6FjAbif+PJxnMVEL/Oa0aISSK4MiFSSSpN
z8m0kLt5POQX8lXXD+0oU+kiDA1T0nZLmtECBCZ3TZQ5FZLe6zbP9lQHCKrPyGot9Q1JbfCBlfTe
cOqvU9x8fiMjZKnTJvT6gst6LoC1bXJhgEIdfKEqEw6hyEOME8/PGcPYVrTsivY5rb9kb4Uag8kP
aEilnfkPu60Kwq/rSVPLpL7tpbh+5zPp8lAyKHeRZjcJLT3cUpc7NHTqXjsdFg9qCQx+W8jV2iPs
lh8EIChCTz+lpjJlwU271qzSW06iZU1w/vlsPzIUukSVEGXQTPcxujDW3fNijm1KOvSHaIbkGlJd
itzFTguN0TDVneVGrTB46raw7NvWoaK34hOTVCMjowjFkAQBanE/AEM2qhPKBEtytGbESsgb2ouk
pGwsYlAJWxYlr75jYpQKwclh+pVq+Cc6HQq0zohrhKBqmTRbcUYe+pAn0ewc2uFpTDfWN845HgHW
qesDFZ1FM0l32zb6bI6p3O5nWr7isIbajMRKZCXs/yKgKdg6vEH2ZYO7KdvLwy3ZkB6muWjmiwgx
hwputOBXxKQeayc+07FBdOu4UMpajMuhL8eR7HIi0FElJgl993oUOuc2F9LmiclVqfyBGiqNPzOK
o0hELtIffvsLI8oCr/xr3VE/wWJ071O0OqoUu3Lo8o+odbkoJPMUIe0/weaYSuFtsb9kfE95LGQW
I+z6dqMwX10DtW96d/F3bGSfu0/FGFGwKi7NFDzj29AXbhO21RerTHSlDoJAwUpLvDUrfhkr91OZ
AxtZTcJgQ5N8c+TB/xCGmw+MTZJcL0Y/Bekik+hUKQMhrYecBEbKoe2SlEQBXmjj05BesOg5o4bd
pZ6iWza7Saiyj6YAtqBuy41conialbjz4flx3kSvxNSLdzq7/Mo8mP4FV6yp/6AdphKWmQRJce2x
A3F3on0Zu1q+8dMtVqX+ejLV0u8hp1atgTQkz36+Fc1EyBzhYKVPK3zO5AQD3A2TlGOlsTS7joo4
lIZILUXJP/kOU2xwplWpMXj/DtfHofDvUHRRIsW7MTo4uv3t8yblfShOLJ4kys5yDx+D5krJc1Qr
ijdSARuxCtur3dBsGAAw+saPBmTvO17hlZ9PziZ8t496WuGW/N+t6+76tJtyTE7BPm50/Yl8XTS9
wqTbORCXcONr6AkIwoVdyUrYfu1kmrrMSmgXMW91dl6QFpIaIKcyj/vFEyNm9Z/e3xM1JGQZgvOO
i95x9xG3Pv6kHJM7/DlpoH1cT+yxRK8vO5+3cIsFbN9+PwC+n3JodHfkxHK2XE24LmjJJma7k0L1
/stXI+Yxx/GYArZ5Ux72cmXVy+MNS2pVF1j6vyZ8WVYdI76043+OdWyWIoK20b5yuM5cAAzUah1e
ybXZAVBEP++813Hq87DNY6UfX8fNjYErFmQZNeztC601Vmu6WFZuBbTaqmw/p3Nyb4JB1JUXSu1q
eWdP+bzbfsCJMzGURejvm/qyjX1paQAEouNs6gqDWOj8L8y2MSPDoQ/pDsR2BI0iY/btGSHDQoFU
h3JSqpoS2M7T4gZ9gtcVAARed2cvXUUM6cmAwnZwa8cuJXFX6ZdvSwrcIdjRbGvXEsSp5a65zCNp
nYDJClrxoJw5UOfYhwRmp4OJBbJ0VnbU/nu0v4qEiuuRa+xnDPRCu7H9JksY5d737jnFG1MqBjSI
xEaAbO6omPiWLMebSX+8demjkt47qjjRVDO0xQC+MqI8ghS95cP8qFPeRUtL0WbQngkkeQWJsOfz
8c8+hYczuS6ktHzlT7sfO27zrA6LuF7wOR/M/7p25DG2eSC5Idh6TnwD8EvOxC4bMyxySDD/30js
HsZtnsw/UFnC7kOVaATQBJEHzz2iBYj5Co7A1+xWRlQZcJeHCJKDYNZHjoBEd5kYFXEwbBEJMV+1
xEhBLGIRS4OBbD6LhZNNQ3hHHhPl4QXfCs61eBW3vtyVP/ixQoZI1mRDq/MyKZjZxH2afoix8zcb
UyzNC1w26iKKQh+rycHp6xEr7wEfPNr2XQdo906sSP1zJlChQASG5gzty8nslnPGmGBhmfjv/dFL
+zx3+PpNLJkjFMn6KbVl/VPBmYLa3IglEZTjsg7Rj8PYJpVbNw+1SDIXJ/6mA7VQHAKdE2T7ci1n
UWGDk75nFSZMft+NfvHLOr27vFrthWtDMhi8BM/SqxfcVmBY0swWqZhN31dSgUflLF2grkmubojc
rqqXvY7QKuW7OYBm8Jku3jsJgNQNYRcH17wehcDPWqx0YABgtQceDMx8nY2dyuEcdupLMvdjx+6t
NsiPG7sFFNGFjOJ0Ac8fLsjEq5hxZ//ofXvi18OjQ9GZT8fyM8vfUTRMx0yPMUbh8LQAFubJx1f9
niq6fpMRL5wSNB6I2bJtWfDOSeRSmCV0JB2v6D4Y873uGB8xyWr+dPz4gOsoNBiqYyErznjqsPer
99v0pkXbnANWulbPbAwi8k/pFZSWnB6DY1d518kJjKV4MBcF2XpheVymPdTEjUDiTbfExhr+6mvu
yUk8+JZkOERPtnYAAVZ7XpHiKr1+o+Xhp+Lc8O1vkgqgy746xYSZl92yAxPvqWp5oRrEuQjFUFcL
XcwimrU1YAV5T2xQC2KmcjAoTaRZgtLbxK+cntkoqHLIJUPzgn9KdbBAWHGclYfxBltUKWyvLihk
veBTjKnpFYXFlEAsHIgpPIMlbvNO3G6VZHtL5/3+1v/qdvKldOUiKUwMhu+ZKBCSIuTjDS/pDCuh
wk5rAlhWVHWNk14cds3WeFIox9L4hEFEL7W9J2zoGaR5AvZOxjCOBcgFqhLvAW62jTBtBb1RsO2N
07z08aOuuTLDOCs/xKGNvaC53VQdzgO++N/t5o+pc5RnZDsqgY8jAdhQMDLWsRoS7FGMt24fLLnP
bbTo58a9w7FeofIhq+K6kLO5XUtk/Utj6dKYM5CHL6tqnZtf1HaEruu+HD++SHkak0DT7VemRkr3
1ggsg/ro5J4yHzzSyTk3DEYLrt6tC8+zOnFv2+fmm4yHXPioyJA+bTQPJAFauCAGgH23YmgZtVIz
P9YvAT1P518lk+uAL3Rb1Z6fzU80tLWWIjjFRAKCwsA1qA1IMVReWmRouq8efhfNcC4GvwX11kkD
X8ztSeQJMXxDFgpT16xQrmpGDKyMVGUi0Eo8CrxaCgdNz5N6vGOOiRx/PVpWbDV6BPaO2eP/FN86
OssZTWcQmQ1PqqU2yUXFLFVwQ3UxokYrnN3qAjQwiN/kektpVh2SXC6cuUhhzxPjXMRPfcMJiOxP
8eoJgZUNEmUFkyJb0U14ADe0AxJK/UQOli6UWJ7b02pZFZPv6T6fwjE+sM+HzXIXx6ttmfQHy2dD
G+xLTDsrHJNT+wEXC+XezBrkrRHQkVj/5lWMeonggiiwBlmdgAg2Xx+BkSM0oaSGhcgzcG538DOX
poMmvFHRYYB92/yxO051/PoksQ0qbHtcG6nYeFw1REGvJ+nzIzyGAuKpzyRgAK1jiz9jOmKzo+3N
gtQqaJnIVCiiRvr1e/rsJ10qB8fyT1nE3ZUrGPpX4lUlFB3GngPwhp+xQYb/gAPxU8Qp1LzFe1dw
dP8Z+RKccNTsvPirYI/UhG3ia2W0pKGLJwQTpxRI1PRnOmW/OnBRdUFlMEWUUb34IHsq2r8jMfJb
xFcWCOagdXD7CrzqInthQzQHUrpwyWljbTmduSxuJvc86PQlxmnGy+gtzQuTcpRqUI0kP7K5+Bsr
Zp2Rf/YHPZoEGftjo6UBLLcEVOVN+xm+4lio7lzOXWBUW2T/hgj5TID9YA3gtEseOZdduVzD9AMH
2ua8c5QKQ18JXik6Jtbk4RvbovFgl2a9o4Zxujyfz4i5zxVFfcDmzEpInwidQEokrS7csi1HQHxk
8kk+MPcNRW7N4PSG6ZcCyeL96xX5np1VXRh8xsk3txNp61x9hZbjPViUDHx9qKO0ImivUIgtvXiN
AtDJBSKMWSW8Bp/414ICzmYlLYhXyuAaem3mke2SLpTjF8YarogXAuYoMmnQCNSXQulUc77iCtTR
ZbnMC139iNJ0RxBYHTPRxmLXpeJiy2TzNrmcDfCisH74+jrr4AVpzYWuiZ5fHPgMIQ4/+UHPEhQa
MIVpQDiSSvs2AXblYlsJeihSw++XS1BCILhsdrM9wd5LckLfh9l+M2nO6FG0It8XQTGlZh6tgZ/Q
5eRsPqt+bcXt55CamvfWAygnzz1pAK63wcBt1YgnH6WI4qkXyH9e+c2Q/wAuai94aaQ6HZOwBr9D
XhafkaxY35qLAL5KxUEWLfr/3qBEMcS/cJI7IyZPRtQa68SANcNy4D3xMdynXEZZYkjZZGj/7G6k
5UIOdbcMFKa6lyUfkmvVF+q4U27sM+F50zLhwuMcjP1TUOSDaZpIUFdi1LgJRvGO8xVdV/DJErH2
Xd5W2rRtWbqXvr3SceHnrwp7prqHnE6Ecuh/jxjs0LgqFw+69FVasPfffbUDBopCkw8+uTQUsxVC
QdrFiEcmLHrmjngFuQFRvZwKhl8whsBLLxdKul3Pu6DLocUOsTm+iL1ZyiXk58Zait7l0MY7orrz
3Wz+YQ8trRnVBDHgex5WXghJdsREfQ8BS4oQrCA06Bo0nAYHnbmCfHDa+W2qOJcyC7OdenEB6/Rb
LMSNirMdDG7wLp3fsSrTdIjfMk2ndTKenF3hnzzAeynoIsOWPYh0KZzfFJFhyZi+nu06+eOPXWfl
y/xpqt3ZCJQiiXZKwbrgBgLBm50bl1Wg6t5rIpwi34NVFy6ryJqUpzThr9mubaXcFgHE3oTBz2kA
/ZLPOYJlsk4drbTRhqhStKU0FfphbOluKezjzpHaAwWUNEBWKK8G2xncGQqTfMcnYwkhS65pD252
QXw60bdxzfeJEEFKtEnGPkQNigwa+CKdsrXn3W2wqP6GJFzOF7e/zwBPwp5XkbrruPOEYKvRaOgE
iBMerLFw6srfbK2fYxGYLFzO2z7x3uHZJIFs0u5l8XVT0W0PlPXKrRksKFxCRyyMSNHI52xLyW2L
njfn8ZOGzvVyXe6GlfsPT3oNojir9JehKYzGrk2Y39XJxrFY6BHNlsz4Wzbp4E2vqadyz/QPAevu
ODMi4/A2Q6ZlM3Uh8s2wwaL3yXUSl8Qwc4fqKlGs3eX+ZSKh4FTLZjEFgttvO8UJ4EaJHEpz/M1E
3c1wIqMVK+VhnOE5eqobneEBGvcLwIHdJ103FHALsKQQEl0lkXq2Vd/QFBnAW1R7uNEie8zH9+q1
PRm7hWtUVX+BBTwktMQtuA/ccSKwXPIODgs5vUH621CHesiPbfCUCqXfsqdrPQw1rBh9hZR+cT9X
1DKgff2+WjVgUh1x2LhgO77fr0qmo/NVHoX/wvnO7HMhlaxIrQU/dRQDZkw1dsWzdoRIENPz7YqG
NwLVctxTDlFJaIJfpAwdyZnv8lgv2F82cbGaDAS8lNUplTgRL7mz1U7Kx4RSfPxMkkA7V8eoYjZ8
GNLdg8THLdTEmenU58PU5/10HUU+gfjj3YlP7k7rMAaUBtiBIK8XvySLw/tdl4zhzWATvKj4XVCM
C5zoo9QmKkD+MvRA5EhtLSMT+6T1P+CNA5KL3KTLuqYW2BEWKWoMWsSquga5HxIakPxWbz07R3VR
AC0S2VJv+5dZKXG6l3+r1+0q/PUaQTgws1iioLpLjUEdy8mLYcaPJFLEAmGRoBv2g/czVkgcmwIp
hCuFza8NpKj95ntG93tR6W/cUrGAjWdniHUdtCIvomVuEsRE0ZAfgMcwgqbDQqgJpR8bL18by80c
qf4pSET7V/gKKG6tJu3Pp8MjeQKhqcfCNtWkXW7xjV6yd1e1mCnDYdN7iv4D9k2KHooWFRm8wfoA
cgs1Qqjby3ddSUcxIRsFx2nGKzdYg2BDFNrV3DNgXJZIZ/XfbSdwZSTIv4kTP3qWdZa78K8qrgNs
tllay2SutQO/l4Q2zFMQVq0qcPuksnDPY5IcFC/xQtHmKutuuHniz28HdbO3DfCYmB/uc0n5ltBz
s0xBIWNfU79LXbyIoaNDVDNHy7NBLHVdUzgAqPrlImM7LrzLNq4KBdcwrlEBL7MjSY74pExyYyWJ
RnjeoNVa9zz4F38K4glc8H77z3rneN7mV5ljIGy3BVMKUbIiSuQgT0YkFUnL7kst/K/ZOZfYv2Rq
bcZv3QAlcbxKQvB4+gB0v6ZF7Q41+DT0XMCAK1EdLgMnnAxd9zk4M1BmdERKLMJv4wZDDL/QK9RW
Gg/2hJaZCDV2OD3l7pp/aXWeYK5H/lGGXYMSTvQoFsQfqnBHlybxBURn4dKGHs87vjfiE+JWDMzL
/7zdCvgTkr4c+RJUVYgB94cgNB9ESlfuk3XssCGPDsqzOvTu3/0w00eDQWZ/T3w2KpCJN/dFcRlc
bXpsoNUpbN69v7583FKIa+f5ipKxItorfQjr6kqTkFdJFH8FibmgmPWXwClB2sVyPh3PmmKnPzSa
kB69BLkpqmyKYmr4hDstfLVE4rWrljjBg6YimBRcTg/xM0G+Az1IVBYKukZRToPsJMUu79dcNohO
YtQugSjVVZdpbteyps03a7Mv8gyvHbDjMfysKWLvZto7AIYzcCzP/fLgN5y/kFg7A1lWkF4FIe9n
U16b4N5AJtzyblrlfO6NqCmVcDjTas07/vvXIi29G3tL65De1gSPeJbWleB2CTqlcYlRONwoQw5P
7a19h31/fuEvoeQx47SIOEDPoHg+Rklf1YCST+/AHT+Kxjdg5+UeEYQAcCFs93hEdYKBpliYO1TV
B2xREFBWoo3PNUCKLcuCknO12ldRBPu0VEoYyTjXABKgMwhLPso0WONcVaRXC9pwSA+fXAR7V9VK
cm+bB/gUq003Iqv6SO5/0XsfLZXtlEzwIqcFpbAZtYbOW2xD4q5U++GZrls75+FcGJ6e6p0dURYD
3fFf6UOIeVXs5/68kY7dp7GjKBevS9uBENxPF+buzaC1JZ5CEzHiSLHC4wuNlLzGL3DsDsNAegs4
592ccV5V7CF2+4/bK/lG3P8qwgQxqgXQU2OVY6f8bY7T4L3KbW30b7gIG2tXrDwtY0AHNHpMCeoc
9RPCmBBX781NmOCLtC4PwKFXDB6Aj2ohTTKy/OW7O0LaZ3sAQCI8iE2koq4J/y52QPd7caG++fqS
3TG7NHgYN/m0yF+EwKbpYN+U4Cv7kUPsR6tUg4Kadptd/On5Y+D6fzyEREo9969JqfYVCTcCSxaq
+gr5BIGOeeyzQJvNWBUmxJxKeJ24RjqxUx4QmGhVoF9a5d7+OTBH5crBXF+p6Qncf6E4hXqkLwXQ
A7uMl0EgFRJVT8vmx4K1QdKnwgqywRbmb9UkHfKeRM9GI1BMhUOe9+/WmbpjoJlOV2dUzig7VgPI
LLfP+OnCedDicoFdouOjEMF3+8Du1Mbu9Loa31puUS10Dd7r7xxePeL+6g5pAJquTAJQO3kLT6ZX
+koijrwbgDiuCP1QgF3IbVJJkDGxTuQ3nAMESwGBc/AyDq0WjoFxteKwBnYXJth7D4lV+AASgqaX
2A4AzZVXIsefWGGvMH9p5cGeMfCiFlG3mtxfDDuownbZYef+AmK8a/GyAG6P6lldduCWWUQm1+T+
H100XPrtRBmOAsQq6owNw8piAG2IJu1d5I4vRm6vKJt66OrHPwxBC1F2uI6X0QbzLAvQU83or4c7
RAxDT4DQbifCxR5EbVBTYjU1u/ETEz1nyqsvDNV40LuWBh6qhS8pKTJiFPqgsoHb9rM7SPqKmn6R
QzUhNJsQssV51CcVyKewZpvEN1FT5Pz5uhAoXRetWPC0B6IgdfoBEKSxvp0trivlJfE7EqBNfIhz
Cvd7Ei2PLYve0Kp7xg6umQxSG9qwYNHCjcdEviKzifGV1bpGrSDtKqarT0oiA1FbxP0lTSV8GhRP
mir/pKEMBaamguvoLXCGatZahivhOfSyRc51A9Db3e381Od6YUFGCmGYaKH/HcvXpV+TbKcjN2Pe
ofCvOirhTA3g2VvqXOWggaPRf7RNyN3svtVuPquH8y0mUE1SvPI7X91QqSKy331H+fydwcpP3HAo
lGbrTFOrD9wAN8trv21WQwNg7736aZ5eK8aJHMuftDOXjq1H76sbRYfZkS7ItxWhP69gUYD/7gU0
n/02YPXivf4toDiRk1FK+4AyOyoIj+S66yYKncWwYPf8F84HAms4sYQZ/adqv92TPhjpnWKDrQH2
ofeba9R14x6g9vvN6j6IK9J+czU9zNLjOWjFwFCVzwXHBdp+l/iSX02YmAY1+q0kHJy5TiGaLyl6
juAmVM7XVepITnAS0jRJ8ADSZ7FHBVbcar+uKb5hNtMXKv+/2yzPzf+eRf6Hx8YpfZXZCxKuZVo9
TNqElzTJUQWrI0aFi+FHUV0vxmIoVKu8oXnuTM72BM1ZuUzYbSBTxcUYedPu26vOpUOk9VulSOIn
gOZDJ3nF4VuJRpt2x1MWr9KnNZTCtvCI4NW1q+xsv0e4+Kr7iOW1RmLNG9tOPoYsCsDwn+o6bT2J
hdDAFA0BF+msb+noviNUgCMpDPlHPMKqkGjGs4JJzkokna7nIvb5uExySkEAK+aV3e0p4gI+AxvN
lrsqXvoUOSVo1QQ+Ij5+JIwa+s9T3HEQA0OQ3KbniwdSALaWGz3sz3llTA9b8aasKGzM33Uk9Oki
wJcTqvB7DHMM5lXRGfbsLritwge4L4YMAuQhKl9pK9D38sm4fN/j2+clC+DQywzSoLIgiJJMKJLZ
vyXMOqlOIjDOgapjf/LrGpy2kclHbD1gRZmUI0tu9tLPNbb2xy/RaRQWr2ESJ27JPkwhecR4Pzaq
jxOj6vSZ7eaF/a2SKuPwQ5AGOurR0bmrSID0Ma+zXGl78ZCSpIv4jA37uLIvVxXSCvSb6FFcbjd2
GLLa4+9BEu+lVq04N3n9MgescC5Zr8x2mrTXwXkNNamZNPAmHImVEgjbUoI8gnQEiQjza8PkF4MD
23GAG6PR2n4ZLj0ryHMmtaiyCBQJuTwrn7S4VCcCXxUh/i/TmaXWZKRtgb1L+5NlwRydcq2IUld6
++0ncfLJGrZ+tdrPRPSW5p1uGv+LIRgVABarWGNv04nBmpG1gkCef5o8/pD4QFfBK+Viaoz1BROn
0Qe/Ag2KDNOKj/RSze1WQxUAGNNUmJpRPhYGd6Ga7MwlI8SlpHY4xbvNncfW5uoxVX1LfyRmJ0TS
sGq5mvadlQoCq7r6F4GZIM6Lvg0YiBlfocqEFc4Pt4ijAjbqMOTjwc3i7rADL04cDuw8OSXnMXR7
W3BVGsDFk3k9s1C5niXmywTacmshHQrFAFu0z2UToFJeNS4/Wvo26v/kF7cNx5+6NrFnSfKhjjRO
/s4o0Xk5TAbNOkbntqBG1mc3ocEs0znp6PoqSqGjXPEjvrreyWwEp0g+NLDhIhF1pfZDnlXDcnYs
NmUEZv84ay49RXotT0TF3Q0Dj6XMEP6GLt7aq3of65IFVNLWsZwREAlX8MAc0jMA58q32www0TLO
QrDVB7BwdArOLraxn2v/se6jyvbcnE4/eSLNuDli/uFnjbjlZQFqiI3W+Jg1urUPgNDIiflzpCxJ
/Xrw8OKyTkB1SXYLDU8FaVxOfaj84/+q8fWcA71UVIjq42a1F3NyPn2E6BauHQtQ/+9Hn36ZROCW
eiySVV1nJnAC5LIOLFZVtsUjNifZjj4XIv08raJSvkC0CfW1zJT8PdvzTkvzwo7kDoU95CZ1vnF+
GfPpQx7JefXGevMna1vwVg6I1x1SX092yHpXJLOvqPdYpYkM8jdYN4yUPq2yWjANdzrIHY9mesP4
jsuOysyXjl0huyH15S58jXVeoF8hBbwrLu+yD29bu5QZDRisX0e5IkSTd0fFtKTNVoly3plY4JtD
KiFsQHMW7dHUXNqlviIdaXZ/Z3MoyuwDBILfXLA9a3JeGpoVAgwjNNWrlCuYzYwWCWOqKwWf5Etx
oV3U2Osij6C55Ht07YVayp+A1x4ZUopeHo+bhwLY3Hxhh2YSbhqEPVGu6ngQ3cprMy4JhqwrPxYP
jl7dzD0+xuZoERzrhUeTcZ0k6qvRmQluLoSQnqeSMTgZGcXWOnxWozEMVA1oxcYBnhKBS4eIr3Cm
mEdthAggd/sGkCmSHgc8AO3dF22c0ACKu2ufDLcrZJ+PDiXKyBOIe/dfXAJcJB9abp8qMQxQoVJB
Vj+k+jXmkzeXifSS19MbculUFT0nYid6YqF1us0TiYNeLBbTo9z9Ekjuf2QXQl+IzeVItmnH5NIj
ZONSno0KZFw2BdLiaXMcbNm86ZS/w2Zi03YEac8B8DaKVhZdzwBJeJqLIzF69nthzKE5U2ut4hzS
6M9ie7sh14SG1PbP7tzfmaOPQH1Bhh+UoVXRGD4jcsQ5Ki7eS5T2J55aj6ZB+6pgFzRc8tNAd8gl
eo77jgveROUHoyAnmgjdZEihPg4S2OMm0X8fhNRqdSVrYl1Xu6D1fyvq8Az+xrmhZ2lbkq8rz7LQ
kNeTUB/gvkee3YrgSFAGRDYcTJ+0/NRiwT5YQeRUMn7MNwavwlVsjRntcB6C0xD1Klaq4hilp5ji
2kmPAz5tsl5IEvaKokvRYn4OZ15zrF4LTx6Mbm7T14s1BMB47vyDR4MLutfgczxylT10xGasH0Tz
G8s1pRKFh13gM/J0OC9qJkGvaUopfITzXgIWsQxxvddpMjgpObWKuyMivxMNWj1scUInCmoCinVZ
0GU+984rxk8Dfe5mHcQBGH18q0jP3l2OU413t29+MCLGtsRrRpY4ZJu07ZjEexYiYo4JLJwtqcfN
9TufhS622z4XVIn94x4thjgXOV8gUDfZyut0W3zL5mZfIf6Cs2Tvtf0u4yaJUOPAkHit1qXj0mul
e5G/m0DopXlVfE6FxvaCcXcVZuY9shbfYJuIIBMJvXsgIgjavYaGAAjIbA3ceHn2o2SetHDXOyS0
rW7CRN0RauqRB5Ua/dwHQ3cjuyenhcBasYsEVw3S4VOd5kxQ5IHPtTwSxEuIJmcAGM8Vmir2q5Au
iYNShSyh4PsqdEiKkOI4gtiAcmRrOXhNqqfuxmmdMg0DG40ElWlP015fodcbXZf7XpouZyHo2Du9
pCRj2gG+LaszeowGzVeqYh4uDsL4ovrX5xgmoVqbuLjXgzm49f0s2bCHCf43fziNr4QbK8f/arSx
kNwf249AmZTgK7HWlB/c
`pragma protect end_protected
