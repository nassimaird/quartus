`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jI5JbuQYxycp9QvFyarS8QpU5KKDe7UmS5DcbBVWB1bhicUPEQqFWAhiS0366LkU
xcZtSVMS0wpVvS6mpMNTPJjBib3UMLVEMF0sZ3uNMt3Nsgg04+OZXFm21rw7lurw
QzYCvvJlG3Vc5R10pGo1uAeVhS0vgOzlKAtc3Be0Qpo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39216)
ebHJAS7qeIbZzNyoJr1CxZPQVJa+X1lwlJVftTVaOlgmquR0N/Di0dns7VSh86bf
kFDkNCm3gfYMqfIXWuBYqvVhVwE9UQByd3iKp+Mat8Kmlgd1U/pE+bDPf8X3s374
CoSbtS1kZHm3q6jsS6wwN/K+pcETXp43fGTle+bpGBbhsSDhV/6+Nsj9B9pT9zqK
UrNxcpx0J/6b20cxHsw6Yw7PbJbKzJc1R/TMONARCc4OoMeguyqvagyXI933Tx6X
nR17nkBOvJFXJVifEPlCHV5GOcFaeiqdcyytLQYG3bI/i6EZJZ7kQBBaQWMPmxcC
df8QwRlHN2Ud0tSv7eCVfZvYTayddJI/JhKqovJZTSvldDsORkHuPnZF7inIGU1b
OlOJ27QVs3AYogIZo1sTcBYy0DL2klMccd8+A3mJzCJXU+rT5JlSIP/dYZqJzTOG
zS4XXN2qWI5MWMyWbLMKo0JjZl2BAS/NmvNYaqmYMz1CqEb/q7Vw1MXjteDtH2ij
/5jP/Dfe/1llfvjMi5v+kboU2fsyrE2L8SuFxOzs7VmXTE9Z3MK4EOfsSR1Z4KuR
QpTHO/56kWRiQ3Tc6NArx/+cDp3LiAn+rsvl5WuAbw+DFwiLgRBWj7hfYlp1/ZOY
4a/WHbBrDEyi1XWegpqMhTVAWrRf4LmihunFy1JvMRpNSxpXVcbnp4H72NoMfth4
CZQIqnKUMxY92HkBTLT2k/RxfL8ZK4hV05mAOCEN+Ua6G9B52f15tp9Ke8l8oCWW
0NU5tluXoIsTY423fBffG7W0y+ogPMWz23y1hms2Mq1gQoA0gcwl6YyA2LBPjGVI
EWkQSlxQEbuC6DiYZG9mqIqGkIPUfk05f1nSr8f6syzhAUAgeOARnIg9poS3kpTn
WHBhzrFY14w1rQpUOIiT3w5MirIK9EHT7fZDGYcmlmHeJVn0tvEzkaLn5lo1ZsjA
diHZ7xu5DHsMnKPFjOsv1xb7E7AOmUNoOcaDui2iDc3oY/tOiVsnGi7dAWW6J5Ou
jxcFX54/PnndwINGld5rrspIWO1aicxCk4eaEbadOEG8M8bHIgPaRglxBtza6QUV
O77dLB3PwrxsnyvwDwFti+avOnczp/JsIS5jWl+oOLb9MPLltoXbbHOxzwtomChc
VjwztAcOQRc3X9/VJSOhNthiCPK/1S0I3pqhX1bXSltQZRdn4pIfAby1nDAk8aSA
SIfJCOVf5l9iqxCZLjMWiiH/VJs7JwsR1bRYiO3YrbUl5VgsAry5ScAkQZra+5QS
d2hxqhetEW9ZzFg6toM7Y19JxJGIH8HCU0fee8+RAcxBAbOCZQqm+RaLDV/bfIYL
VitHBxyQLQ21nqFZMGUx/uQjbPjNVz0Uf63uZG43bxYdf8LTTlrboCD7+i1TQgXg
cGCgGeHH4H5sJOapaBqXipHJOJWwvjHqBgPrpuTPO2EOF/XmeaLBXQC3F7+hGhAT
ieEobtQUN5KQ0hwpWWke0/87h5tI7QmAq6kFkS3BP1/1AUp4A8He2hKT0CT+Ok/p
t32Qjl7dmAx9ovtZ8dvCoxG8jT1A8cMd4XuphLe40W3Vw7Jsf0aAnXDeyeeHfI/m
8APdtdn+vtymhjHGxa1jOYavcepssqK43S2Ya3C0yhc3vKQHrKcajgdnkdCfXb+W
zErTvNAY3mGMBC4JTBxT4nWUoWGkNiRpX6G4XSvLVcDIRACWems6HwMWtMsoCA/2
7qI/7v2nAa9eeHx/6YWjM515o3WMCaPlZ2cIxMDHqGg+JixICsjaYpcSm0eGr9hy
Jev61s4yvuywg7j5uk+2yUufPgTmOGSCnmMgd6X3uPKqZ3NNJcx3O5eZxXRjU7zG
27AS6kAddVtXaRcsCzfnndSUwZfXS3UQow9kz67ziTkdsQ9wD6lMaAUg/e+kgP+f
qauf74me9Tt3qrrDjsqpFUAUi97tYZOfj7ws2jGu24kxu+4vyQCLwYgQ0eLoB4MZ
ZdTjr9ORYy6sE9sfb3DXOECXUYGiWyJyfmkrdn+pnabte2IfN994xkZwWUmonVeq
oXc7+Oxl62HZ9LLDtuKjPUzlNcCV8S7DIVB6I3+Xn0PBRrLFgrSjjl9+SRrre1IB
8jj5WKbgqhvMAIiHT3TteEExBn92B79xwaZqWs+SNJRsfn6kBvqVY/GJStWkLXy0
V91xumSjnjOemabnbcJq81X+O9LhFk4G+iymPsqCzSn7Z93PctEXICm9C78n8tGG
p0WDbvgzfs84YJbciiFJ4OISoW4sWN0kboPq7GqmoZ/sRInOzbpr4razE8ZDWsJB
H+L8aouIoDY7b1YTGveWW0UOE2y7r9QIPAHMVHc3nnYXdMNxwWbdV39kF4LTo7nH
XBFECAMZhwfYpEPGFqd8igzpMtDSjMNSyWn9U4Ltv31wXok7bte1mlHXaYdj0zW6
RyKDaqeLhB2wakHSnmsep+G2HzRIM7fgTZ5dvQSvsQNpQoGYMXACpwFQO7k1xjuh
zIpnKB5dfOnyHyjP/eL2u+oOR8vNnuTXKRdJd8djTB30V2EFS+9T+mEh08KQbest
wNjlDQHuQqKSe5fTxJdmF3rDIdJmnyadEFj/3AMQ5av/kBl9ondhUDzpLMjfiir6
5WV8ai2CdUQCqPs+s+gDAow7XCx0RO3fn+LhhNVO9OoHjUc2K7U8cUy7qwPn2Yh5
XPOBpedUJ7qJqJZtA4/fuxi0Tllp2TeIH06WGp6szglpnsUVZejz0u2EA/tcK1xz
rlTbUh0+jdjY07bVy/c0tmVAALfii4gf/YZmcxdU/DVB/ghh4M6Vbt6mFr0+H6+L
Ak6fBRI3XSX/S8JBaul9kuth3/1orFbNhJhLRVqy727aMIvM7O8pNGD12c5I5IK0
zdx8CLpNjLN1fnZ09YdsNN+TMP+xIXygR0M5YV2zprOv1wbre4LKMREffq00dPym
7lG1byiaIbeGYldL0kWWs8bzPJGur/WVsy2bot7E0Qe4RnleCeiqI6V2+YE1NE4T
Ura6wwBq4x/PUN+jMNkmopTD7Td7bDlqZc0FljARlhnhShsf7Y1PblfO8Joa9qwj
P0c+iz2mt6c13a5nRpXroMW6uG0LaSFIAfubri5t5ehLvYFB7Bd7fMhtIvR4FMF1
20WeThPpF7dPOZY5I5ou9UVDlk3VvQFZmFkHc3PEMEvB3jW4YpuookRTyTjvOWTb
IorHHZd994sltIlY4bhmsPpKjoTeN7Sy/JJn9Dyz7kteiTmUDDyTYXHpHQ/xg7oS
YGIHh03EomZEvnnAqs91sfTIBD9038mHq5bTumrCuPXxPllzgl/B41w6MguYmwqU
w4BLYOCj6G68ocJjdT+bL+74LgT4DmC/yHGBOFSVzXqSzLv5pIT1eZWQPHGqZplV
3v3GqPl/FBivXWIJ+jsAD97EuOnb/1EuY9GSGhZyJ9eqHT6Ucr02glGc44blTZih
z8MHP4DFnr9Oh/z6w18PwUsQ5Ua6+8dlSg4Vn7ulmmsIHyW6Y/IiMgRVgg4tru3s
Pzo7yuN7sPHxDAZutFutmTVYrlAoumxd2M2miy7gTpv82T0bjNacNi6cCUSkvrhF
GiVW47pK53WxB2YZSHm7kBWsDgpTB+JGue2Qc3hZPqixhjO4Uz2zqs313fVc6jTw
fGPS01R0A4N/T1YpDK7Fg2Ps/SMvhTs4asW69FRlRzj/sWJI0Mc9qiBltaCcl5EY
s84SF1g4xxb3Rpz441P+c4KS4IEHtt+0vIznoBqKDTz3Os8W6jv4Vng3GWmpjq7T
4slQ4xkkKX8Xw1oHQaXuA9q9OtS2dgSLC7IDmlREbpWVNrGvJEFwdIpHbt+Meo/L
WrnjThElZj9zcouwp75nA33G5uFljkPs03ZQO4Z3k2x0OeunOz7mxlheRoilpT/i
8NXvIZV/58xTS5HkSz0rYuC8Xfqx8uqOQ5vFmlq03cbvrtXc3gnCSZY+u2M3tBp5
aQ2wK5yWbNhRDF/Y2v6fuYH9AWZSZSathCqZUwaGWMsEijvRS0Nl9l+5SM4Asd6n
+0gwfQZxEeL0WQOCStoyq9AZQ0kZXUP7MyGIWL1jYbAYw3zaSR7RdbKXFPX+v0vI
fhl9EQmS7sX1wDkmkNzLLzIYo7otuo5Y20XGQ3HY2wkrbhORT7D0JgybFy1g8MEk
L/QVvdR51gSXantTymtp+WpS+KgeBWtRDZCurtUicOEWbtDvRDV3MfE3+bq0aFYS
3SjP4R3Wc8MvP3F7R4xp/0UCUIyWWu/PiO2P2Nw1EQMyqWjGt0R+x3V27/VXAExZ
zaAlYrsZJjFlEtaQmPg1l33SbYO+Ny8HV04vMwPO0oNfRxSJTOW7J6sRdNB83Kt8
4oRKpV3GZXPctp0AXbPeR+yR7caIYncdkarGL+4HiWPPUiqi2jdstWYAFdAtrF+u
8ddjwHIP+xZC4gbugKZ+TzDCq6VcSQOKyyuoIfN/MHDYOnGIsCB+pZ9B1c8+qajh
S3p7Wd+nqZT/RvXtPrU0s8tHGcrHc8SmH7Ci19oaKh6FnRpGI7LYbw+bbzU1sp/K
d+vukyyvqSBh3V0arQIiFkUjkZiKHftgAPEfAoLQ8bSxDi3Rhks293ZKdEWXEhDe
PaNKfcXZyvTZF1yrEmjsGBgP+4Dfus00Et5K5S/ygdo2svBYn74jeuygTJbdDALl
q+N00VxC+Ly1o4kuoC0VprsHtyKfwT5/ngff3o8I3dJbM6sB2ecu7KZFi/J9io9m
0wrLKaUjWHABGqc8e/h8Ho5ar3BL2eaI6kJzaT5g35U78Db0IgLyf5JQA+9CwJ6/
yu5EEt3Ze5Nrh/CdMrCcNNH2zh3LR2PlCIcnaPxrXZF6XEmZe9HXFCGQm67Hscso
Ov6AujA3Y1fDAALO+vBa/onYHZUVqfyEDs785sqGQHnizQ0jAPC6mV1IKtDGaO5n
MNT6DeSrIZuOzn3jGKmm1PJFIYRlY3nXjpW0Dr5JGxf4dazL9zSScYRvV1RzBzGV
ny/gAXV8yF3ekIQ6cDXMEmkclDbY33W5W/ng/LPAZeY1aWaYmTOBmtlbHEYJzWMZ
OsJEXAQFaUlojeMHtZpVEWsXiPG7Ky2tttTbd2/VvG5lGa9ldaqWw2ydzaXctggU
xv2mA4hAKHZwNw0V7mjps9Daz9JrxS+EAlAd0i1aUK3YxxkCt26iTuCmrkN0YEI8
FvcOzNKncChvvG9jOqBUQk2m8QT71pbTSqk5K2Z1jt7dNduDjK19xOX9E5sw1QB3
Btc5YhgMudB6Fe42ksuP01XrZRhNBP6ScENun8h4juJxD4v4bFOuuOlxCE2TsEx9
doJ9n7Tm/k72z5y6s2EG7a6555UF197732W0tPKRZDpiisF47OK5KjhOYAvJo6bH
Yhg8w7FVuqbpGrkM9oHNlIRv8b8Q4dl7DBVf1l8cpFEE0wdQA8fRsjJnJtm/ItMZ
aYuVOJLuNlYPz0LTrgE4fVNutjYbaJVGd9RJmmq056OYuow3rBtY9DeSQs5+tMpS
KRDh5UM7e3f5Aq3ub1vFqBkM8ZF9W2Qc2+QfaoRiKAOoiQmC1dq8PH1c+KEAHfC2
JWeqBRTOGoRQxD8ivuBFX43+6uhpmbQ9/o3NwPXguEYD2Spc+uClRj0dRbhW48C6
RfBIyb8aOo7NSv7BMZeyJMl4AiOhSGu2ys52rTHyroKkJyECdSjQ7xBeqeqqC2rV
q8wcA58OLMeh74ctefHg+nvAeQObsK7L8EXFNvY+sSooc8hXLedrc/xoMlvrY9Xk
VjlVpJNfQAmdbAQsV28yk/S3T1e1PLZ9o5f9bKbSQMH/TyOsY20snk+UNnlukp8r
p8FhwyDuw0/1lLxPQ3kWqBqAu2+1D4J2M1AWYBSJYlBL2c9A9/MHhK9+m0qLtfHX
91edjZStMUSMAoh/Iu6pH63P0bl/blt42TYM3GXarm6hKp9gAoVXUEKSejg3L1/H
bKQjcBpqzMXZdNI4UEWHeYyrnXFWUfeuEr9BE6pr00kv35Zza2cuWTrkj9jjGPvI
5se4vxuwjO6yryhvhhrF9ehMn4ZId2DhCf/Y2k0rG1MHEcvkZjJgspcz0GBi0bkI
lbQ6MtJlVgU9MdbquBCttRXvhekkXz8123aHGVjX6+1PPcVUPCtOXgtrXFrlxi05
D9XlCTujhACJNNFv3OQC8YxyJc8jOswEg2Tc22BA/FxRINFVktn/5XmEPEB2Lmtx
FAw5BviB7SA11icN2KKtB3PnCawEa1aCdRtHoMvSp6/W6cX/asSCB0ptd1ClpaZU
tI7ClmKABwxwxezBoQ8oyKCL98y4516wGpUnKQQBVgXMtVYiJOwvqJfkSQ64+Nr7
4yGydei898T1eMqHobK3dGpwjulpp0iDQoVnQg5bha7NaWluzhgPJtsKhMqyuP9a
hPSMcEFPen7k6nGH6vIgw+2Xm+2NpsgmsU6Abt93A/Gn7DUZhRCaaO0e2jGP0uLu
Cfoi1XwTQm0zDKUOFhgdMqz8GJAbW2yyg2c4GFl+b7ANuhZqrnm4CJAF+i9KqIvG
BF6PCyg5kVTbxXfoHobUM7UfHCkOHOgi1QzywEMkmhC4U79KPc8IUbEwDcZ96/vT
+NrgQKd5WHfC1d/adyqu2/xhhajx/0E/oZ/qft5kotVzTaHUZNCmxZBLwaWo7hOk
IGKgz5ekR8Jp99eK/ZBqeIu/jmk0WSPGv/bfd/skCEnJLe0volHaNnZsz0Ooiyxq
g17XoTFQTN9tBP7JV3SFfp2x5887dBo2WwzXEJwDXx8Hn1mTEzlMHqj2tmkNJGJK
1ORKyHwT9GuF+ctgSgL9IhyM6fQxdNm8g50xrCtE0IhK7AajGXF4SqdXXVf1BhtM
uQgcQ/Z6VXSmFzUov7OPvmsX4wAzizFF54vNRTEePJMDMwpjOgJFpL0XxujRDMpy
TPBt2+CYSOXutZSiachCU+ft3ZLMxMLWvkCFHy1UCGAcztd7t9MXE3r7fllgO8CO
ruQ5mxbBhg8Xd9YcE9WuA5zc4dRHW1CTB/FNTjjSSA1yXa2ncmH6wBApO/cjoN6L
pOvXXD9rFvvY4JlPGMDE3SlEg3D4Bqr2vNeOqWIj+1C2KmVHBcT5AVao4W8zHyYA
KrZ4BUxTq8iiiz81jiKtu4BGjVqs4bTwjNIPZSLyA4ouvc+7K6gZrhg7u4C7ftU+
HqGpvXJ2Am4Ji149MAZLQi97zJ9vogd0B2AsrNUominEakszyaWaaEmk+V3ZLs3H
Aj+62Ld6yb5ZXnjvrslgAK8nhPORymT9juo70NpgEf9MAGmPErWar2E4+bkRYlkH
bTilDfGqkBJCezyOd5rqJLMMjKQHIS89YCyVYmc+okIE02OgrqMRNJh/9whAG86i
sWeFG5MB8MG374Vh12sVEeOsHFdgRPkIL9a6sq6/nGzq0kGgfbxs3lPjBOia7ZME
M4BAOhBXNlp0iKKDcYettj26Gx3MrDJh4VE86BPtJoPQvEhcKWdnnqjpi57EhBj2
YJetRV1n/gp3g6xXNUQ2na7qpxQMDpmsAr98tgtwczCWZCXw/LAevN+C3IFTQRGO
rJTjNe3Mpzs7wfJAw9vRTVhxTGJABHjf2nsXUsEvhOQ1Rzwa01tmIaB3nMrNEaFs
swKggqM2TTN6pq2In5vzKChoJL+we45POkuK1VN/J3Y6D5s9xuj3nuOV5WOCT8CI
PxxYDQgyQyYdc5Jt1Rwj9gg7iIL35cdS/+yCJLr4C1AkGirYLyGOn21xqmnvdeHi
S9TEbGjQdx53c3wQdAb4IpXQAJ2uxXbFZYqpYGECOhi8Ub3zVWEbE5U6fbVOFquP
Sl058BEv+yy3T9JYaebPxC/zRny0kY7XPr5ktKk5yqwEigPfu2TRfXMBFfItnGSF
tsaKAQg4gqC8nh9MDMEEAKDzeo5HbaB1eUAuOzVans9fQYPyqQL98XVMYkASOjMD
DxGWSElxkJHuXksGSJk/132qFBv6zgxooxLm4i5pGV+f2RGCzgNRlxjPC2zs7cIK
B1SwuLmuh79ZZViaIQLk4RHBchUsVPmwMdp9ttpAlrKU88h3ztHk4T3AwGtCehEl
vR4sV/yCODppnNlwtFBFdzIanIZAGuXBg9TBDTNg4wInYhrIXbVYwOC6g9AeXF/g
B6B9Q+8PXC3OG1FwZBGFpUMuOQgxgk9mIx0jGR1YclZwqpTJjLGQzD2MkER7he4H
xuvqMGAS1gwftowmxzrWRN4BrdpOIMuK8eRlPwVUmG253ehRyJYa7YmOyGR/vF1c
27hIN33GgUA4f1sLHf9T60O4UXzyhffFycswGR8vvtCJmsKZULknfhPLtsNAe+bh
B9Nd+l607Z9L7FsCFnjXd9H1Z2jFrovMUMQpbaOhyoNz4w+yCrWPQZPCF4Le0p3m
/9+N2SKfZbVh9heJoGIhvq0d5ZlIDF8MSOgzIq+l4aqnXR5mg3UhFdIcETqtbfVd
gUvlm9Leo5KAWMNMG06i/EvAcyO59o5lndaN+j5jF5KhMAz4NgpaNJ903vffuHrw
VMkZbFoCSIAJakAqIUw+6jBpQnnHPYBIftb4voXqrNylm8XI9iK3k9FQinaqon7q
DpMzZtX6/OvK1YTTTOQ3a1/Qry6ikZcknKbfiargxApvBt54LB05wuzZvh48/lLi
FX6ZCU5A0DcwmLvpHCLwQAPh6d78Y2cjRVqPIhRo6mEyrgld92EQ7dDbS5LRV3GC
X3aJqOPDULHf107WLmIPtLzPNqrkdxMe8V/yAA0XM4grPcEYRo3kbJsVdnfE9IL4
CCVy/3Loqf32MEAkdeTonLSOx1zQB7pxOSe0Rwn6WcUmSnZyB0qB9uPrsjJxwq6w
NpWWJVhhxNrEevBMYeb3iWivy9JcJpsRwxYJaYT+6vfxitdUol9KtUXlF8wnQPAq
mq6V+//LIBEjFyDeLb/jb7lANo+Y0AFNAZFIPxEXAWb1f3FL1px3pOG1SUyKAimH
Xt7Jq4mCisKO6ok//vMvmYoHhIEp2e1APfP2gYlLmdpBnh1wXaBsO6MmbGWJN+9z
B2dji0rdXKeHaJb18h+IugJ9Bv3tZM6eZnIMRMJDxV1UMWm53i73ezs4ejYBVq9O
zVtMxCnJ6Ua4ATPh6tdoE1f66DCUVubRMzHA5QgVxQ1Ny32NIw6lFeNq25kBfqMZ
qLvIzIHnF9pZq15G0FaeeXyH3f1jx1d7Dosvpc6V04W1R7pp7Y/Dnz/kZXwvxDkP
sIKpuInnt7Vlcw70vGhrRfgL9DbzIfF2vOLX1x24u/sworn1YaDRwTk/MBEUP0yv
Gjs1/SkcaD17QhEKA/pm5hM2a16bXGSJwXaie+ju3lFTmsGS56Zd31NevbLXrgNP
ythHDDDITtS8ql6rFHNZIQXiX2QrGjg8oKjlUrS502JXHAvNrsifzIbaeYT3PheX
LjhXupbTB5c246hWFqPkK1H0bSLZ7+tR3u2A4o4YKtQLiN00SfDNu/dBl04CvCoD
cWkodkOYmoSiDNgMjh6jFqAH+NhNNJCAa3u0Ge4UR+itJM0t0G+M9zgUC9a3VENO
GWHI0sr20MgDQOTmK5/8CidSD4aDFLcl44haOQ9//Ntil4sXOGGmDcO6c8TSLn7L
ux1O0kKF7chZndMDzDqWmnd/cYe9s0PVfUfG556/Y28lneMcmuKabUILdrAo1tpY
Pc/+cZ97+DRwaAGoVgMJ3N9gMzJ5IiHHhwCOj+fr47YVyIK32++WHNep0Z+XDqpO
VP/exBMnrW9g0wPemDh6aNhEVhwmJBxhYZhqG3hKgARou1YIBjwjp1cT664+8br2
Ee5mkpcEX8fGWxb/S97HVb29+2MXMTJHg2gXXRJWgCr6PeRwKDugTtbOnBWUAbAa
jTD9OB8iIH2iBStCBfkOShmqWjmczu/N0dDWrWX6rk77YG7hUnACPPfquHthISEl
CviexzC4D6kiqzZawitbf/SBL4UWMrjFgG0JVLqBACJjl5jaq5KOlMQTN8ZPx65s
naF8V/uX9bSxy+6zHgV7NufaEjDi4VoQDme8q8AOM44BuktIDDUAFryk3lHwop+A
tqsGEzOzvr3beWFZbHHPEenUbIb4/XP8PcSJHL2fKK7k8trqViWAQw563eGIgrQH
SQzHopM+O+Oc8TMrH+NwdU/tJe9XJFnj37QQJbryGYoHGk37PvmF8ldy//+V9v3U
bykHWlJkVFWG708ICNHwqt/wE85U5wKthsNzm7xGZ43UJfNJEnwTrF/f+osKm5tF
uliPrqLOZ34IR20B2gooPUcBDZNRwn5s/16Yorjg4EdvxIFA8PII1MCktZ4dIvE8
dOX3oEhlY3WnkHWpxlHyZf8eoQxNtXAEzwtzZCYmn9TAP52tNgbwkZAxDQ2npF1n
dXWzGm8tjbBCGGWzt7X896DtM3YGIh8DoJpQ5FWLFURTtVbeIR4Mfz5+cy/Yt43F
FDxo7Pv8TjLwjV7OBKN1HgthygNA6j+7FAK6zVeFqpcHyzE86Ae64JsY4VurOeNH
ZhVa4wSw19btMS5f3wHZ1OMIYY9P2tZw27WTK5YfajAFb50sXAbi82cVrodOKdGm
WKPNEpw+KRXQcRWPXK89YJnxpB7CdsPRAbvJyYspF6o54tHPzeaMPX/SgXLko1NA
XBzpSCoOcLsT7PJEg25l8YhVLRNATUlRCoJ+5GBNM7ejSlWE22CjqevKEeAyeIPr
3OME+uLrr+0IknaJBdHnJf9SnQCJx+2j1StQsGuYJ42+OxmKR7fiCrjQ915TfKZ+
YaXKzqvR5udDnX6m4+WB53QrjixPfK7AMFbxqCqg7Vm4h2ZNFbiY6y/lkMRK+GY5
U+XWKdwF9z3T7wzS6i2WzrHxnMC9GzzDtHexuXxwFWpv8ohu8RnJZ50j6Z57vixX
8TgjnDW65CwOhInHqhMJkhdSOhzOKe+gENNNKC+8BJOBKrSGI4q43IbAqLwfzNZY
0/keBtbNpqmqs1uQb9JsUc6SMiQSpawSTBdViQg1zIhaicvuIh44sQWLnvpBi1LI
gC0CnLbTPtrEpULdt1zh670cFox+Zs/ZN1JTfijKMH4Hyv3MyM1ySp1qZbMihTu0
U8fbBb5S9T4rI12/HIcJq4rTqFboxM/wh/lm3RZbm/BIfbGpz4laElTTkQIDTfmG
hD9YD3vCOmcXT5urzHShPkXqz8Ezu2tx/YJ0P1YvpXVWf8FsePPFCAA4NRnRIq0Y
i2pQQ6DzrvfjvoF6+WdXkL/UIzF7BKnqW+xRgZQ9PQh9NtNir2rUoGxEKMBo0qzW
KrupBvOUuL9up9tvEqnFNO4TXEEKwaiuF1lZ5yLS5ybgDhns3661mTV/qitvVA4l
xwZOD01GzdtT8r+ZgPL0bthOI9/XQAExaci/l/5T/Pg6sm14DyoZMu+qQREopExg
H9Yp6mPVfyez4qyvrILLHW19hAHwuqxVRIkIYcrIU33nr1Ji8ib1YKEPed59KGrU
zhGBOmqJcoi7JAnMSYvQfbmnBR2hFEy0q1vJp88aHR47plu1QNN5UrHkA3LjTGik
OsV0/AnSwqy/zfZkZ4MXFv1OLIq3gw1Su2zFOCbu1pqWQKpCigPRvxtTz0RrF7dP
oR2i5kpPhE7BFPjMSXDKBe4YyZiDP4d26Cy4nGq7cTB7Id7SRRIFdTOirmsuU1O6
NTSVW+qgatlzJaP7aaL9N6na2TdFkthrkYH7oxIjfu5Ne16NBMA6Z3zmzj5gwy9J
KfO5itIKUwkAJ9VCC2Ah+++45ZSdK2DGM06U7FtcrTsMWYNtZkSzjzegadHmnGSB
reiI6gh5y4cCGew7qSn8j5X2Rl8jwhHnbizWrp5c83q7ctcAtoxNngHo+nxIg+vm
cAQAuxBh8kBbrXlmMffhUicMzwqDJVgAyz/loJrBygb2eORcx+t/Gj6PfoaF7cn5
wr7cDv3n8xkxutpG4N4UkU93BVnqrbe3tFJKwlPHEc5eE6vL15eXKDiAPSKyCPhU
J4yh5FfKemswBmAMCUYba8RZpjKTb3R2OKu8x5btV80D+wpQCNQPMzaYJv7t+14h
qdZaV8k89frusreKNVjrsi9n2ChP0qwonv19dxIPh7Z93SZ8DKhRR+8fvl9apoRe
atFRzo0vRk+8DBmPtSM2BArenCvPMikA8iHEF1zEl7a/FHMQ4jxzusaMBfK3CJOq
asUXKsuku1nC8MVeNojQQXzIvGu8p5vIQY+cQ0TtNs3uMD6Ifz6neoOIpzPuuFe8
EaRr9Zfev7BsgIl0ahic9J4f3VwKTfWQ3SikdUYaAKUEBA+rCzE88kN+Soao30tt
27glcFLXsRhuayCF3WFs7+s4TndKIx/5gNxgQ8b5ilxhqldTEVZp57CIA+c1o4QD
kltAiWV0g/NdBSk3Q3fMoWQ3tSHH0N6298BEvdI5Lkw3unJONl0aCfllaa4pHVZx
2WgPqlVL0CYDYCGBOKeRjQjSBUV/+V+tpgQkb9S81uVmWcA80F2Jq6OuKXmid8pL
6i82NDhbyFGeneJ40ZxoqxrNvbKjd9N1htoIyWSRv46q2iqsX4TWS7OiBlcDkuPd
jxScRx2GA4al+XSBUlKxfza5zinX+BHFuLzu6OQJ3VmZGVrkZ9yYdKYLcvoSwp2/
NV6aMxKZg8lEV/DxTvjL7+nPEx11L9PrRIhPYUC3hIzSEmUD9yB70tpTRmaOhqzs
l/aBDIx/7e9twsQgZc+LPgp5nbRX9IMCKadxtMhh4ATCCJL4drqNpvivLSROq0xL
ibxllv/LuJS1gC8zqpxIkb7VdnfH67sdKbdbkSJImhOEn7mo0zHIe+m5iwGbDQfr
XfQp6IcW9gM5UgSfR/BSx8a7/JwHcd6q85OBulan/55GcSUTYEhTKfwGwQvy5V7U
sQH8mLsoO/STQ+iFuUHzjKsRWOa96YhitDEGDEemU9SSPVEU4dcl1Xfk2/Fz49B1
cmRIV2fjkwAOFExsIoAJvPM600DKMibnmgAxBdGF28porUmuX6zKIBRQkXO4zjnY
FAYtU42JE8GdSZ6RmgH3guJ+Qi70SGRtwryaqQK8lK1VIa245MYkvq8AKwDGLJun
HZGoYCLVqBL4a51eWj5rn+9DAgk4wbMS1ywrMnkTE+ianQnGCcy+VlPcqIADtHEo
v9tL5wDLoOj3bBhss+PzZpTuWcGmkum89nNuxUfM1CxrrVMeAvzR8aEp6V8n5M5e
Pk1v4DCgeGp3Y5aDUwAMYN4lDeLpa9jwmijLpQbRSNF2c+jp5Gz1XMi7xs8NQDxk
Qm4VA2gSIfNmcOocj0pMDuhoAO+4b/u3yJjBOcgAtcltfRpikyXwX5C9rScBU0i9
34MV9OvT0KQPYycEbxb2Xpt0iAO83IAtMZF13bKXsAy2mOd8PWC4xkzV73zUqJue
F5yg/LXDYVit1iTMOACmKNi4pc/M5C/PGg1Z40Xp1qusG8HLtcwdedF4w2yMsu+6
h86jTFg76zxktueYxbjIGnif2Z86wQHQhrAaEYez6f2fykmoiHH0+6SBfjVve6UV
76lh90ywa1de9Lktq5cYq9Vxm8uu/b5y6xmAfql9V+vOXAECA3Cw2+v0oaoTB2XV
zhb574Q/RFXJo7yF23kFOsfHIJ7YyNTXehfz2eDO98J90Y5ch+hPTMJkAL8bWIR/
tL5v/R01ohl/5SlWz/i+VsDKRbebW3bMwWUNGQAGXKhhSWKNfg+ZeA84oJeWXQQC
ejLAulPNrs9MmIW4yUvyAvBi6t0q691qjgemDDA0o2fmjZJPxS19P/skAyMBs/+k
8XXDOO5yS+ZTXKVzumGhpDKYSe+WoNg+OeKjFoUuEzxOqUOtkFne8HGGh0lfSIH9
fxl0mmzMOCoi3o0qD3OyTRaFG93BhOnyzxzxrH9AYJjPXOwcaaDc5DoB6rVqBpxw
T3MosUj1JQzqqZHXOQDdVyibLYJeG1IXbZV0z8z9H39kTxtH4TkrILELXQr4W8vJ
vkZl3r0Gv/Bfc9L3JIMVQhfi8lpt0yazxE4iXQ2huise3laqN2EpXsQSF5Os8p3q
YTMZE9mKMQbOFnEO/kAg7FjRAykrj7/GOL0t3OequJtnTIT2M/ByMLk+YDMiCn3N
/1LZpbytGl7eeNWUaf6oKQhyIVTAN4l6e5eH8ngPSRnn9vMzI/73pOuguD1ZWOEh
E8Kf7++gHBo8mU3T6IIPixy2wYHD7WBymLBQDk8xRfXF4vlzF0SFN34nUjlsIm6t
kgXd3Cm7QnMUyQeeb+9c+npN30L7vpEIaozY1FzrXsW/JPMNifgMA8MT1GWn5Krk
oRS57tgk8rtmwgt0+ZDVKRB8cdPQbmKVt26E21pnYGQ8yxqt8MnLO5uNiSp0FSbE
aUReeNiwrUkj7K3cTNAUyPvzl5WDy5sKsP46yCI3pmcy1CrgugAjYoIr9vr0wtJE
tjJJwJOpuORwxxSjhHCgAtbbJRU0MAbUpxZ65gCi5EyaGfKTDk1p1D6xd3YhKdXz
I99qChSCDcYYvjCC6g6S1hkQFFmvxxqwfp0hJteWIKjfW0RE6Xr/RNxFZBgIcn7t
NOv2Znv0Potqb/fqZhvzChRN7lJyDUDwWCwFtK2Waub2LLT6e433UpauK1lar0+g
ZXoKuJazdscqcu/L1jtg2+qNWzxJfqsWRlVY5YpHf2UKMAiAgRquAL6bgb3K8RfU
T6W+bx094zY1JGlAv4y12fCiV5brkG0lDEypjsZoZZa+mDzQqwtLslGdKPShtHMc
h8+9VLy22eJTGttCf+thwjgKzcUvc3/UunswAuCnR1KvSYs2HuZvbU9nh0pY8N4s
8NZHtgKFt1tl1vsSJhbg4G874wvSBffYdMfjLi7dOaAuPNv4JGL467BeM3wlXZmS
BHh1JG4svBhI59bbqeHbYvYVpJRYrLOqnN7+dppZTSYidvl7yYSRYFemvmEBnBhY
ApTIadIZCdsLuVn3prx2bZzxFlRY6eJzOckT6piN8674+8iqy4tNIfK8DRNKGhu0
Pp1RyRa6eqSaiZCBz42g4plsewto6UJpqOGmyAe/T2Iq0bCFZ/v4gyQscLCtTpN4
h2QKe3q5XD4GN9TwI6IcmbPMhlEaOoytye3dcHxV9IjG9uY2xX1Wary1Cb1Y8mpj
z8+c2SHE65wg+BMshQSu4DKDF+2L32XOJqs8BQ0CH5A8LEyQEDiO/899o4EQ/nJU
4Xg3QH6gYemqu0NdDI03ATPjHKcC0V9yK1zXqhnH/z7fcIeNxCPVoKMywyX9NoWW
XMuzNxpfqPF6AspPwRL2U1nzrZrmoSR1tpjUKlVYMWRR2JRPRY6OH8dHFN1saFUC
tQ+fndws4+afhQF7KZ79ReyDI/KEm9XYC+EMgF7u+XEhW1b5ohd52yUztEFXNrR5
lMf3sjY+dXd9RmIEy6TdvRrw587M1br8apncT9hBCkSCiMs84g8n0kt6jR3hWkjY
pRX5veev7D/3uoyu05BS40zbMXhvJI2rItPmUY5wYY3asKxQZBpXtM38rrcQ6lNI
3kNLV9dNCowjFM7iMIsbO1jvEhUfJvp0kzQQOENfjepJBXnvAM6TkfuLwKPAH63D
Pjblb0QiR3PwUICs6HS3JQ6e+JwPjpvHSQ2f55BWUVjDe7TdQNmKoQo2mVVKM9Cj
CLjpshy3sBpoGB6t6DvK7tReWbs20MdFREUrHRNWjTCLLMBIXOYf3MR4Qo4e5hT4
m5b1IGZMtbZwVvITo5oYc+wk2B9xzZey9tkhUhlTLqz/Ai5zJLFPHAZYdJ1UgZ8V
tcnncJR7O9Ys2tXOwOlrwUetQuBNbir7foUUiVGF+rszXbpOeJRNVJ36Ad5EG2PD
JXy3w070ze4cma1WXFWc/DstZaKxz/MjMQ3ZCw9gSNYNAvk8TossDdSLFgiSphHV
NAcKT8hBBI6Ses/EcXPdIU+hXJRbE4Qk7eZq1wZbVERam81+5UaCwfw9ftyr/PJZ
QFwb+jw68WVnArzMOdGXvvJTzxHyfqFumlGiyW0sJd7GNMvmuLzbgqF4Zt8vnJk/
s7bCALM1vP2ulpthYMwe5DF61cNykIBc3ftA6mpVylpi5zs8HiZqUGGiZCjDVUmI
c6Of8jZ4XYRMD3PGnL6MBjfkOAbtDLg0DIlSMMLKrvZ0z7BUiMZdtAx4gvgwBdxe
jBlinxTnMUoezUZHirO2MJl0RJMZYlw/lYklftZr3bOWyEqbi0ruC29qtQYpxKsB
UwLAbU8Jr0MSytQFH5J8EcDwgq2CW8AzNWvzbFw9sSPkxtqQ8+WOwbX78tucbBip
RpT+qdKPsZfUvSvsrLn8G//TrXR10TvAMkMXCSkEfZ+wEmvhSzj5A8PsfMABCsd6
lV7a4DnOXRrxAA/9RjPdlUaTCLkL/OkPBIiYctmd/NB95v2LMq8MNZhua65FVaCN
9gpSU7Y0A40RvBRiXgCEYQ6dcgvqPceJeGug262Q39RiyySvo8vf5W6cX+ZujL24
g8kxnp/pIP6z2ZWvllIufU4QEIYNzQ/n4sMYIsuAQ0Pt1aqkhms5/i2WjmhZ+tV4
OfpCVv4PuVfyUqa6US+we1q42PbgIvjN0eHQucQMwjbrbIwIlFBp+6x0+xjT5amM
pubRgM1MrDBR5rhocTjD1ARbcJUeyaRCnkUkd4Yad+85p75V8MFF03MMDLmKO6A9
Bciw+aDzL1JAlnYpB7lESQGYubMn0tB8zKdB+3JdeZ41L8lCrWLUXhm7dMeGqPFG
aFdJ0wAujiFZNjQqAwt2JvScE2GjSyg6MACQdIrEQ+RiLMoCMXdUbfUimhI3PGZ/
J8h+iGYRuxeU1eaKJoGqgt5+dirAY/dX69QamM25HEGQ99pUnH/xkVerM5bi/e7H
3Zixrb9zUQmaDNNmMO+WOrtw/lf6dkP+N939KIS2bqZaeIERnft/UUogeIrBJFhJ
Hr6YOOzdqTeRSFTpWVbUMrUaMegKXSQyBBisw8zeqmvpYl79N3Wg35tv0M8Wvv7W
0PAk8OrJkl8CWXiZpHGCVsUJycY9ejancXIdr1giBtJqMlXTvb7y+/XtqtaYnmMb
MOY0vCs35uz3KNJh1laKHwiJja2+60Zl4qkwxa7+GPr0nHyothcDN/W0eqxikGV1
rOE7TwAvbBlakzeP5ISoiyAUh2GieMjX7mG4FP+m87/dOsehepL/Rz2ooKrRm/Zw
cpEzEo8sAFI0ZDzzD9bhWID7rnHyuuHwYrl8ab5fBbYsrip7ZyeBnj//e8U8+Iho
XUJ9t98A+VU572JZNiJ8Ex2OnZIDQLoQiVVSWHinFGi9Q7FOea3EewKoJya3Qm95
N9M3cZeEjDWWdNb2jXlFoXcyRsa7vDYu5ltkJMZx23wHbVrnpimThBhCxRzyGrx7
B7LdBD8WiE98Yx4EDg200VOX/dnLa3J1nmNKXmCwYhBIj1b2HdgBdK7qOZ15Mq8G
uixx5ebY36Tk/XkYGu97W1IGe8621W9JEwtVo2DQTZFP7cOnakBC7ds02QkWKgof
EksfQjHroxxPudEfeX/kKt5YCc2Oi6TG1XQPB9TCgHWdLAwqd26hgkp+TC6qPgok
g41nunZy+3zJE3cRHBLg2VHQuFgLlWt5p40fK5YSa5J3RxmSy9m50/n1T9o9GGft
SUHV5NXiUggoeMjKnKhRrICm/WLq5LCHTepaKDuA2asP3ueJ5PwsMXaV2hR+3JDM
I5AGkrtv1YHseH3juMX56dyKurWs3DRQo34MRijSDeG8JZTtqgMMouPYCZk5kDtt
hGlyXKTis5MQ2DLH/cs2aYQRpWl/m8ZrNR3QNNFuYbcypl7enj8SXyaK8HyMin/H
eJPYxkfouvF2iu62GrBR7bbWDwXvTAqiwlLESjnQG/h9OCPbB8ZrH1dBrcA0/RjS
J85RFN9e2+L9x9D8migFSfZd6ONxjz9NnxUUmvIia/LurrlpnaZm/NVQXpwhijEw
YCvbn2A18eOJ1NaNgsRXnP7eG0KLgu0zlyvysRTENL+aSWoRX5B87MUqtcS9dfS5
aYE6x65oFakcPRzo1etxhnVztjW1spdDOtPJ/NwTcYltdlQwxmIzArkE39lfQ8W3
8THQrIEmnOHKWNYxDtpV4GbcXxv0Iya6m1Wb/AAKEy1XmRMRLex564o6qM9hz3x2
SyksAARwK09+nUhh9+hfj2mW7ynA9T9ZY3rsRO8Dtj664nxYAg+HJ8ijgTx/ucq2
zDCrFsNgI5Q6j0Zp8c0XJWoJU+4Q0vdjgdsEa2p8/JbDW3NGPkHZUUocEAGH/dsP
RoshkEVLGNnlt2aqq6EGCA5HIn+3BTDhT4JXLy6+aKIIAfN/10KMrDPfrDlhgY5F
TQSvsiMEEKQSaMVmPYas3AYMB2SPUsDRO6IEM18tZZn7nWniucPfermay+DknS7T
pLXh1jts+odmAgzwFFBhvzSmt8GkO2wAefh37kvn0rUE0Epjzigu22CeNLju1ZPq
BdlN2LfJqlZ2L96D9xDybuShDTureQ5sQSGH0vS5eOCXGWC0jagI9xlkGMNF62+L
/wkI0l0Sg818gd3YKuryDZBcLorKA0Z9jVj6VAhFqY76xPaBdl1M2AlaJRu2vHYW
1cb8O6fuzJNMz/qt7PABRMCiBbPnHR/I4vqNdJIDlb5uvWASYRPKtE3RuOHCdPYj
bru5HcvMUjncKIotanD59HHkT2W4t3Bi3NPWSP0oYkQQQSaZ38xfuHVekc/EzIfa
ES+L9xvj9ncLZjBPKmdwrhAOSN/BUB6IUNVW0RN+HELw8Yc6pkji9+pjIMoxfXSl
9+V8APf/67btNTt2Ra5mLvgWCXKFQDc2sVTE7SXF7QPQOtGrE5Lcr0TLBKXBLG3z
dkQwcrMqi4hOYPwmOIdgKL5cy2lL3aNedCB3opgxjFctdUx46cJ332HNYYR2wa9z
4KuYqp7yGexZLAv7VlHvrerSLXUD35EYYN+RKAlGcauR5DdbVZ9mMPuciGP7pIBK
xVXdRwjjnm+UpP/3rEpfTs2O6mrm9pf7ntsvcmztcvz5g/CAQjSknAjl9TQL8t//
LselsBimDHiRhCqizockm2Uo3C7azV/HEeo4BrKr9ot0jSvhUwH1isf34h2D9pPZ
F392gyi+9jUWo9a14PYybAUstRqMxFW3qLIyTBKDfA5itwb9toBcYD73gw0CJBVc
1HlOmP+FmJ349/Ua6irNj1yZnCr6n7UcXOlQaXNB8kK/PANumW0GcqHPfG37Fqmv
GnqAq/Atro+MyPZOwi84nNK7t1WuiqlrBMdEAOLtzoFpUht4eNIC4vZOAG5DG5Ti
312z0wOio9IOUUK9q3Mwuq6jjVagUaolbKEQpQoPaUGILdfcOzwoK9FmGMv7p4hb
gmYixxWzEYuh0sSq8KDWP++wDuvRq5+S/qFl9u8KLbG6XUeAy1oh83aPekTqHbJk
QdT3eNDK7gExPiwofKTDS/Fk6tEtu2iclYLMbfeLUM0J1eZfE4KPOWxPl85UfrS6
Rwy6bGnfeokdpLfXmke3qGgkXqiV4K6NEBgCPEHDiraxr6NPuTPEHvZZqMzy5bCm
4WCeXCc8eA6F5FDAKHTy2jSps1HKcOH7PT7f3wrkvUScRmzSuqxGDffXe3dD0zPX
ZmKOxFgnaH51kiwQ4YalQMpab/eOPcgolfWr/oJlcGevIxPePHO3wnol6jGS9yR8
DwQGGsQ3P8c/gkKpd20KCrCsa5zIsSLoj9IioIxHkqLvtH1LLOhS4KOEqF5msPvl
PKDlnE/vHlfLzbCLLw/EkobvzaRe5RYSVBxbDXLT0zTT65/OB4FCg5ZGP1h+EtYo
8j1WfrF9EZC7RM0MAdTzAb5/LWxIy41F/dMciJ+Cu29XQ8EorobCqApReCEuuSCD
Vc8KT62A+ev4U8FrVViDJjoD9Rf7QetxMQY+y9jAGjuXhvpecUMtmEi8n/JPm/tT
QKLnpOUrOmNcwrh2NdOFUBWpxN5RO1KyCW9tuCSxHoNpd/vwtAn22ULBiw+UTfkK
ai4xRB5MQ28D+Di/4aP5jAMDqGzqFztW31/5ly1xrPCyWAII8Ppk1N4upZnpUZ9b
da9HRIFgZPbX9r6XvlhnawBwtQ/RU/bPJ7mrV314iiHrWrbd1ymWDLbOM0bAIwcc
lzEnT9PLjJzwE1Qv1NfDIYNGXqKWqmqbYj3JCjEW+P8fEnU3KDb3FPTN0Mb1YRnD
RZptRaXYorS5DB+y73DuBoEgEaiNihqiZJam3tCn9qbxNQn/jMMq4sVcxqwnyix/
u+sL41DggyGj/RYM0iy0SGqhwgdJLjyANHc4HudPnph3TKxcVKu5Pzu2hDofWixG
FiXLWA0MYLo3ZQmibBp6rSBLZ2p81bxxIfcbaj7Qvx89x9wuIMxhXLQ87219T9Nd
DEcC56Vu4cMTtpYiNxVLNGCJ5JyrSqPtXsucX845Vh2KI0vgkwmIoyI2w8YcDSd0
lfFujN4qtdvjmH5/xONVwJhv5glRwjw745w12TzB+J93v5BuaVG3RhA5Cxoktw0u
BzLhKj4ecQLtp7P/MkMxhjwRbK8JajJKZqvr6520/9JgWBIFaSEgFnaPAXqwCy2w
wth2sLL/XUGR3yNQOQlPMMsy6VLJw66Ni5KMVYhwQZExXrPIXHiwsM2giztXgQz2
YLfZ1wnN2Y2BAROFxAiSai0qv4Qkbi2OziH8rH/ChpbIH1o+ktwED8bG8P5RhRql
AUhsq1rxGTv7Skf8OoEeD/1eZWZ7fgu17P5tJpfEQfoc/l8FcNBJ4CsedvLACmhu
sDLTyhfneiZhY1H2jSKMiu05lyr+0vkZQ3kb9cnC7jR8jUU/7jrRI5HJElBgDPZs
ipMRWzmaKBxX1MmypkAUz1obg5SpHep+//8nsnQ73vemPoVpfiPINcNO6oBnJu5g
nNjTvO/Pk00xnl/bZJcHkCIscZ2O30HBkVIhMrwsuke2BT6xyHkvMRt0zU7ndLjN
KE4pChQO1v2+GRE9fgFbTU0ZtcJ/uDivkHlDe86OcRWUy2vev9BEYuA3VYgmJtxL
UoBB3FSP4Fc6h2nTMa+Bf8GTQYGBjYBtzKKbaUzEudRinlrvB7+a9hIodvO5hu7K
rUwQko32NDs+wdjFCWupcjuK2Z91ig7TZk8JPa4fjUt2ep5nvsoh6183NVXYIvPp
4jQTsbLi5p74wp8EGrSpFMgNO1OmSA50Gmv07SYOEBDiZ4Nx4Ncul+mrbL5+jS/a
pfGZ2ZHXutB11VcpmfDj9alnwju6Zvp3Qgw/tDiNPXiXiyz4a70a5AZJ/tUSTImw
t7iLZFVXuiHDK/im1r0USugr9safz+xjNg9p6+Ss+6Qdw3SpsYsa81201IIVB/DV
uto0b1nerUNfCdNKuMVG07E2Stv4Jm1LOdixLEk6gUw38p7xGezM1P4em5jXkfoZ
uj7CwE41qkw/skGPgkArtOwBLyQJz/ZEJxtqguOhwsb0BENPtIJnshZUsXeGHJJv
X8MZDovJKoiKgID5Vcvr5n5VZBdxsAsuR2gSJB6eAVS20rf/vCvT6SH2np9OYEyu
QUr8vjUQnpxd9XZWvYK2Scn/q3fN7/LRHg3ZBdPZZALBWPFiaAVAnqnEAfmaSFNW
SywD12JEwNIix8nm3CqMPFaYWXXZ92CEZx2p5Fct/rrqIo1x8cqN3NWEvGuzWWxe
mtixWmfilRk6pVYR/1DYWslnkAQb+dxRAJKT6YDygRxI66KwhzvxbLCvmObDhug6
wDvXWBhaa/Bf7AsRisUsPlVdXgfJ6QY5g/axLVcAOOcbqyVS93TZHU/t7IeANdLq
OVYaE8J/ahtRZbBJzVRTi7FNkp74ctAY/UX1KDiL/6/Ul4c0ajB4HKoHY3qQPnQP
wLcCv1VoXwK0n3Ppr/pTwiA4QXWhzLq8099alsSm9TIF/YwScYT2CaRkcDTP36fB
fqo0P4aSrwuW0dyIsWcPmQxjSYMtO/NFxishZ2jQT4KMLk6qMcz4hxbGl0Epdejg
S1f31iI0Tdxes/wu/wQxmYYXoioQTu8+4RiTZybHvhKsedxgPDh2kuPhOs7a+tBg
7yzQVrrbIEA8noryE3AHB6BmWJ0bTb1DM5k8pRKIUnKFpu9Jr3+EDe/UflirSiVn
YetCXmBRTnu45XIkNcFTIqY3SSpB3dJ8IE3nOrzFakvTg7co7R0cO0yAMlHU0VCv
lprfSIjRJDwLASJYCNd9eZttX/iAJg4bdg/bXi1/988MEOgot4ecP7f/y91tdex+
i1Go1Ijngmdk/Ehf519d2HmptGoRpAXNdDu9IuD3tPcDm+CtwylePmCa78xxizxf
qI0UTrKQChX92jxCCCDYH5kRcx3JiO5EdKbo2yxoRwdtCic6DI9ys7C4cNGDUDQZ
S2OqHqhKvHjtXypMhm2T9/9zuYYGaAT2M0X+w+OfpiNnbTOKqqTkjZqx+LTsz15P
k8HJy5JC3pLwFU8/euSe4ng74PhFHth0TsuLZVZYK0E9NZKNjIXaR5DAkBoHjB9W
04VWJ04ZORSGLfgyi+9dirSKKtj5o5QFLWCZjMSgOfMN3/mSq3gv8TmMfshgUpBi
0KBhN12Cc/Gc33/lLMx+GkKae7ehjf9962X1YCdvQncKSK1ex/l2Ei42UZesrLcy
ic7tWgaQp8DciFbCP/swa1JwmCFaTkE4Vvc2S8cCiHbSHUO6NgWexIEZqbhF/CSJ
Phj0OW5xLbR+L5G1vGZBkCCqpG46LPu8aQRQofyBnfKtd5iwhqCZoz8orhWUI4dS
L3M2Ou90v5VU4o5rTgqOeH1HmkjCGbzRQ8N29AOOfRnOPEo1uzdWqV/bLuVaS7e1
eDeIcBQo5Hh6v0Qw7D1aGbLnV95zcGJyC/Q9RBab1uqYwEg58hWC5LvnpgpWil2Z
5wv8w1plno8oAE4ey8HgvyOlLQFnH/KMDmKrPP91rQ2nHs+oW2LZOlaRHDveKuit
ybqBF4Yk4wGswVEWN5Ope/Eerzg75IRgKkbsJopWdEpt+WLfMAzsvH7TpSJ5k298
sosQER1XK37xubv++nX9HvupsTWhd+i5DXZQHTikT/M6S16BXENaq4g3qNdsRMc9
kP7asL/6a6IhkLx454No4OxIbvDulrxRlKd/nZQaqImK8i5e887oxXE3fzQtvJXm
a2Azcza/FNYSLp4VixJJ8/oiRqFZspvpED7FhydLn6RCJdibMR9iLuWMizUHdNW4
JAGxZMQc3AHuOyGdMO/1A3AS85opK7PYnuvzbc3kdDnUvflSpwYz55w+J6AE3xcd
UQgvlolr5gOa5Tgq5SjqtOVMLCtGTh5MJ3p99YL+AIVy68efwJFRavctEun7Ij9w
Md5u8Q2pCTwB0qAYoNb5jJLnHgDtVSmQy+fklliPXC7CYdsP39YOzf6qPaNEpL5w
3MhzlMc+PUEXG8RkPLqrNG1YsJSaLY42ts6XdcwpWJnxCFPljYX/TavL1UOnzYgh
DoDfz/F3QMHgw/aLUN8YFB3+07ZW7ofou5hTyXUDRSVIh1v6BL87J+sSgHvHYCTy
Xzg7OcJqiSUBqTDdVlqchr86kTIiqXj8FxjaXKxVXM482fpIjPBZsmMmcag38J2g
DzAp8pwa/n6GiH6Svta9aE+xc9xUDTdT2TqIbx1TnZLgrGM2WdmDY35dvDqrc/Me
lc5NfZB579vtlTS/CQsvbAb857nTrWYuNqd9zQC4KAzPHDSbUeu2C5m/XjoRhszt
Xk1B9KEhvBVhLPEdwimUm4YK4k6OiVHK6KdDp1KgAHLyDTAUyh996exdwgoWqeea
tcJ7tLLHLYje8n1x9dXF4aJFUYYF+nTsd1UD3IcXaU1Dy/NKIGznogVZ+Bgvxgsh
utpnKPcGx1UFJZBwbhH7R9oYx6rOVSqaPVDGsV+ekD3nO9iGbM3zZfYbKPD/hH+9
52p1TsGcnu9bJy/dlF90IeCTkYF2gcWetMbdtbaNZJp3f8Z1Ha7ZLv+6peO7/Rw5
YahEcQbcmDpBaFpWjK/h5FklCL/BDvYcRp0kXkEqY0as7a/nqDYjLSFbI/gzCXNj
+cepTLIgldhhMS85tFGuvXpMR8nvuB8miTs5w2xsogEvY/s9561pHQsqrFVOBw9t
8HOSxaZxBO7k8QDyFKujVLmheJ+FbA+1z6alb+LpDMRf1m6xKAR1NTgh2Isqr4x6
0W+26x+HWc8/Cy0XVHQ/vxInPvdpmdAk9Qq6GzEoS8uDp/Jzd8FOjDGsl3fcn1Xd
87x7K1EpfsUXTCaqu4kt1b9/A+vyqG8zV0EDrJT8paq5duu24WulSHoN9p4/wW2D
oDURc39BNp3cZKu1NsB3bDBSwcxIjyR594mBymgsvcUq649LHALU/WKhkMWiBIyS
CzxfSjNiqANhU1uaOm5eNfP+ttMwQPKOtt3WWKOXohHjxAVhDebu586vaxlzytdS
ylzkyK/ry3HADYCug4QVJ0hSwBuV2/AmYCwCilr1jI+cF+cqQGiez45qMK8G7Ybu
zsQi4OH/6Ril232v4uE2eUgf4RYjPzYO6oSslfvjCXs8bdlJ9xBBf7enfv/o0L9E
+RTWe9q8PTsleZbRzX06FNrtZZ31WpXIiOVjSuohMkXmgzIXrBj2Z7Y8Uouq0XUb
r+Qo+fvYpyujZh9k9/Y+SdCNh/Nn+1ag2LtWpmLWy17qWs/Ql+QJ0hD03k1CO+e0
2jYsDEUoPkEa8sJeXXfBs9k0bdrYnbwMPr0D87YfUDvzWYUCi5awI7+c2L4eeRqj
lwdiI9t2uxZeHFJQxvi6+mlqjkQDKUZqjvV504M2b5IZ7AI8psbbekzsEtfxTvzo
hQkzXYkmFFcR834jZM5wpM5sM0ZTxEE4rAV8UFIionZ6LCtGUrWJcU6Gffz8lhEP
52gXIydNWvm747btJ1ImN6FBMIv+LGG1L+K4wxIaTu/3Q5FtQyivvsecptTsGtQx
lqfmsv5g7CPXz6s+QYjji71kXq3H07BZuEHzJCPty8CTixLJqXkZjqK2VZg7lJei
mRjsc4gb4rxF7X2MbHukcbUsb/WkcgPokBp5hE2jC233p8VmIfHLTl7iFnJSZ18C
x1hWei4hhnZCW6U0f4yX+9WcZ9lf2vp5zeyi9obgpn0rS1OFB4PXzQhmOkxtWDTC
nwt/yuHpWrDSiTzW3InfKUKY8jKbWF5jOudIAVmBx8EWz3Q6On+72WAM9I8kGAoy
kcejNfHucUHmP9MRzzFBcqITNlGwjttp4W99ClyZ8h0cCpAET5pg68SATdc0yzlz
b6/JICIJjLjxuUSdPoQq+r6phQxrkUaPEwjFKQgH9CMdOSMd6SNc6amaG9eRJpEq
mUEbVcRQZi3NH+Hi6QbpgLiKGdtreVhcnC4zuO973btY6BdkyRm1vqrebqAdvoDJ
v/E//DUJRlv1tVvzduWX97w+jdJFHmuUhbaYXKdhFQxqO6yYSZGaGp+XPS4i+AzI
TVl+0102hvlyc04fc0eVk5gvz2+BxAA/Yx3P8qdApSp/pEJC7gv80efKJZqaHo1v
Y6Ws3lytoGNIGHA5YCsZVTTsQf7DAYFdwjcRlxLWctOmgv3c6rLWR2s8YqB2TZn2
XEpYuI99ga/z/dpVrmu2moZ0K5VlKgmxkIvrg4DEgTr/NTbjqyPE4Z2Ar5G2tAtM
3ebLqwkeIc8Vc1zRM3bcHJvhCZckTGhh7R3aWqdSKoNmqftkHAonFGlRqd0IKfkf
ky6Y/keaD5HzGMmNusVFnoVMSz3ntfdxRkibi54xfigI8Vy3gJmV2Lqdjaoz2W5d
u2BLg7RXE9Cx4abRIL+gk9XDbGtsvGHqKB3Kbe4z63EJ18r25X2eY78gCBrqIRUb
U37YOtt6I+dyX0Xv1Io30lC3zDmANZrt/9jAcTuFvzG+U3oqh9jmfNwHSfF/sXly
4YgAB9lCPfpUq1CclZvrjDkevjG77W/TBxeq+2u/n6KH8x9PN735GZRni+hbEycG
O6tqwZkESF6cwdsIeX6rWkv5DPreziVQCvk+JYxcUSJj2D72Z5QH/sh0E1QacI4G
V2psa1YOtRq91iUI3qplJx8LXoplqpoqLRumUVsH1k4yv5/8YJSs36ku93vEDCU2
lgTHE/Ul16NHVqQdmfDZmtFypWTkVxfggEYYAUptGhby/VapADtEeXX4Jk558hvE
eeEGkH4c2TAr1twdQ3gyKj/aFEnzAx8TVsXAOi50VHzJCATTyba6GErbYDI09DkN
hmMn3VRiaYWO9JTRYbaY1TW8A+5+0czsYF8nOReoa+mhHjqzFuRknQfvtCzVb/xC
V5ld+vur4V1hGL0FbVZFbaXTssCGB3yi12afc1PbzVn+VJRLDNujAjsvsYdUoXfT
5TM5sMWIbyKdDQ8RFCldh545u+mCqWCLjrQZuJ3CZqoJlpnWrUHuNqmQ1mcuzAY2
BoinpKkIm4FzF9IbidtTmrjWs09k4UjT7wRLfyqD+tpbbqgwQqYhW7fmLm+tNam/
PYUCl4QaMXJlE51o+ls2vL1ax2K4SNKHhzqJ2iB4MOcHOrSt70cTj3D1KrHpeX9I
Zbejn10rVi4Oj4HrHL8SKB2TXvZD6V7CdosHCjpV6rPLihy10IevSMUKUjXNdHJ6
cZ8xYkElAHMMy49B6Lb0Vdhp+gW7+WNUFi+zPJr8rcFD/CM/DsIqFTUO3FqbLLOt
ISejVAh0B+74EnnuvQskYotK5CJdECa1Gd2VfEyzfI8I6/lyVkTjsscE1CCdy3Zq
HXFqJFfLVgSZeq5h+trcvf3MbxVk/eZnuKslMuDsBj/KQhIA/BFUVdISHdVadXY5
4VuGz7KhhS/VmzcATTxIOQaIVFZEFX1HFmtAzwJ8GLhdPkdiJZA32i7wb/Y0YNBW
0BlN+l6KKJ6BtOLqvWZnqa5+KO1UzUACa1Pg7rXL11KvkByvePP92sOVRa8LxW8i
+RA39E64OFAK7ujzs/jIMm/UKOIc4my9grV4/4KqxNzvYMlN2NlWgzp6dMZFy+bO
pCfqC1v8AAmopxkIb+958Qt+F0krwAK91goabmYHDRABRC8Pn7nADGnzXQw/Tn9i
yiekvAOLcyHMIWxctD/PlhH8X8ZePnsri1gRBE/6Dr0edD7+mEZHgalrtk9nqyY9
yMbffVoSJ/r1S+SOkZT36Rj+ZDyhkHWXwBjqBCP3pwFw+2xQJZrzDUbJv+TpVdSY
DDMhJB+BnoaWcRGBjrqnBh/7YsrHZR0mv8VHH3yEz8fVU2X9Szdv7pK8rTfKqvR+
6yWaFY1/Un6wNvK5NzG7QM7a7OtWJQ/hHwKxwJpAb1kvFt0Pt5UFiTOdptqisN/9
dAfmDdYhq+Zly2XnNK+QYHyPdp56XDQj58VD2mTaApnMSAzkBH/BqIxS84OmsgbP
UPpox6ZVQnAuRnq5bGREQ9NyJvH7jAS+Ds/o5dStVfgeMorg6qK7vDjlnyCiqe4Q
dIocHaoRhIy1k7T0S+N3+gqfaXDzsiO/4b6WQwYGyXOaoOM/6lrGl15SWRpVBXfr
GcDzxFJmsx9k+BY4CTBrkoVow3eP+4BtXQy+M9t3lldPFycds/pFr9/xkLx0X2ml
Pfm9pItJa/ZXIkziVntuFp5gPRQB5aPZ0h/PS3JPDa/3oNDL68Z/tJvt1thvpNqN
O/FW8gttFnWvYGBTcv2+VwFoUDzdepaN46jgyyCC9Xc2nDq60vA8HPyrhKzNFExo
IQun+esYLve28tC6XlX3nQT9eEX6bKAaWGO80ny4kLQxJEDyEKAUeKlnkTpfXEHq
Bfb+sHFajvScVbiUeYW/3DyG0A8YkbtqFGPIY3YFK7BFASSEU9IGz6CWPDv8Fc57
MDSB5U4jbTZ9hkHqkPJshWznxwjlD/c01bcdre7DpEr6N2jbS3kQl6sxAss5XjZb
OZFyKKGPW+fFu4jdcktBHWEXAumxY2cBFpswa+TElv89JBYBttW6Xh/gQZFjRFMV
Qp/ohPVyqIoG7rUzahX3XDH3FViNGG+o+1ZKjPmrQPF3vMovCv+GeeHYuwfMRmKT
L6PwUysbBhQE8lfbzox1Eq5/FYCOCjAfmRaPcnbh2wP7dQKTNSnhgV4x+EciqWT4
gU1QiM7RviA9UmqaUtoIXqRqO9V0u+2oapJifIJaITFqHAbXDbk8/SGHy9wSCE7u
/lAgryN5hMZDSkhiTpeJMMJsfR/AYvQBZReyT7Ibtjp9/BW3EJ4RYNuXqgZtbkCG
U448CnK0QIjyIR5OhI/K+8kdNyfwJtAvO+oalTrrZAwCeqKymOFWrogGaaO4g2Gw
01SSwzZUUh8Exv4UlZzWS2myvKNfabudmz19NGrqeHCKwH3PWCY7pXqi0QaD6Ljk
l3m4dOvyC1gouzi0+D7T0D5gx1oWBqYju8mGVbmty3QzZLz1HAO47zhOC6utBfDR
YErZ0iWTiRNNhnl6UEDCtHA0TforH6ErSHGNCGRKtpKctmB6XRL86SmM9JGXtxZx
Z+HaG4JN7XPVvqMCp1fKa5/shy4f9JXSuMctor/gStO406SS888Dv/tOOfZGrDQP
YFeO+xcFYtyBE1cLQwsHT7NEOgBM2Xn8rg1fXBQC4Pa9rDwQiBo5mLP3prraYoiU
nOroBjboH7+aE9JHqhGVliMMMicJHi8iW7YuLCxEhTksjQlYYgJBiINm3nPCAXfK
hFE1sBRR+lFvEzgUBVwLrWgJ0tMH0beS2JRsWmM5KJIu/OfSkh+G8AQBVFYnfIeS
pElM+6aQz98ZYtvGDvsmq9Ozc4j6mV3szzSo6JGD4vJ9f84ezKE26iiJmIDLVVoR
ByowRKZYmx//DWNhxz6EnjrsCxU2PCUaPOIwEOX+4u7VHVbJjO45ye/hapFHjHqI
lea4/LaQt2BtWDKu94OYowzO8HlnyOWSqMn4wZoPpoZsufhQPVo9u7naJ1X21a9a
RcLHGe02J34lGi25c5/1B0Q/5HKUQRIqVPC1AgP44gjZJEHQWzVFXT3jrHpoACea
xQBXN1eJyDc08urnS8oGoADGNTB8mqMDOCfl9E4FF4ZHmGICXyW6Eq2zRHLRSQ/T
5k6VzHB9SYgXNdMpQmgS6VFMmoWFSHp4+frWhliNO42JsJQEugg5amjDlRgawVIX
dXsOm8osg1o4e28hXygAlm1BetCsRb1t++WC5OzU3eQ5umvHwCzuFfCr9z/XS3rt
N2GUgPKhzulCD4vI11X5sxZbN1RmEvUJk37vT3nB8tKznzmizdth1kPd5gf9Z/Bc
aePOyuuBqmU7U5URRpNBe3w3/N/ZDrk+h0djSwicDIfxQaTpo8xd8Ydcq6yXQk9z
eXGj6Z8EWm/EVk32nxKC22T+bKv1+U0YFvR1AnsQk/SBxNS2DkxvcAiELinIF6UA
Ffrmzt7YTOaDNI+1VeoPjhNzRCtLA2c7Zm+XdDiu8gXYtX97FzKf48xkvyqRubyL
/Iwn3DPxeB/8LVk+Dn1MhV1Yyl3FIdIAoRA3Cfs2sBVh+I7f/M53dpdJlIRhQ5I+
9TScwPZ3HsRj1eiPBflpBY5GrVNKH8fI6mNN7RrtHE8YDOWlazjV7qtEcFXXXstI
uq+q05GSsd3wTVH8PGLHLj+g4PYVVDwcaxcF44omPYNrgyKC7GadvbeuDeNfY7bU
gljQNni3zDbg4PhSpw9NG8CtjJa89lux3l7MinpxhJDAs6/It/mz0e8fszDxB/tX
D6RrRZ0e/a3gD+z1PZnnA6cyQNtd8Q7b/MxqCC5q/EVxiPRQAgLSOhS5J3dgoLN2
u5zHCYE0VJRgKbAYvej8ulxHgAkwV4c6EmoIzfePJTCHLeTRuOsGciisCYb8ggRS
WsIipeSONTBIdSK/qdH0RXf/B/xZ1kVwh3Kad6ItseiO/3wKCreTWI8PUWyCfhNR
z/uTYxzMDOTkNsGYbJw3a6WCMNEjaDcAte4xLl/FxuyMQNyWUuGtuYoJBxFEM6NF
qZjbfThmPdpd9ZlvNO3nhy7nccQR8mdsNzCi6CHsinqDUT++vo+GjIULm7jSsICM
xfWziu54SVeEC2gCRvzDk6bwhxE2gAjdICMB0zHh+swsGHHe4zeirfCT9b1fdTbU
JpEvItp9D0By8khEtrZS5dnls9wagsM7bEail0IoSdI8XakGFO0XGD4juwN2H082
1EiJ8Kg0H+klIsarYI0l5NBBUXf8hYaLl/E39FWXq4fKnjdeu9ZXlr+TcgaMZFrG
blPKQG2v4NLxwcS76zXMkiB5ErFqTK4YAMSSDPG5UH4qqmTMMA+ODk87c6a1dpMH
7FeQiMNSbUCR773skoNDww0NFNyEE2vteZjfePM1MbBao01K0L31PbHQR26okR9s
RIKM5gXR/XE+QVy9IrB1fbdNmGzoY2LcME+8K9zoV3mvaYLwSw6DT1u3MD+ajGVr
Jox3v2LCd0NWB9Sfr+s/YnJQzteKw4rwiZCcD1gZuCE7/QbXsYR129CaOUXO6pzu
7EiKwrlCH+CcyTULbBPTjhUFsNizWFrqxVkeO2Ud+jLpIvmSlR+EHhTgqRkWoPMs
OzNc6lr+n4bUoTLWc0RVFuenuUutaRlRyC4tMgsxYEDPBheLWok5nflpubCuSVqh
L9/jngyynX3QHQV084+HXkWQcl2rO6aLAH2gZKeScCQ5gs961+LbJTKR5KgjGJ8y
I7nBdYpd+SPzm8eiQlQgVTq60YB59ypmWVqOuWR9x5Y8HjGAc5CBn1cS5cXyNcjr
p6tJ1GsDkuxdrM3PAVOfFNwqSFR1Uuzw/uzdF/yf2nujGNj/tlwglRlbjVtd6ySe
3TkIZEikYLKxpAkjO4Hib1MUMKEQPfswglzSvEdMtBktu2q6DJrLlDTsOGFmILyK
CHt8H850YdO0QG6PhlukBfqo/cfdrWKFs7QBk5mG4RfRJUzlnSok8sfQl9yHFjKz
cxjXITQG9X8A2yqgALa0Xx6jdl1QeZV1+N+j+Mat08FKkW/Tc9L1pxKXkOnteSDV
GLrT/mpCfT7gMh3RoL0XHuNqvuMwLBKs2Fx5mc4FHXmi39ECd/LDPqjYM2PRkiiO
TxFG+Nn002Jt2YFdmIlk73Al8L/G0G6AzLP75r35r/yTOKZeLQc7obgVhQ2kTXJc
otpUG/hKbU5JVarLA2lvoXt5Yrij8ABEDWYMFscT8udydf4q+BAH2Hb9WREIwwvH
y5qlEkvrWndrNMJ2I2o5YmEBEqFNGD97VJfwJajVk3J1KKtwb4HQmZIB9T63A6/D
aAKdWTWcEJBmxr28FFvNiRtDGj+Um/RNotiA6pnPHD9PskiWRCx6993ulQtPzEdQ
GG8mGpLvxB3I4Us01fwFW8oc0KtJGx8q+LmSUN27IuJrIFq9XPq6ztugPm++2rtC
Xdgb0yoDlrl8FHBZ8wznPnUbdj3ST9ihwocBzgF1Siziy8C8UZP5c91G3qa015fb
QlYlNMrDyuUjAH4rE6lornKNOAalZGo0M6jCmJXeAnHAkmPykk40gGltFlcOmJxW
n949Pytsw2jtRxPi1N8ZxiEcKLNHbBFn5InKhPf5v1IfaFAgyVRj+2g2QQUaP64b
HcvYajlP/e03DWh5rZvwUjWcOdAxB0n/SpJBZR16K8G4564Ctvrd1Sbo2ggwrxb2
2kDnhxLbi2UyepjYXRfxpdwZWkALfse/tJSUZiAKlcEUJMv/RFfu7/E2Abp3u5vz
smBGKVJZ5AiPzhpH1Gmvt8/VH7DVnR0+CtocWfnaOfBO6VwQ+dRqKdItT0hmIja7
Rha+XUwxerLKBB3wOpy1uLJJMJ5UNqTECoJjsUWTI1K5OYTcIVbGNamNZTXNnPl+
5Z6NXzB4zDX9zUpQcK9T+rkq2Naifzf/eai8g/yet43KDyleP+YWl0bvLJAEkXqE
nJ+AgpV2B0mX75t+3fdDPDok9yPqQd7ivOWRIUZxhb5Y28QpLncsq9JL//aXeiYH
vI7z6mz1/4p3yOxOn08sSkykaUmkMsKv6sryxNrEcx228vH6p2iUz+S1F7x+gCMV
IYKjKvqvHjy11fDq2AYSu82oQtoS6E+Na7EP5rIVuOTCFDULPJP2h60HQSe6lhNE
7Ih7DLxdjPjPXLsLVlyfw9nju8eugRRoyn8ootmhGkouyHU6X+2bk513IuvQ7hdL
Iug+uIrvDuzIQbko8C3eIUW7zFgn1P8RtPZWHHb70RSva9SqMxmHx2ysd0ixvv2D
rndxN0mtFT7jViZtYLZPMkFM8aED3ZH8hEpnFaOQxACMDKpU8fzrKsjvq8nUQOUz
6InDk3TAhPYBrbQ/h3QoXKE2NyFEpj4MD3MUltRPJ/VdjmOkUX49biVJTG3U3m9A
wOSZU0gK7FVsX0uq+FCBbEOUmMunkGmsJ0lahmzGsKr7QlBsZCZMDdpMyaQi7o6b
rc3nNVRBxovUu+eoQYFQpDhFE2XTwgalWs2EmVuvwtC8YHeEa4B12wC7d3Gnay3a
TQd88ucodmi2x3/BMoD8bP3gnwvQGLrUgXb4k+uY9By/wGkpHy6vcazHHppQtI/U
A+7k0k9v23E1N19/8yvtECYKy0yAZ4JUzdSP9Zx8fEhMR13eEOlwkuKNCD6Lzw7Q
UTZn9BnyUprwc3n/p2R7eV5ZAVMWNAt2Y0uRgLezckpwdDanOWho1bRhPRSS04kc
/Rz3UwODQffRZeM7FN+sp9xx1nJG9MH6Xx7X09XCNNdCSZ7g22oQJCpB3c6lz1tT
iOD/OOiGe67DzDElURCsV7N+MDjgPyPIwmQ/ydEPDHpiuMDUMRVwdTTwbg9S+5l0
3/CrYPonR+AEqn9Ei8AG06o6tYUfHukTtcCofEJLlv/gDjGY+39FKhshlNCOHlQ/
isCxHZpEYLIVB474CZ2VYv06aT6fhby5w3vnf7XoGGodz0An6ctr+g9PosWwgLtz
1CqIVRwr2ZzPax0Mv9eyOjG3BsFVsApZ45YtgCPtcDJXvX2cSk3uMF4ZbvIkbnaY
Q/hRKPL5qprsom0aC1t2IflxVSxLB84wcFh1PsUCx0TjH/RX+bsq/St7nCCC+4Np
XFJo/AFCcmjsG7LyMy/oISnPkaFeLOi4cDIkv528WISQ2VrhCYvxfbYPbqN/pfMR
aFnXpi0A4zYdpCZXqBkFG8MYDErx8snsIa+p7j9NT18pgr0IqcvY6d2d68C8BSg9
gPSPQuiJzpDtVDVryavl2dzQxctUn44XuBbAkQd9PAxnXH8xSdR5Cc+n7c7/Iop7
9YZPVPgWgQ5GquZnotDsHGcwRSVAJWxs3D1AtMYPW9L6aeilaQypafuii2a8aBhB
incrhH7UHO6yic7Jp+41e64/5C5XVsi7kW/LzPYJzuVEPYsh28JR3T9rM9NUzGa6
yY5oNBCNECx8kaLBEP9P+lNnXgJCfgT8kIeVN1RdO5TfBxvEfkKn2acndP/TmqAh
Yv8MyB3iHwneu4jq/752PN9t9ERhZ/n84h1VHMQbkpxjF7sC3uO5VHlJeJOZKWfe
w0j5cXuPVL5i/6/XWnwAFc0tBLozzAp42wGp6EAe7VvuNPBgJLEqSQBukFdEaGZO
kFG1vnQB4CfXFT9ruJPtWyKNUUIRQCPPg/E3BCs1xATKRa+4/jahH0PK+e2NL+xV
YclbyB3OPw/ZqNTy9A+Pk9y0E4lHNv2HzTTgTAoowZwNQU8IfROb3lOszhVRU20K
SRT8Tkk45jReDTtC8GMI1QEmVpjCVBeg9EoMAzLQ266dK0NZ7SA/F7m831d9RQet
Wdcndiq61H5Ugo+n0+KZkBXHMKbrJP8KuNfGY0LuUGdMrdSUtG17OC0ZNzqz5mdt
MsD58XNDsH8ls+4biJ5njPcvCRRypROH+NdeFTKBNVw9/HkENQ6oAkXAChLtgXmN
epO7Nwh2zLLCI/8aoQaoe9GgafHH3U0rp3lehGhn7AbdwrtdTGHDBn1YL1r7/e50
V1aWpebdjPXSMrJB94zM5Y41T/2i1fZ2+fKKdpRu2SyOI0+WYPY1WSGg6xLUBS/d
e16xFs078T1alhkX2Yf+BDyNzGPKCdoTyDWpUgRXyVr/K8QFD2gFbMtPMBTHL/Qk
PK+5kpm52K/TyEQsuheqjQbT3+Xhk0+ewiXlV6hG0kRdAtwUSXViNS7tozQH+EE3
1I126Q3hd8jPEIfoaAhzn0Csi0Iru9H2IMYfUeF7Mw+9R9ZYu74pfcZwFEA7yRjS
QRzHn3JVxckoA0DQhFSDFSZmwrsqbNmJvsENHHNFkaPBrjmdwsGkgnQJbEroKwpR
ipHxSyU5/+zyDvzzOm4KMc0hAZDdf0Dj+uF8ovO+aBXYz3sl5MS5sJRsBq0qJKbB
IY1g87EumAUrAti/1Fr7ZXFz7AryG4Tb1JkBICKzidi3UzTATqw+q/J5HVXFm3IU
bdWXIMbd1QvYG1znX7PcoJKtcBzc2TNOv/kHdY4x9pVan9xxlweOJQWaSjClQUDQ
hgp8LmhGL3SzdYvf3FV/AIRtFEE3U+tWe0AJCEVhrFwC/QqVnm6RGQCedp0lAZVv
RgVGF37lbK3GOmj+bE/KepWVLHu22uUkBrYbGxYD2bug5VQpEpk9WUbXK8BxTftM
FKp3ywxnUDLc/5QOxd55+I/8T75nbuODuwpeB5H6nNBj6reSlNDWAhBds7ApZ2vH
noNyrGT7n36DUmsfqh9WdgS4mu063Ku7tv14ybthfK2C8YNrF9v4+o9Kj48xko8H
pEtyCCV7TGCRMD9U8QcbPat6PzIK31bqixEN6yvun2s7ZxrhQ7BzCUAaG0XG5Wyj
tOvKY9+DIr5Ggiya+v1pQAyLy6neKHszI5S2R7eCUOVDIydGMwjbnk6DY3eL/1xZ
NAOYrD5sdKO35h8ZWZ2h6uANdA/k8nlf7Vjx5HVQPj7AJyQzAiZ6LcqweCiTLmwJ
Joofe+rXJFxm6ObD405AP3Jhg8OyJgN32qlXzTJQewBcQTMKhVPpUiOePupuJpGi
28u1mQx+zzXM69lRRKAO2F1pdCHOB4zKJG1GT52pRdk5pEDI67le8sjxHaMQmTuH
sTk4QIxRglyz4/z90489/AcIg8t8SWJ4fGi80/Zii3cnUo/AIcImWRYd1PbeMEDN
ed8YfGDxLyPdQiGzB/jPeYSsNls0skThbCCLkLOXRB3Re6C8r/JMtFyesp13hlVj
U4vPFHJne+0M1lbrVgVrVk6bw9lLSI2ekmhaMmkEwufZOEZkZ0nbLMeipHIMQ7Qa
MdYaJl5p7kfTkpQBr71iO//wC3CXfBSNU8MJLbURqh3GskLE8DFLnFHzHm6XcwJQ
omUcr+nRzzfnHqTNywBpr3zw9x2iY8iuGsGjQHwDWtC5YX0TLTvnSPk8kIbzKIFK
lYJbqem9d0lqq2ZtB3UaalneW8c3t7vbauYzh7oRvKFYOWz9XPhJ/1niqamLNZYF
1KUJUXISAsztQKXPDrt4mCiMD5aZBiM00N5sdagi9rMIYz0YSDKtB5nERQHgc+6f
htwqYtv6MoV6rk4SP4kHJXsXfDxnzZEqY04caXqx+zH6EnSu+0yLUw55uVN0cvrb
JJljmLbRWTiy1CncezDJo5ciiYUfzOGiRqtyHXPyKy/o++9XzIjr1yjsMOG0ZiXX
ve8F3zUD40T4vnsIK8+fvgEiTEMa8ZzlPcfPNE0B8AYx5clFH3fiWTabFXn3miZQ
0LAJJGZgBENTjDn8w5CG2WJV8ZfSoovDnCye+tM6Fvf1+lNV+Ca33sn8Oo8YLJgI
JvSPBaGh7coTNV6Z/n+VbLwY3Em9yaYtptv3BJhlDpEzZTuckWZUq1NzI/80xnl5
4SEKMOKAw389Dd2ZzwUNFj/+L1xxI27U7M+fbvorSkKAeQRsgzasMttd5UW3Tnmk
d3tkmqbvPSgZvTsZ+6t82WWdXGQ/YGA1Be1AMruaL9Fu6Qz9WoHOQhE757+m1hRw
VxIaUQS6G380SrD7QEjkBDD2SGXK/o4zXxBpywuadNO4xk+8tTi1OjqMyMhak/9i
TKpdV0bWVXZenVuNqISkmSe9No970GADL1LN1shpRb44CmL1wXlxOAPYnLsTWe8a
miLCps2kV730gI5k0b/M7T05beeL1qeWmvqOxLj+Pi9RUDuuHfRrDb6vcPOHQkwg
7MwawPFYt8StjV9U7ScYCkUVGAge62/mej4U4xMwKU7ybgGIHCuuYJsjcEaKcSLa
w4LhIAixWeZhxO6uTVdoQRHn4smvWpTl949fF6bfQkZiduI2TFQqXLytqKRkWwVn
3rVgT3342iU/sOQIS4u7YbwZqiNFy6rW1Ubervpq2AMoLEFYJqBaXH/deWZYfTfa
8MhRGLuY8BC34BiPCkByt77mt6+/cbKaN258prumv7RGPKkDMt8x9273Izxnwyj8
JSw5taTYeUbm20+m5lRIXRlIZgY6orFWPfaJiumj8DnNm9mirVVqsHhSAtSyXTmD
2AMMC2wPUqsKcPR8J19y4ftz6qQ+O1VmJBR0WskdrZKtFm2aykplBjSVSZv+mYst
SZD6KS1O0qZVL82ofh4MErvSlrCHhoMF4qW+nOtmb0Ukwc4TbnNscy+PiG/exOlI
pPBWi2se4qJX3RY4FREpzKQfGoP2UbB/F0FEUho8M/FPuz6g1XNrv3224b2qJpbL
y51PTemXvjvtMYI1MyEOHN4vxgUaELifyzOlQrwrC8+/OQoDQAq0ZJHScYnLYeLi
a8wN9EIGHv/yjWUBz7TGmbc/h5c/JN5fPwQ/nCWQmrJhGaxZWXxKU5VNYWoQVL5R
yYENkJt03hurYxiL10Pe0TVOv1631m1rZkDDtieTxQ6+e1LGX6Q9gXvkwaMT0YSr
PBBmDlncvcC1VXWIV/k/CWSUKhhT495Jeoi3Pf+TJKBEyvoZYZgdd3rZU76jIetU
zMHLYwq2mNytdTvUfd1vvzI+qNqFmtsrF5T0sDA01h1wDLSkgB4OvHzNA9tS5Ct3
F4fBAU3BuQSafRJmBz96V6zybILSR7gFoQ/KZxbTmNmZgQ96agFQKgPOIG3VwBqE
ytB1WkekDL6aPJCpbOZRlR6p0BxjyFqYHDjOgdzxglAy6Wtv1FIdoqQcFj7m6+ib
Pr0+c0HopxbZh3A3lu/MUYms+siH/NOK3VrmWWsSRrj5yaZ0rS8ljPOeIjjjjlHU
cOIheN9p1uDFAOBZdWPXUG0Gv9NA58CDQqFnH/tcck9H4NjJlRZdfRjj4Mp834xy
5XEVxdBxtDWlWOL8N973J8ZLfKwvbY1trTVDhx3YPShOa1m06HqIicLMmLM+5zz4
f929DqwNDH189OF54XoGVFb8/znOWnS2BKu3yEPl4zWMau31l0qJg+X683B8apQN
LbGXF1DfFtrOU+SC2XcZoIt7t0oC5uATr0ENPHzu/JCmqS3iae38quqc6OkOi+Qt
uPUyS2Anxk4KRnj93k5HZm6WtQ9QyELylbUBmOlMCH3D1V4lXKseiqN1VJlJ32SM
e4jaDFh+Rid/76sAdf/jpg943rDTJlABk5Vo3TAHCwH9Vx8vIHqhIKlCQlzHe10x
EPAgZATItigVFflxdhlGRxh96Qjf8YiQzSCX6EpTbPTxURK0GxbnRLDrjQM3ZqiN
2urcGlBV1cta3iy4NDFDr6LcofQDKaI/QfwXuJFO7vktqoBQ6b9PKjUUFVa091rW
3Ex95uzkSUdIlB5NwzOBOELoj8YpUkyuzR6HHtmCD2zUGwF6PMXy/WoASDzYCqXQ
+2cBpjHdcRVJE5w71kX2CU87OhSxcsOiaTQQFlEbMxrBuPxfl3aC800bnS3t1zsE
2vH+rkPZpP8ggjNnUERlH3MaeZc4yAj59BrObqEHLU+HOJ/ZHCJBQtIu5KWRgqBG
3k1D+1y/+3/cfXZ+mVwJwdW618TZGFCX0gDDEr0dHCgA2eM7Ma9KYBYIkxeZdBIC
42SPCNWqrK72eEUF8CKUTjy0CTxcl6uF2MWm49jTLJ59veFaQmisUxsiRU2tWUM/
2zzBoMppp3x4r+ybtEEW1nrjni+4MRbJOr1+6ZRnHTGmP2yFqEoazL1aWJvPwwwK
kH/MX9UXqwO6pwJnSF0ffRxf1WpKP+GUW24wUISFi83RluRd0H4LyY+3a7nYEOG8
OT6zQJfqcwRdN0go4wnKz3M+/gUo2e1WCnA5jMLT9JNnK48VaAEAZNFKIDgSAPYh
/qo2DtrsV3x4muUAp9aFZkr/i77IIkieFITWnCnr7GtLiI4ok5Z16qA5p8KWTpv3
kjEW0SAvh/xvOhIeQ9IqSXkZAgPJ2XTpCGHot1pYgvYZY6z4O0NCN8qKc38TKV79
G/Di7qzNIG1k6QzFyzmm43SICZ9gjnOfhp1Gvo/v7xfi/1CpXrqWzFhgla4IfKWL
8n6xkLlHxgucqXJBZ0WgMvKf8DXitGSiXzIrmZAzo/iCV6y51Fv2/0xI34QuHKJx
Q/Tz5U+BchcCU5bmnfPwtqIQP4DwNorAGuCby4mYDEnT0W5kfsRQd2nnpRwcSa5H
Y5mJJuTTzbmloKoKUUe10JlX63b1I99rZ4mUUTnNoiISVNKisJs92O0RGCoWhhTz
nORfVX/q/EyQLKKdwsTZCD0bI8bqJ6iPpIx300AGRscYLcV4kv54u5z/e/EcNWeG
KIzkZqZX0+ZY3g9XC6Mm/UM1LLa490MaRvE3BX7Jf5dI9ugiZp5aJ6kXe+GjSCrH
fUzbU9vfQSeZ+XV+r7ZQ6xkkGj1UHOPfsdGCRTJS8bmSq4jdOc4+Z2Rp86n4bAZV
zH2kNWoyIhdvmUGVKgz9CeqSPr08sWfMlKtU+O6hTF5VH50pcMODzQtyJHRNTFFa
57i6T5eduihgSO7q3bU4Lz2YgBXD4MsWPIyGcq/paak6vQpptkEQF9Qrvob+C5Gf
+xAtan2rvM+GLVA2dYF5R2LONVGHDTowewynAx9Fr9dBUjRlfNuMuWFxnf6DjSRP
/UcwXaPPBHgjxMOFqI1HCXsmlj9Ceo3TEqfTZ0t0x+R1w8cYR/LrBraYxWyKC0Wo
2OokC0L7XplFAs+u4EOWeHvIvqJdDVOPf31JhqICmN6CiJYZTymJHj9yKoFwNB4A
I9YUS/N/9kkLZ8+iJIKlIrcp5amYD+hOhUdcWfp+5CevZH1kKL0sk0mcry8/dTXk
p1Nq3WQ/L1tz+bxzVHPiHcEmFoHjiNyFAUyhoTNjnuw8UZ9184mWWgkUYS18BoL/
+gxXN+YgkdPaFk3TEx4sjX60X3xy7DcAI7Qjm3OCqaslvM5sjeeOpqF0oBlTxGfQ
lhhIunDzr0x4a7qWhsvrU92qZi80RvyR/G59PKSaGKlP/382wwYj8dnyQ20ObZ5E
sJWfPGKDj8JmJZnvnyWTrgri4tcfrupNiRBb4+i9864sL1szwXkExmiQA5/ZIcuf
EimxED6d8uHRhFEM5zlYlSFrJz46tS7kwtNB4BdkNIWvFH8WueM2scUTxBKfpgmc
mvhnH7LXwGCor6tCDWlOLJpr5UsF/Lkjsatoz7Cqpj5G3c7bE5tbUxMjtdaFt7Cw
Sv8fptZtrePeh0P2jStGT9Q91IIVWhl/AAMHWC4JWqjZb25MHrtihyN9jstB8shN
ZB/A4PjRIM7Hp/vUkWBg/D3749eH588iUGmyHTcJNLxzWQLYWbkyCT0SLnD38rxR
tZkORneCOKB+N6a2p/XovCmEzcc7dpqBCD6F/Q7rUMnTWSg6OvWXQohBVVm0JIpX
eABiebLwPAmUmn7GWKF2A2iLTgH3Qk7Kal3wVT2E3pGHlSyOKrD3U9KZzg5/EvSD
+ZhML50fEt/PjaNSXTGYMKwCwpDcZSBP93zUdIufiU6ACXFWTZjeUSBoXDIblMU2
cQmyvBWPKsIgMWOC13F9U2qL9uv55Ia2RwMORxBkzdK+XvNHDBM0s0pU98M2zVYR
uzaWQ7+linNuSYO86gybGZouJpNvxoKpqDWvuAWbGX6ioe4ns8GkyiOeyiNLVW+R
FIKs3yecmjO7BVoZhWvDC1gOo7jydHxZs1u8TtnlhAI6BOx/Q7ZT8Y5rDIDRAvw9
MC8IApFB3QdYQKmkSj1XB8+MVtAgN00bPj8CgRxLF/UUcHXQSzAm1tl1+pwutnjw
fXW5ZqrhWviIYf4Ebz62FbUFugbwhUDgdoa7c/Xbu0Vm6PBclmK3/XrcjIBxR61X
+BUJLpN5IQv0CvjPC3U6fUq1sI85HUpOiDezDklvm2OU2QR5MH/ThXR4k6wduyyt
ue4gJ/hFjksAWTjpbNXVT14uixIn6hRZ8UNB/n3eAjpv+snkn9lRiCjVQbavfw5e
2F39Su6GgxgO6SY5kvYNk/rGw7xWmO4ickFFIj1GB86/+yiMbek5rjOA+uwjcFiC
6gI6+oq0qZPOfitH+nfGajW+NQR+Myb+QBFjtiA8D8ISaZvVKLbakolpT8P13Ble
KqRu8BgKrZ0BAb9ukLh0H7zU8DKLuknkUXq4W8JnzDfqvIKPgADLlHm72upE7RP9
LRvtSeppbPnm5p48ez4Dw3TTKnrxwKYi9e+aF0GDxYv4+mYbaedDgEje8YTqJLoa
bfT+wt/1C4RXzoOaCWSyGTEaydMelkfGUOh7bBdkXBlzB6wB6NVZALwEbdHPctLT
Eo3+YxixSkJSRO6rSa3NhgsXujPQgSPa1g4uaZB5anFFdmldZLE6djs9ncp51eWZ
iEEBR//m2MXQkcEjUHtdz4z1K7sx1/bwb5VumAhjdJuTFO0hNOfPF0MY4pC6oHLi
mDieJ7N6tb9wOmspQAeuszR3ZZ/1r7euIl//hSTOJ3wKtE6FanZF6SXKcFqwywPp
nP553H98BuNWcRAk/0oX01haAte+u02GXZC56iNxd7X3Ds3kyHqhH794ZNJjOBtg
WqX+1PPsrJhemRlLbol+hSmJ1qvZvHfuxrWFiacFz3rPV7LVUQ8AHoC02gACNJUq
4P7ePv5WmNwu1GGIpG8vVLkVMK1xYZbWoRQfJk/jpkHTkhVRghRUa+x1+mO1Po1P
5HPyOP57nt6P7zYHQS9va60wPo4Gg+sjB5VR7zujla8/BvP9WZeT7IfNTfHS36aq
EG2bamDk3vMRB1lZgfK0m2jluA3lm0aopywhjKRmvf+aCpX4aZQfOmRajqiIoKfy
CrajFmykCYQRaHyrKK96HFebFFW1lwe6LYHua6CvHTQEj2EeLA6dwEGcRXXQyeSV
rSZuCD8mq2s5+BD2D+jeoHc+8Q3958glkoAE8AUQerDito6ARkJ+GQDrpW9xWtWm
cTy/mhrHmjTbmkkyxRwSs+1l7blqW1whhO5ncHhuJnjoLrQ+yx0lcr1/TxDKZi1f
oDgUF1ydOB8pWgXfW9KUzyakghgwos5NrYEO/JpjEeabGErY+2sl9KVVnItFQ3YQ
J9+suhJYsQ0dYpOemasbvjvD9QP4fYnuWNTAfhR8AvfNHwTghvmO3hRQkmJNA6vd
VmgGLyMabN2qgkU9eATt3oXl/Zpp6a6VAW0ceDSHaRV7ORDy8JhyixY8BuUJGaPO
kEsa8g4QhKa3nXF5quGAkjoZeJqUuP5LEQSsIIEKbbf/s3WNVQx14s2IwUhcwtTR
roy1TR1sN6jvqeeOzrsBx/vPGiZvS6ZZZkPhM673uzeV9fpp7REcIvU23dt59XNB
E5yBg2+XqRtKGfNGwDTiNh163WfZiOj/077ai8IdhSr1ep2zoyIR8wDejaAQYDkw
GCKBjoMgXSTuawBLKX64BJsdeU5rPPRFyYdPY491clTdCXlF4/fpJrHstyc3NQEq
JipYLaQ0ibM540HrpGWkUj3lgtLihZQRnyfHCroYDECU2lqFduocrbvcs9+D17n2
WlOduTUMW6bZtsZj9jmdswatExhrl1eTeifI34OXGg1KbDwMIW/eo7t5RjncNsfO
/6mhVXkHZeU6NEEjE54sVtOQUrkzJltGd49orz3DAOiMxvZK/H4v0gATmpkDibhd
qzH9N9dzm+PMtDdIF+2Ktg/OGdqfDZLXHSiNHXmaKOaQmV88YPgQKX5UWZxgifsK
y5H9dZ24bZd4eZUhlzlnK6DG5Hnc5fvhgWVR3VJMcK81r22kSntO8CtuLDTA2NbV
OxRf7K9G+xyHetH9M2pqDPkr7eBDLZeQY/0/NxwDv4Nt6r5uACZku5+6wAtKQgjO
egrkPxpf8ynyJPl2dOVMbddGPXU8PSXpapw4bV0ZeC82VKoZ+f4M0xa6ibRtzvJy
39VvZ+z18E4UXjoVwPuMbX7lq5JNdHhMq92xPLv2ynI8sL4DQFY9DM/P2Dg5D6JF
6Vvv9PGh7WYVmWd074bx6ZWNBMqefZCXMmPOKkc6XHDgyyaoxuWBKzEbC86Lnbz0
q7mqFLURRjzrlcdwnvaOJolTT4KT0IBqMbB+97iPdapeGZki8aCJAHqSGwmfIxU7
zeO7uY9h2OhH7ov+411i0KdEhN8KHwJv/TXH3rWhksf8hywcT6Zm6R61hEFkaPvb
LyfkXq5WNf/I+rJw7L+UHKNSn9NJk2lrKQCHWhsE4Enuc3SfPz3KGQpvEhYVC0Jg
9hEoLjRej+Arx2+tWjOvUUHRfbnoLahTV2tqWcOG7Pv+j2G32uY/ZBE640kMpUr0
fUXu+R/ezZ0j+YWmRrApA81B/ItXhaPIV12rZz/05I9T6x+7FlILeh3xahKzPGmV
XXBTs9ZCSSCsuRBrNs6r7VCuGe+SfbRHnGHLSx2yeP9Dpcyn0G9daeunOl9dxbOF
l/CysBtAznpwmvoNeVxuZyhKelNwTMczM4LGKwrhK8+oaPVvigz0Xp9F1NaNdOSG
f9WbWXVgeO7COV7DaXcl3rr+0O2JKT3t72ycE+jkHWMAWnNcis2vp996TkZDioGi
z3j+A65VNSEuxKip/NZXTA9RvbB4ZVArV2ymt7/Wd6SJWsMZNkRKs+my27Xxv+La
+dLm1YTfD6dXSo0NbwCHrYAn19a9jFeXDQwRAiYhfWTnG6YOPs09NAWpNVtMUgKx
ODNp0Ptkapfgo5Prfm6+G4R+bX5N8H8NpBut/W7Iix2CKsFWF844cBzQU09N9G3q
b94bsb474VE6uuSFsFRoRYWRm2uGb5sXyMihb+UZvb8hm3OOFiephIK/9pvsF07h
BCNPDY8y+0Pb+7KcDI8yyKQobtbuZZsAj3LFal8egmMA8yHKdsA95GW+bzOIsgMM
RAy7xUo7CtFMbv61JIkVOQ0ZSFqDq4TZOBG+5/uliq04AFEDblT9rainogIL3vFQ
I38ytZUrd7mrKl5OP5Uh80M1SSbD7GSnwhUErzD8eOL/nY6WW5pSTDuKeCvHdLqB
8lai5zzrsRj5EGz5MuXwmKIQmJgTrZqmPgGd6B6ERorF5sSFDiEv/zLd58MPgb7W
0UmdavBZTLIlxlwiatpUbhod69WfCXzoPHr+wCrMvjtSzZFK8lvb5z99f0MZ5MOZ
aos4WNZDdzKwaYQyzO9LHCPQDK/YcMscfKcOgLv1FJgzUXZltbSMFHcmeWE8cesV
t/k1qfIeBbDOu5PrtpGYiIB5qNRuaTROD/hSQhJMLAhL767g35Cv5mbxa1ehvwJm
hpHYnZcY8YSebf0hiP4ec/xKXYqsBfF+2jXRawNN3D3L+I9X/4Kif4JrGGiD1+Ue
2fLh/hi0NGCWHjC00PI8UlcDqa/QJD9UjqxBcyj8WmEt1V7pa9p4OYn4mfYNTCxV
1bMdH7Ywnom5JCJ12F5bwAEs2RvMqmR5qYm2ElqAj42ZlRg5AKUkzTa4PhCdnZFZ
bxkcLAh6F8AuMotYKFC0OL6I2ggcVz4UU36SA4H1rrlav91KYkypBokYCpK1KKk9
oSa/h1vH3TtSCiYun9SviISBfpis0C2LshtCyp8HM/7DmrNLehCpuWrXPOE/i0PZ
Whe5tuRj+pGy5Zc87sppYD2M3yEXSyEMkehBuNQpIG7KmzwRASma/QENJCea3BoQ
w8O/pRLqWjN5GM+UyQfQIFrj1NtQWfc9MYCJtwbI3Pbmzlh8CDePUV+/p1eGWuun
jQVDzlPL5RMDLWOSr+tG/UAiYoWaVgRvU3TiqFzEFaurFCY3WxLtLv5asODOTNCs
40BUg9zlUuGKynvh7aiMxwHoWpkxx9DjwbjNRQYvHmSPnKPOO6iTo4IiRCihokBp
cfk5Zz7lazGthz7W7zDhjKAz0LIpYbLDfw2aEqZE76x6gJnJ1D1NzEb6AfD6ALW8
SF7IHjFHMjvIJG5rXD+XHXttXSvwL5oKJco5LvUbh3yCjXmX3b0rs2x1IB6kTMAj
hGbMB6YNjUax+52OBMAXRbRnzJ/2u3P3WZiI5deIzRfUF3Unngeo5WxB6MqqMXI+
vVXC05xx9CFy50IyEYXfUUyrR9Ag01YmKn/u1BE+zXXkTuZiWEHwsHf9B9PZfg2o
0beZ7Gb/LivBzdSpWvBLdmUYjteOue6Q/IpPDMwkByO3PHW1vGgHgxCyQqUl+lMH
oQxOj2rpoJ6LKH+NQcdhbTQygXIkCyIrsWpvT7iVKydW+2Tdcm1dcealenzdPaiX
uedJjKo5mkRq1Owg5ybMwVhwx+lyn5vmQOHrQXvNGa2eiU6/sqTckp+QZ44Md21u
lWpDu5NpNdC0ubAr2kwgZ0PDlK1drV1SMOOjOrXDVtTRen3guduVRi1aYUD3NPk+
S638wgPbzuAMfl/dR/kv5C0QRMH3XM5P8icdr999EwtcTgNrPEKh46bRjrfcfpza
1zO9qT38WEqj8/LG+RhhNFrYiM6nY9lSfUC5a8eXilNuyD/bHGh8JcZmGVU6PFC0
PZWN5KW+aAYJM+wC/UmUHsPpCID02GQ8ecSl2DK++IUE1MM+cFHZmKr4j30dsMTE
ViVZyCJNu+zTvJ8jZK3feAUShCtYS2ZCwu3qpFamKv2KmQBmpPAcQ52J6Icwrkkx
+dFFvgD6uDEXqcDql5PtfH0U1Bz2R+1y/awZ1/WNHrO7UT2Q8ZC5F6dNUE2H4Yiq
vnafQrOpZ0Zel1mFkYWIchWEpqDWbN3f8eLi2kDJFGdIlEZ/9Xzkfb8oVC0Acbo4
qx7MfTVYlITN+uBaVQY3yLonCdIAE8YcKRNyRZw0zEHgFbiSWZ/S7EAX2a037rRN
841Hl4GiBF3G4WsIA18bCONcgeXQfmnU5UoVwDlmaBh2anNWso9k0nP6gSCCFVtK
Sj2O9bU5NL3cU1yj62jwF8tadxxM2FLM+HEwwiXc52HaUTFhnr5aq9VEWPDQt5hM
IdVWmxm2OZMQcMiuFB/OU5R7Ep6NMgJ1sDmeY/d53hmnjwLZI16vMxQY1lHqgM/j
Qq43TWsbNDyi6NSk+X6MzS8WyoQFDUJ3FZYyJGtQ1gbHkjCKixWHRfEBt4bWoueS
cr5v4iffT0dc0YaN40JHZCM1J/exe9JB/WKGhxNOpCrlAkbQI8F+9Xl5KYRAGF/Y
2+g9Y3v3f+xz0bNjNZYO5bzwZWPBpwwASFjXjuWb1hAelgpeWc8DS1BmR+JlnvZL
GuclG3Qn+iM7e978L3j9oDk1uFnixXQ7NrNyjNrpKhjJlPxhqrSVWw4IGcltRR9D
JODiXTSBdm4FgWeH1MUCRNUQSfRe7RCd9K7XvBB84XeXAqV6EzwncXyN9PsUbI3f
5ceOjz5PiAsHwgcT7YUTftQwPlScPF5OPznZmylZ/psJFEBmzOC5aMLWTI6aGg3L
H9SnaQExqdlV8QdCln7WubvZirgJcHU46hECQAwBM23mcbsnDrb1saAla36pv5G1
oRIUFPkBHEFv5/IaTwPqLYgI1H2P8HFqMMdBwVd7eP1+vm4WX4XhdVBJS73nMaaV
IXBA0ZQC6jXWNSAvXDTqijEQg9xi7ACZjjvgY/yF9PD49M4556VMMhs0tVs6k1hj
cRAcOdqIuJMmEdg2kBZsIiI/KqtM1WAW4GwsWVcvM2BJJJWAZ5S8AvtSlfM/8u5i
nAUMUV+Rq29FTQ315GZ3maS/N8hkIeT2qYs4HMH+aVjNzg7EUWHUZNmgLox1K5C9
FgVxt3KVvvqwA5lLkrrniL+sr387kIM+2KAmDrGKkGXTiKBzWt8HSbrI1CI6UYHF
nakEpjLiNvu+Led7PmIe3YeKjJOCyxuXMs+sVmBBH5mF2B8Gn+cObxdg09L0rVO5
MXyQbMA+m5AVOppfNxo6f/Fn/3WxF1ooq2Vy7GtuJdCuLzFQ84mKYQ2hyBv2IqTj
pMv20jfy8+pf+w29qyO59AzvEIepE36HZC7+6j/tew9sWSOKmS3Wb4II4QnpysiO
MJhsy5hWR3J31fw2FVlyzZFsGAN1RFQdH9QcPPG2qeoBPIKp8izpGUBMd6t3bjh7
pX1AYULv0Q7+z3/NY7HH4k32DDIol8nwIM7WBzndH+QHNRvEi9LC5/6p/8xRjgKr
o2tVEserTsTrgCxM0JXPKHVNXwDWjQcfcAucBSwYWskjk4cZE7ckoQBPKVcWVLxz
wNbL+ys04PJKw610/xS3mkUxBQJH2vn/AMmHRlkaiAUMBvFYFTinxHqXMMTLFbMP
MD1NBdgKaapzgtk6Am/W6Gz4xXRsGzKKTCWDtqyxakUYpZxgrf+eF/EY0sURQecU
RL3yszSgHtfnoDFXggJ/QPJez/AEw0QtQxCiK5IeUqr+uDXKO5r6J2xaqfoMEXin
DYjLuxw0azk4yyDllnyZlnZgt1LmXV+cUwdKlSAzyL/QsiBY2NjzVde6KxDWzPAQ
HfO/sGjeKyWE3OTVhF9UQ5XXRK+XvrRRQbv9uh8UFK2mYA0YHh+qAfMGZkxfCoKF
n5CZbd3nbDsPK7vaKaKG5H3rD0LbwyZeulD2az+cTEEiCtZOFiJVnN1Bf/K52N+r
wmwuPUNHoX1gMYNsbdIF55cdfylH1S1LE7oPLNPeC95qMdENsDmvd21Us5YNDXLJ
bEYX6iVL4jUUMDfsIiWjFJ/9FfXB3Zlp3gIkwzVLRuewpXyLG+//jwD0cUeVrseD
BgF9xPKXhAu4tifrG1qgZH92xtvdT6dMUvI5ntluVmPtYvb04BFV5h4IRERzwW7T
9CYHM4DO48ZzvFsSe/MYBBAyYxl4kni1C01tUaKW6PWOSjMw1p/pJJQDL6hH94AG
clq1NZKoTuYGqeJ0pJouyuG7ZDewWoviizlaTT3OA9Ff2RkRtywPMk+/N4ugDqYf
39WuETQYplnYZMYMt7gfzpjpfrn11XGvYfw3VS1fD2NdvlUfERY1bSXhPyeCh0/0
hJUHTzAGLoC6q2JgAiuuWUw+q0vfn8T0dMbKV1k28GspLrapHWs4P3cAaXq97dGg
qmf1uJxmje80e1dga8fSi/tI63PY3MeMK+a2T+sAA09ID2QzZXm3YJIWWrp632+X
3MGELF0ODi/wSLJtF7a7bjX+W9Rd33JajcUYbgcLwU5FBE8ERbnMobkXHY8cueEQ
wka0I6qZIf1diWIYDlb/WYPSDihJ0E9sBL6GBcbMZwh0qoaSne75bSApg3C+rWCe
aQ5evh3/q7isuOPveiFb4SSA4fCGmCe05ZlFGWod+qkXT5rz1bjb6JkUMPhqh+hO
uvsob2I+/Zst69ZlzmASrCf7djURp7OSL3FZwdCXzgDxnJ5bxyv/+c9n/5U4PnLK
tQV4kO0lh6QHYesYhj0iOQ+j73Hs1o2NZE6Edm0ehXCfR7xM7wlCii16CoJNtzUb
VefMlJOQo9pE8HVjdrZM6tk5z7MozNvMpubpDtwenz2LgZNlqIdXT6JfJiqoKdCB
+fC1OmuQPuPlLEwbvfz+J6Qxz6BRjEmQWkP3eIuCOBDI5AGI/kmPNFDIB4UB20gF
ANa/EytH2Nla5wXiJIZCcFDYeLmKjd/J514Gq2MWW+5Sec160zXwXP4G60GnuqGY
SMz7IhYz61N5BM9C31Z2YHu2aVOZNV7IN69q5OCl4NZDuaDqLAO6QU9RgbMP0QfV
Qnr4mKNodeywuDfPYLtLYehy6VF+DXJ32otjOGIhIDw3Iuu58GxOX+iLvfS2I6hI
0ii3kLr/Xc01k5ts24KJCwPIP0QHF34Y1kKvZw7zOw3Iv9qeMZQtwW0dlEeU6cbH
adn8c2py5ZoE/ZO5iZRS/ZHbNerrXu2700aRwLlMlLH88uinRynnUtWfMwmunatp
zD/q3kKaepryR+QW8vYrS6I0S0nV2KeEih2AlE72WB1yxDZzkKgWqoHQXxTVPFT5
s+VZVVvEAytcRhaWre7xHIZMWIpQazKDa2go+W3gWaQR944UtM5r1VA2MncUcHAn
aAdCT/ynzDyziP6XX+yksgLayEhbbYOimxWlwJ6U55hmQ2g7agYll/rKNIrINTfR
tTLi1QhqXDLf7gruz9UxYcoYdtBomB98FKw7aUyelD/kAGOTM6nwIcaoKC0p2IAJ
5mQzp3pspZsR6VeC6GhUiylfEEWP83nZ+YSOd7Nixju7YuJ5R1UQlFRmOK4PmsOS
+X3WES/PJsmjuL1yztrGeVB9VbTlnA9mJ5R9x/JNAZyZnn/Hy4VK/TNy20g2M0Tm
D5JIkATUL24onyf70OxMmi0u58ZB+ylcZFeYn+HRbOLo+sh9GmvGlsRtS8orhFXY
nRlQVG04zLmSX/u8adYc++ltBzveGKmd+npRDKbYD8M5/x2ztR4TNWdRunIV8ixD
1yEo6hywXFVqrVIBJXCHehHt2Vr/bJ4XDcstYEW9omCGTJrN3T5Rg+pS7h8OIhxh
gN+FsLY8T1cuVen4IiLPscXJTphYGs0C8rL2Vj8ASnjCgu9OUUlVcBTzQCjWExzG
yWPxShuFHJDryPy9dOeDBgIjSqTKc42qTTHKKFOJkuLyb2d/UeSlYWlbQXTJAQuH
V8xfkyey9Vi0VElFRFS9tprJVg8FOY+uZxmFIyufwpkl1io0lTh3p+BDrHgjO7Gz
YaXNhv5sWg9i7doyvICCCWott45Kq6yfJ/HZ/cqG32cCbvpiILpBlZL6JqJavdqb
eXapHPNnRNIcRZ5XniTsbWpatCPUTxwIDuD4Njk+a/YwXDEc+JS9B98HzG4nxPCL
d1V/b59Pxe8qeXjZorivFAfDdgirlGJ3ZBc5fP87ihbCTHhnDvbcrOoKT3ccM25f
P/Aefw3MJ3Dq0sCx4Z9Js1wdnX+zTm6L584iYPXhiz1/WQ7EnZbishoToDKciqwI
RpqR4JnqTbqbEUoOTG3Di6AFDpfcKi8OuPn0YuI3n352xSR8HWQ/AQ98o8O3J5yV
i/5k7I11G0GJT4CzF83GAESWWTGew6sK8CL2CgRLh6ZNC4CPwedFBI4c9rHS6AKF
loEzkm9HCYUknvv5NtxeoZq6tzS78DIdlhHcRBH7Xwag+uYc9UEjqI9SSzFzjuC+
AN8f0mbHK07OedeD4Rgo5KzJ4SbBIS8W6RFOy6X89gGH6/iTC/uo2dcYgIn7TnsG
hLzYphKzPztwD0xqRADLHepedkkQvjbExtcjw8sR0RHJ8f7g3hOYCcnGDslXeLhy
u0k5VMzru2Xyjk79TDTe3B/93akt4kaBUx7E/f5sHIjZNrd1IeughAiX7w15kuTr
NoiXLYV5CNCBMoiURulF8//vc0Oe5PsQNa/Hz5Qjip2zXA4U0aOGf+tnFjteZpoK
TuFDv++dz3WwqZbMzFGRt6yEMS/HzCGnhTBxzKJPibzvE+jE6zsSyZWbCX3CofO3
8iG9XRKVtowU606MkvMG/z0Pm10vqkcAaYmM8IeSHNJbTlRYOSEVyqCHrXQFNIvF
1HT1rKnXGauvXmw3DgA6kZCE0C7bHom5To2646tf+JHBuuoAYW/nJ6wImSp/jZZs
ufy+04V7ugNbdNi2mttbuwJLBFMb9chS7/DdaV70btmvOBfbheGrA4+C8YctMmam
Thjm8ELh+8ey8LLJik6iaUz9T+VP+PwdVw3j9YVROKrD4K+nNoo4pyt1uo0Gy/kA
Zw/ys5EpmHjZycCuGX0kI9Hr4g26uJQKDm5vYmyyMjFRJPXtMWxPpsbNTSWSXrsh
8jH8AJwUrXk/syxrpKBIixGdM82EiKMblzCRb8eK2LaGIqVDd5v9IqhXz5BAaQ7H
Ib2BTO1v9GrTb+rQppnZBwpmkQuiiXh4Rek57fcSKUId9udnRwKmk//m8hP8xwXP
b+HMg1a+RjicP2tw3lYB7cz4e2dtq4iIG16Mzd2v2cgkqSsA6ofQUtoYMDNRQxGj
sXt9QE8r1yONHSfxwizPR1l8FmEa4Zuk6Nx7ep8YL8kuwQzGwpkb7BTS76g1TZZL
/DD04WyhbzQWv8Le/RyrMdOFiQkulHelpmwp7aX2g1TjJ3ZSm5CUfboDK2o0ROhO
fRwsHlxT4W2IPJgMIoQaVTqe02QYQEPfhO97+PJoWSN01j6/4YSTLykbe5PaOq88
uyG5yCbCUZdAwvZdC1cBB1oR0/xxmCILS27HkWMPjfY2zEmg2jRRrFMvZXCCAp64
ra2I7RBrIqnPTrrAHW15xhCUIiYvRlgxOKb6Vkz4WChWt4uSAp8WuMuVx+QYHnH7
m195f+vVOqJhpu+exAeJvnUBQNkQ2uolWy6WPzZqw6oriV2D0+apBvFCY1auPlG0
l5pNIeFGhxA0JXtjOSUGhpPBypdC+GIb+t2CjwsaYNS8lafZ9WmBsLBmBu3tCtn6
gYjH7K0sghHxnz0XsX1VfyIB1QBSxs17v7lwRg8I4ySw32ifa+xzY+q0X5TB8tgX
XYK361e9f4HMIT1K/N2CzxJYSdI3xgEf5wMvpLmVrF5maFE1+lCRqlnqSI1L6LTV
WdpWCD6/931BBvDbZkRvlkH3R7yeOE9haZuso12+zHPkAOpbNkUEZqr/b3aH6bOz
6vAT+w4qiYWta00P24sVDXef9Ao+FQlrNNDAZbsP9jUbV4ho2x3LOWQUAMlB2If7
8LAiMZxNjOA/DyiY4oGNewP+Pekw0oflOfDRgZ7WtAUBxMXD/C+8ASQbfmmVVTQN
nv7nR9xaXZ53My8bZtMC2njwJm4mXC5F6SLbw257CEWxu2jjV9oWoUn16yYbtBOl
Y60sZ359aKT9YZqtII+F1sBU1N37VBUwxLPWFdHTvUMPmHUmGP2JoFwDo+SurTFR
+1ZO+6VhlfO4dQl+kVVcTJNaYhj+nIQWWUMN8v+Uw69tOHaesqHsoTJrVIDAAZZ4
1SjLmwGgSZkS502RNbxhA1U3WW3cuqV4vdPIsT28r31Dta0Uwk/dEKBcqC4WaLlq
2wfzwpyJb7v9S66PzXy6VR2GX+iowBlL5r+efEwMSy+nfwT81cKnvNLlOTfK/vgP
GDROGfgxvl5esg4IHFZf7y/mQ1TnML2sKFgTfc1V0PBnE7+jpWluvNnwphmrhthF
OUFbRVXxfXLCPuQ7Sv0ybJG/6MVGpIGECglvYiUtUj1uRROFVXaUovveoQhvRpSG
MTGVChIBXG5qKF4HreEgj/GbIWaJaGeN+rTrKoTOs553LB1ppNedAfDhwYXJRY06
CqhqOF9/XT9rXutUdF13O2YqK0H/zf/N7ry4Kgxc/k3L1j/EP4DhrG6N4ph36q1H
xW7dz40xGiYx2xwQ1dd5xfXLdYRL+AU5KBMmzU9f9yjExcPbLrIJQCSabVl29PiQ
AtzR52QQPkXxb9m2qcbNx7uhjX11DLMk79bvULkdvCDTXgk8Frv7DMM3uxG2S+lZ
j7LSatAeNvurrgUrc/Zx4BypkozbNpXl7Q5HT/oHcmw/Gh2BHTZH0b8beLeSoSwc
II07JL+q7+RItqh7IB2L6thcNq72D41ImfXOjZXSrjLqVtAeg34MyxHcLDNJ8wYg
+GM/RhB3quf5DVm9Pj86+I1Tag+o9UNCi5br/9i+c2hoS+Ziv9lUhiKb15km4m9n
P6L6Vkr+Y2INQO46vzyI4aMGKiyxeCgPPA8tIFfJekKCrQMYc8UccWn1TG6kSOx4
RKYzsqfXJuaeavs31CZBcrp9BjiqgQDD4xZX5O1dcAjKKaEuxSKL63AeE0LxcYpY
Zx2redlNP3BzjKt95ICiq5lq4JhRUGhIuP/QSX536YtfeCmqmjtlYaUAB5f59sUY
VCzXTOjEO7zOJndDPdOcSYLi3bcfbNxLXr85ausB2vMz6UAD3olS0w+xNnxx0/nT
+DBHHpvUVjj6hiWjxmw/UTNX9virhpdAP6N9Rin6sCmSCq6gW8Fi7CSBDn6M1hb5
8JCJfe6JTNw8TorPfns31277A12qlYhm/zJDAf18exLAcNjCvjK7TVHNxeL3Y7kN
8MHptAaTlbqly3NV94H+6KskHi6235garsrhZepP3DOggX+068qENUXxMBzV7Hc+
aHnpnNxJDAL2xd5YgCAJCk3aB9ckMTXyobMrAFjJXCHE5WsuqOXKpuKDpd+hweRg
3tH+eeylbzCitUBRBZvIvsOf4/X3odNnOWllkCQwn/zKrOGfkRINsWhgiMVOU+rV
`pragma protect end_protected
