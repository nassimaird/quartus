// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VJRCfArd4CuaeIWOwUYb602HQFjbJPJej5wz1SNl2HQITP/vUJ8gYhnPNMBNPzjpVRwIyFsBj665
re02Qmr2J8r7ab2tcVEAJr8WgT0F4/h3chUU6jUowt264ORfa9XtwWhsl22WW0iArvCH3PI0WkyD
KFIicOMq7MjZE0qF7391v068bIHdhQ//G56/QBs2VeNT8471y46TBIDrFAZvddGW2KDH2+RAsx2J
uA5j2hggQFdqhvH0t59+qIfksVQ65hU93UagArBQrclqCYNKpesBlpsM09FcXw7qk9pl0LYeG7yh
rR+tDJVTmixXViqcXwJ3G6iyQccGemIpgP/jDA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31040)
xb2Dqq/jFDagnE8/Z6GeWp/EeHwF5SBIViMJn7ShEfIUqGfeQ7hKZykmCXLOt+wCe7tajmmIxide
vzugJp9KQeEAdtH/l+Ij0qNBiOEl6+YCsepCHLTdWsZXJJQy3udlUR372z+OwlQl10VEok355QvQ
CFGE1kQX1nxpDghpE0ifov+oKlTf98MHE/e8mpQ5E3dPQcc8I+23jWBFdoSICrhXPGkKsbmF24sK
Owmd5fgAAfGnogeeSF60lTh6s6CGb6K2C2Vf838xC17INIDjefs77qarFTS9OfRZvNYPPCZ4zcW0
lyaSQriKaUS7vOYUS+R225l51lKmaaeABa4OeDF9fCYrwqB4cn5pu1c0iWdxDfKerduNR/TNdZTC
syz501v+I1j9vSB9F6ldJQy2uLgGUhZ9alPD2l+UK7ysbSvT4J5GLaBb5MrCutpaJNbSCYQ4ly+3
GESMcGJXtRF4bASjQ27kWgrxcLxY5MfU/Hk2WEiDzN0DX3l5v5NM7Y1Ii7kF0VZJQwIh5DVMyhJd
tVFTU0R6wedcmZDZ5/yBwhcpt+OXG8S/StzfAq3H/k4032Ge2epUr+zQh6fcQt+BGKbRujrg0AQd
UHOnQfgVXzeTY6DjTD9BiPEjapwDiSIAJJSqQFPalW2Ul76HBFAMHARcZqlPA+puecCJTez1IgkP
VWyxO6Tz+D2TlG9NZ1lAAT0xWnL9Yif7036yYk5fP/2rKhzZNAyFpWEQAtxn+zpS8PemDgscR0hC
qjmPmcWmX67/94jrgY0XpqM9JRlwZFig9EdDHntGhHDOxaPUSaw0azaTryx2h7bqmjDBuDyRQTdL
ZDp2jqh3LkyaDYsHQ1Mx/bJPVrW5WTkp3/xGqIzaGG+oTdNLnMnynJHkzYDmQeCRFOx7rXnTe0yE
GpCZhJU1xHTmr8l88VT5QuaWoB/i09h1NkvVUzSeIRe29k38HrAJyD7Tz2dxN7v5wxc/EeM5Jpj6
xLRygF+pVEzzN8BT0mwX3DgRZuFFUu0Z0NL7syuzWsvgk70Poib171lQWSQvkuO3tyutfCj1KT0c
UqkPLTNvqy1x9/Bufzckb1r7Ak4mFoK/VM0ugvkEz5BXfkpNY3jJ13YK1QggTBjO4+KaaRXh82SD
gQ5SHAzfqVexpIybE4wv2gkre2jlFkIUNjzWktSFEPyRaYRsgGydlZ/jlBXQdPRYT+IbuvtZiFDD
d9WrC3bOoKV4LmWM3eMfvEMaYA+V63DBQ2UGS/zrBxwUy7hPYlGW1wCdKcja+VdCKzNAxFCSyCRp
68MjPzRzPsaIkSYVdEHf7m4QiLAiooWyseGiZlDTGGs3OxURHyxSNPOMoxtEM3daNRcF+NAaqGlo
k5nZTiVLyDTN1EuEi45SqXBn3cOj5VW4pT3rQ6D6fBJliZ0UdKmsSDQf9OYp7WvGUgPym91Nb2Gq
Q8KKCBY60B+LNsX+pdwO7qDMm3L/kyIT7+LzU0mDOE59BeT+aRhk74G0qGyd1czeuJoduzaN3ez0
AQ8YKz8PLXWvd9JUexqawXZq+naYAk5zIn74raDusQMXYU285KEhhUIYV7Xk0pZu1h3w1o6VVKIx
+TDhBrNpaghvAo/j4SkXtMsFkAZhZ7Y9YlMlJ1a7PmeatE98TLQ+vVcUv/uQVr7pjcsJl0xSA3UU
A+SD6C9afkIk9LuZiZ9tlAqTXWNKsv/w8j0JLYqtCH/n1czLSu1Q1P4ERSv9J6sTaK7x5DWZXeVc
/RfsMKrlH3BtkR4nx4r82m7EPMG3F9tD0lKAEr+xy9NBTacWcXDa2QaIscRX/TXFZgQsadCHfcJY
jFjKDZzj7+p5NegyuQQAwOysEI0y2iiZyXjCMK7wmMAd4zzdVsQX/3aSxt1xvm3JwNm20XjvsQUT
//Xz5VjLNF5CJMtFfjOzBL2poZtbG8bOTdrc27soVPSPXuOhvc5qrWQivjyE+zXXLjkJ6d9/cHZ3
gGELAZk0eVWx9QMeDXVUWLMoG25By6UeXbVT8OOjQwiZLB9Z63wCE/CcQBKhzCYwITI8QPpEeLGi
gjpGCgY1Q2+NON73TxitsiWOFB7hCiyhnoM68OvogTybWuQHE9oy2PvW54US7DAW7azSQCT1joQC
rBmx20U7iF3eT4bW4DU5CegdSYZCnHwHnsosK+h1SgKRcr7bx9d2rIvVYk14aibOHghFmq8/JC+e
YSfrf7lK0K7O5UlOEJ9KfvJUpDx9pFPo4fF48dE/BH+2RnFCXv6wuy1Ne2sx8sgsNLdxHF+B/fHy
IiAidTJZ1VCfV4fMuEIPR5aDfrOIJKZDCwNALEHGe74uLFmb5N2n+gpvMfzl7hLw2dzf/TDumI+b
yXQ/8q3w0D9sWQb9I6oEG6UTpd02ECdu/aeZSfYWZMWrUV+0fXWZFNbTkRycdXqORmoHqAx6AXFE
50TafIxNfSqNER7nhcL5n4JIVJZpXJ/obQYjGkO6gumOlDlMMcU8n7SIskyeB2mzmOrKnY+lGLb4
WRpYTIUu5q/a2l/5+B528j3RXe8VVfbOzAgZNMwNf1GrgX8zSGAOa9fsAussDLlrsQQLn3hA2lxT
o65fCXHzdgB/XrVEz6CwAO1j2k9SYWhE7G9aESY27n9IbSHdlOqhUWKgYk+S8v6QTiY1g3ybmMlS
xyiu8BjazBCswoWLpykbvqKugS7FTJDsUS5uCjm6SAZTIPT7ueD5MzluYFpuQXr327CpyHQofAlF
yBxhx7+vrn+OCM3uTCPKaByd4YKD5eJcGaxIkFe/il4LVR3CR54ABJTeRlUImeaoGPvp/lA/yRxm
PL/oeqVxmbTfBfPZrMyYT2VY+NfNOfH4v2xd+2BuotpbkZWdI7eJ8lQFejPqqz0KvolRqFXRn9zO
kta29GlO8yDF6CfP8VOa/RLUG/iKFI85uNyfFrlg4zxM2Tj6yofXBpT5FEDqHyHxy1qy+x+3Bxgh
XgjfI4O3CwMPQuPE0wI6db87X7d9TRimxWmkFXxC9CHzPM8VJ0RfFsEzWB5QtwnnJshOwtYwHpzs
IJVSI4xGyvXCxomWGd/fMeZNC/wfNQ8I6Yh4NB9uIuLUXRGWGo5EwvckQCJoLrmun0RHV3ZG917A
Cm8LcdbOPKxetjodX39l8eB9TI38+WoEQPhwlb9BDkM9jYrlemAtCqG+qOImaY1uFul5QyM/N5rq
RyV2jgYxjl+1sgqMDmG/nlU+oGMit6Uq5Cc6mP4w3E4qMQ59WHMXlI4Pvo0Vu0DWTVqtlSCckeqS
dQdJ+PzWZrkrBrGJkH4B7tR7PSZdcd08olxSBqYElgEonOGIhNF/V2fw0NWRx4iOh72ThHdZhgIC
vubuXlhn1qwouMSlx1lm6OqgvIAq6u2fnLQs7fRLGa2DRZb8wTnDSXh8WvRwrZ9dAEDnzDp1D+KK
K+13HDrQqYNYVvjGZV9iGFvysjF1W8wKEhHSYb/grkafJpHNwyGmdoC3lI4bbTQpKN82luYtOtlv
GVmWBWJmTy1F2EnsmBA7Fg8QdozYYXZpwyjy7Mlg6YmhDooBkGZUX5nqPeAB+dZeD6neTWvyf+cc
pwdJt9/dfDTCbrV+zbl0w8wPOBh98f5rzkw3O29CftNYCAXkGfqq2mZdlXSzbT6tfg/cEj+vixap
I57QboHUJzVFGD2XIkdRXyzLTpA45sBY8sjS5jh68lvSQVVB8zYWVRcbP1QBD9b1P1iLFU91MMVw
BlGjregVERymvL1GW2zV2j7JhgJTIrwGVgYG5OPfFSgyjtTIDcRX7vuzkqXL8XgAzZt5qr+78DLK
OJuQWEcS7k+xre4KmMZLV9aAmgDt8dF0S9t56l2DI4/Ag0/aweYI4CTXlsC6s1DlV19KeP5kUxV+
oV68R/o1fTncOIwk1kWp4NEfjD+PN+cznBOjyMmmONBA5dviawOIVMyFmBaKytw6rZzXlYbdNVqE
U+51CzRkLlMLGhq6BEsgEDMo0kQEEwnmqugH6W85Ry/uRsGZ2uM2j8mJB/swzyj/GL7BE1aAn8RI
sBv61U8oXDydwYvegt/QidD0DgJMPk+ahq9OYARiIbGHaHKo//4/137Au5W+NNiinQfuCxWVDO7N
xweL0dQbV1bpJfVsVT9AVMNDtTGUJ27Kvij2+xFyQmjiGKfOzQvjCnLUcvEcdAxrQeENdzXEcm7Y
t70Z8Ufma6r71yUq/RXfcHXbuKMVPG580SNHGGtAgux8JHSKAAiATL2idAu8/afzGm1oPMWxGsr+
pR4Fr0mDTe/PYG6vQFki2pO2F5VYDi1MxIkZXnYzy6urjyY0cAZ8obqLkJfCAY6YuJqnXZgYcIBr
6+XpxNfAp7dTZuRtnsqTMH79wtavw0+Y4tRIALP97qnHbr7t2yfhTLM9xCWue0GK7djn2NHjvjpu
djFEGxLX+0n+H0PVtrwHtNLrGKr/3dlcaX+otXvVJo5G5YDWEyKNzbu/lHr3YAALQdHc899Tiv5q
08rDz9zYCmgohViY2BVfJnygwUekFiWU4S/YCJaakGZ1hChWHhuZsJBBdwGWpnayB9EAa9wappLc
B4mgTN1JOzLvQEv2Fw5QJHGdD8bBmwe3JKpqGKuzMaDgyqrPAWt7voU/yERYDp/AN9FSHXeszEiA
T3RS5EfdVJBMJtxY8LX2ROt0/8zgt87NQaAL1NvSuiLiAydQp4QBCDmYTjBlKCD9Z6aFSBl6Nito
U7HebmV29+zVWJYY4ItmhmpUGOBFWfOfSzFsa56LMuqpCoiH278RxshFeTVd8hdba3ToK6+7H6wz
hPs9mRTKd2b4my35qmCmgMxbd6NwK4UUPDymLPj/sAoF1uA51/f1zY4VsvxATfONBi4DHpzqIcd+
IxFuFTzXQzPa8DkCSSTsslHYETx8ejV8Fv78ZeQlUJuNce/IQQHJ+AFuHoNp4d1JFRPZmvMO8smc
H9P4YfIGJyoVsSwh6WLw7cPH2iuWHfSTLobT0BLk6azu1bom8xYlHpYIDxT3iBpw71OMehoqIHFo
iqW2v2LczkZ4RR8OzOr6fznJ8IhQHnLfGzmdMH9awV4rsE60icohT4D0tW/l8eqP4Muja6wcYyL2
Ofm7LNdmRFfgzHnAjeX7EYjnC3cfsLAZAb9agWsJpkEAolh7N1nx5wuUH2HSQ+vgTp7Q0m6791s8
Dd/EtXuyzUBIzndTa7sFW4Bh0riEDXa613CsFR9cgZFZTI4NaEok3bKbOC4UoP3T8CYG5y30mij5
aaXQsVLt4xDDSRCcKQXP504YotJAID5X7ZcMHuw0ilQqPvWGe1w2+PobAWTDTro6ZtwiyN/HhNBF
SF34nMz8RgV1L1Fz51q2yoO+kW4pPc8yHW/IinXW8l/Ac7/QOpJhLDy6yToqppKhlwi/yueMaPxF
e8tG7hNDPRzoPZUyo/Civ50uh1WSSW3WFf42hCIY9hwwxiYUtn1uyvU4rRczRgLlJ7bM87WXtEK6
WSfL7amkkQvem9eEjaMK5uvV9sQyzhUxPqkuEyEEQgj0J5rqCCrF671krTLkIfRRwDzVmI9H/mON
8Yv1XaEoOwWxw9D9uxF25FwhdIUJnXZLXvIq7H7WZ3wSBgOozcANERKGRIjH4W5YegHWpEJIfKND
h3FnXnL8XasB3QETcJeh0CQHO3CKR5Z7ipR0TEQYPoYJ6tc8clksOWidoehNl9QYNj8JKfdel37F
vU5TubothI6sRc/nEw3haVeYH2ajF4wYRpxjq+Oq/+82595M9NYr0OJHELm4ZN898/7092fXWcEa
v+3W2vfKKnB82qfWu1gBWFlWBX/UG73Qyqui308Lhq0QSvcuZKGEFb9POuozk/Q6hTRP2FdUEXUa
NSAxxtAqTNnzgKt5CXhJU19y/5Qd5RzlbuwgFuRlWDh0Le9n4CYZGnK9KJiCGmYuT+n7dxtsDjpT
c1hcrjR1RJYQRH0SiT/GoX2vd5dU6qynoTcvrQW4Okd6lEWoAE0i7482+EJSRe+7E+1OdE6SmcTJ
90ceQwUnkcMJ7OjIu//+AZNaiSQ9AAgihaFT1YSTunorvqZsei6Z5IfcjA5W9TksHz1bSP+owthg
MTx6U0sdFQpF38HzhMS0N/TBHBUZilcQDKf9U92nXc0zndx+94vBmzVpJKLbECI8XJCoRGOBhCoN
p3b9AWFbYbdIUDyuO+piJXJ/lJSPBSsVnz30gWZuBC+M2cv0sYcc/Vi0m0XIQE+n+ElbiL/tS9HY
VCYSb6ZibCVr+rhYHQA0rbOWsZpu/th/JSPAlueXAWnc+y2AQbRyUWbh9EC7dG9Y5Ni0jdOa+lrx
qq1m2L1qYEHIbqMXfwMkX8lMcNY6l2A6VZYQncHGwKhBxLp9YKNzQP/0eg71brrjwHrUzZckBmt3
dxqg0UqcX+Y8pMc2+JmV7HHQwp1be3mMzN/6jat2Uh5GnSaABZhFYZE6Nizi9bvyhPvsCESrtTAf
xx8Y0IxdCfusp7WDWMYgPsUKMBTyWYwui6yjU1XiJjiNwZmWCrl9wjX9KH1yV61V0xEYvTNtQZdB
Ns/sNT/xqiH8qmmdkcO85rBLMS68yEUKpt/bucqwm7s2Gdskm73liaSQYoLPU+FM4Mf1xCuIqqMj
/gM9XExqJTOzELn7XZi8Wt/3EfWpQmUHfHkKenUIcM1znbE9KSCNWVfESUFtM+pdsDw3F2mjTqGC
A7wClll7vitWDkiw3YbY67iUFjamfedUX8Tcz1uev0qyrARi0LxtZevt4rP4cav2gGH5VnZW8E6b
HX1dZyv7/f+iEyqqA8jrB6MOtfr1m92Z0f16QoPjZGy+PdRQYInaqjF92E0MjDs6Pj54DXpBsbOb
Zqe8z5PTE2L9msj9w87YK0khASuQcYjxWMKw7GUCTnykrybKM3Ay7NJqwrh5BoHDTuyD7NXKuuAr
m025UkoDF81Epgg/EzW/sj1UDF+feewDdScTaf1bPAuRv4XGRcpXHq4YHlNnzKzRcxOeo/7Dy6MB
HoA3d8egbCgsXOJqJ1qPFwf7VNx0OBxdDK83IuhQ5J470jFS1E3RG2oE4Wsm1vI6giPjmMhlX2LP
b3ARB2cN2ZMSvhBwOA+QKlERlfwKBrLS9cqRZ+5x0eEjfLLPxm7OETFAsoPt38x52w4YnzlRTnLM
P1ey+lcLNGCoL8pDAwuqgI3N+Tk9qPk4KCPzJYvQdYgDUkuKwLNu7ysHs567l5i+hQh1BpyG11vK
fgMdM9hZKZT9viANcUchUxB6Fi2jnqh9nE+3n2NALLQYSRkh9e29TDLBKAOxDJ4S/FG71pwBnODo
mZiguKIjVEJEh77PGR2Tgffq9CpgwkXrs6tq29mdaeKLM6nlbdGf/5NaaKJ0qr3VvY9dsNEWzbKJ
tW5EbMmFzk0MM7Vl6wtW2+VZ3jaYNLh91GVYjBdAeKbnaa0hDjOn9w/9aJ81YunnZfjJUQYfzCWq
vZ/UJ6s3x0+RRCXV4KPSs2RbdVOWRxbKUKLJ2w7gf9P4UYUBhxgXN86uI/PpvfrkagjLkZuDtDJc
NaFXg2v00xSdSjem1MLavNIGAzbGtwkJVAhav048FgzN4+OgUMtCy32rU5chn2tYtkb5TWjQtE/I
4bctc8/8gJewGlgo11n4scV2LwfGnWYtpeBgHey4/Wl8cGjY4TABTdHvRHWglMPgY5zskkCifUUC
b987Qy4ZxmJk8U8vRxG/d/U5FCWqaLsKo2QXrOrXXtdmbeCpZeMr11hMjaSiJFe7iPzbG1q6o43w
/Ek9F+HqdVV64dVRua7ULrA7iabGmzyjnhQmpdZUS87OB25Wwu5pO2Yly1ZH88RI13ny9Dzxbk0t
f/RdCAJ9uN3cjbPvj5qiFj4DYDH87Gc/dBgKvTW59E8njiwgE91+Ov7ykc0nPwYYTloGVZZUBhrE
yvxBtmJeQuUo5M9scnTa66aF4Y1ufYgsDQjqVHbs55Hui7Ai/u+PeURmG19k0hps/5xFYdjiIlXN
NeFWPIhD+mMyiA/iSkSvoQCAe9W8hErX8hCjaXS7ytY2a7XJXcsN/YnBfaQj23NhLlnOe9WVxSxY
X3MHXlmjsJzmTdST4Iijh5iL/+X1rjK8fz1g0Yq3p5cJ6vAwC3cr44yl1qWU3KfgpEFxqp+xQQK3
fe//M8QpaYNV0GglGcePBk60A3FBhDbRJzvc+2wi7s9An/1sAjPG5tuLBQCo3wgN5B9nuxzVkg7q
3TWYKdBHoQAxEbdSMFhfbYQnYPBHtZC5pt3H030ZICGjnsDoC7gwCbv7+FiWap4gNHeSAloygl/W
YbRm/hl3uAx3oPVWFXO+9kOHgGiDvzA9bFwHn7wMZKlas8vXZU3T/ZlAFpwOflICgFITtL8T27Zf
3VBpNWDT6+KDRPKp8ftV+hNsv47W7mftTBJWo0euh38gIB5oaXaFB7S+xV05/NFKkHsCOmiuP13A
bA0JDYQ/PAUpcIvn663Vk6PdnVfJa0QGeJjUeAtiYf+2Pyjtam3+DK3tYdJT7ZjBLwHV8FwChUgU
wjsoERhKBRDfZDm532FrTXFu4Zevnygfcycje2ALGzqGoytuVgkGMf5m1dQi9L71eqbKBjRdnjG3
1rKBv8dT/wyfkDk4N2sYX10kwVKnPbkIELl5AZOYosczIaEMeri1cTLieWWaGWNG+QrG6JoGufK+
4McQbOyLSeGbZh2H/uqtRoipRL4fGD/ChrfKqKiLDnIqOENePW9G+IZJzSCe2+SGkxRUdSkUwBY1
8Fi6NkNjgj3a3Y6+4oaa3AbeaReBszGMNtdLw80ow0G2ENSq/D2KWcWJc7JhbzbWFmgMEcmsCL4s
JbGfIJRZbwBRgcPyZU9CjH3NlhUXGL4zHkCMWXwg20mck53yNfHquaQM6zJ2sHZGEaEdYYkDuLs6
553PCv4FhpxmWco2wyZ0FXp8buSuJMlXppfSURS2MM7ifEqujtJMUPGzE9cOzD5/OhQuFvQDjPw9
zwMNaCMilY1pCiY4bczfcGuhVuATKDyKpQ7PFkPqxgU2GMacwW+QH3sXemniLia+c2f0fy4RQwfh
nPtS6qn2Wi7ggTeuAS0IGawfmGLLXk7Uv+X158eWj5ZpFnwZ5qZEAx7/EjDy7GbPaLAjgN/C6N/X
cMg1oCg+Xp2cFdODU+9UEerfOJ23lQESXiobKghkrnuHZET/PrLqe+KgsaMfqGUErMhHF4Rn94oU
kYk3S/KuJ/HJl+eUOjTT0V6lEnDyNyCJQPwBr2sRUMBLVjK3bClid0hYPE1ltkdP6Zf4I+uiJjBM
8DjiRbgQEA94aNdNITQhn6koLwE2Ked8ZPc1itx8JT/S/Uwo/ZJZPrUOHCpG+Vy8bThn00phtQco
WD2xHoMCeM3I5h3J+ZXlJ1ivUAAL4s9ECU/zB1Ku8E7F+A1rHNNKsRPlQr2oOvvrtvsn2FEyJx0b
C1Brhza6gKBFETpoRYzvNRd7wx9aktiZx7UnqWfe1l2HmzCLiMKwMIWlPBHi8oPnDMPH3U4y/hHm
dyBMTG5KBMxBb77NoyUz6GU8/30R8vUtijoZQxtLG1SDo9A5QUfGk0H0sVvFFGEoGulEowl7Tusl
jBHSnjLJatqiuNkpbhWUZpFRUEjL3gfxuCRfFeNNDiBsBstajlmvsXQUd9rA7ZsuaGyl0ALrnN9A
fl6lwVTPLPfFqredt51Mir7kT+ShSYL6wgdpsweF3NvPPALKZu5eONmakcckEcCFQuwscK1eev++
wU2TNJGxvgjVMV7MLY+0XlhOCtvgPjOgXonOeouZp1WfvCMnA4CzAz9pWv411xWflf0KoUuVbyoX
yobFFcu+0+HanIVXr9AKUQGXdt0juPpm+CfVEUueeMi5RCFFqd5NEQ58WTyMWTztGV/d8iAl0cEP
YojValk69ljmYFQluhY09SGtaecu8eF0/VQtHSZj1bI7Ssq6a3gqMiKEwGkQXgE+9qp7fnkbJPvv
ibNIGrtNpjoPrKEEIdDDpoIVW1i711ROdSiZqL4NCjlmj9FEv+vmT4DgnfZSzJG0CO4v2qtX4tOr
zrM6bNj2Tytuv3fbVzXr+oZrSN4rvcQ3lQ9VIj4hV8JeVjICoumVqzF6Eo3jEhMbuglyjMa6mdCZ
ZPkCkjFpkF74MMm5rUzxDFQtfhfb1sZ1gy2aKJdaHu76ChgS3aF0BVz9yy1lzJSTVfK6PDGN27vw
gWsNol4pYLKF36SRZgwOMzpRMQv8o7DjsIhoBDU4lDMpOvikQUuDbOCL4GtaPWuGfkOCkj6QIom3
wySEK6ylG7qtSqtWeDCenW5bH1z9+LFgkHMC0A6dtDt5cYQUbgb/MywA+Ke/EhhD334k6Kbq96Yu
vtbzx5wbIwqKgtb3+LMSswXNa+Yck+ChyNCtWSLNJlN5bfeI2pNjwB6QRVD2vom47IsS+kG8aWdf
1hxTdI0jGXEWdBPWWv6o/yYJqj4qZNyuGJNpTejnPck/HWCvEUmls6ibPOWptt/QhFxkUSFULPWZ
fG5TtrOOtme23dLV0YVWZeZ+tn0P3VaD5I0FQ/sCC5ccxpN0Wm2izhDnuoZdhn6eVzUOzca3SWYu
lsEZ+Y8optRMl3CV/96dZw8hgAZmBH5fKzAAUL4oYbMhYVPMAgbG4v8q7JT3B0rZZZF2oCD3AT0X
V2s18C0aK/0mgkF9JcMsiuTyu975LaCjwCGcMqiwzTj6ZoiTO3EqbCJf8KSZPBNF9fwXH/+EfFHJ
F6lpJLb4HTlCuEUf/nlUMcb0gcaRg1ggpxfS4irlFUSQQogzGK3DGzEX7RgK2WMQAKabz4G/Yqey
bzLrHT7ywWX3yUMhV9dMBZigVO2IMg84lNjgL5yLae+IMTKHZFs66Vx48pdI0oj7rVOwD311rtic
yGk2F0oS3SaDFh1CeExk2DF7xmDwA91eRbHFsUfaU34OLNvspiwcTjgUM0Mes58hXFmD0kzxF+fv
CHAfVUYgKOixF+i+D8GzRaFWE2N3wHcg2SwFe98AOpQl8Qy+rAEHHvlDfUbUORhM2F5C4cj7lz64
z1OZPwwwMkTneAfAi1jp07IbiB/zSSxZJIseM0qhp6DoobF2F3hyGgKAFWqANJx0xIQKMQxyrFJi
2vkVcSw6dkm+5h+/JwVAoqXGz2msd05DyNLvSG4sfpy9SY8HUKgrpVSc/qz3f3hfAXxKq75jtzQP
akoxoEUEAl00J15xFqL3JTVqaw77yYn6plmiXNig1Fr2WHZX5sWh47wr3vnOTsMhVoYcVwri1BSb
IZFTRGATsQx16gvqTFTqCkS9AdG0Ve6EY0WlaoTepYszNjufezv9iJafxjVTVvNkbykxzbbPK1nn
ShfWC63kqhWlCO7FEbdrxTevDqAWQ2rBpYo2GuE/CXiTKsONiOnfaft+xgR1KYZSf9n8mOzFBT8u
Ia5K3wsF0EMwwAkP1tvEb+VKwyGNyveikO9Yc/dTStrEi5OeI8J6wo5suNxp2PFrXfQbDxyIYpxl
+aiLjvAkVjl1YKPkLeSIK6q3yDm3zKAFfFRKq3g/PnYXTW6CMtOBVsVWFWH9LwVmSKhbuinBg0dx
j3N6D/MM3Yd88UFFFkdpY8AZThUU5Dg024I6wZNsBTX1iSmEN9BXcyUULY5kZUEPWIdnqkkWk6MF
bZgKrJnETOUZ5OJFPgYBBJp1f71OF6uxFV1alNKQpk+yNyz7MbNToGY/JGg/uH3ZATUYe+G+f0Gg
ZcoG10EUut9bkivEXIUDJU/5IfnAtvou/N6NVEGxAvo3gFhleMMkXkF6TmFac3OcUYmEg34bd+Mu
0xrNlqoDwNm2/TeQLUXF7t4xXpVMBy+W52BQIAmyVVFEoqYbTMJEZTaltAMNPwSb1x65C+DJEmEt
l5VeIjMO2z4bETNNE49ae6bPLwm5YlVwy/enmcZo0rfcAVNb6E9lezwqNxkrhFGstDLZeezI6wHU
Ne5KvWcowsVylR2G43+BTUmN6k9+aceFsUmlqOD6VYfqXeyTQ4rtTWSxz5G3nk/FbszF28zs4HWU
tJKhv4vEZqDbWPAikgqMj3CNyAOc5YqZdkDWdBhry6Flx49pqyqA11gtU830p02mq1VEUMP7kZaM
lHXLNV4HnZ+EeApOzFCXWiRXZkyv9uiP+v9nxCpuZ085HP5SVatb4xTuoKIWShOVx2Vllzekhjtv
3Q+UcV9EZA8NNJkpesfzG82Y2huXE8kTfD+1Kk/oIn9isRT0V5XKHeeNTEKlc8s7sRK6f0bO3bn+
gPaFB4sFJlq00tBBMgyRgIZCb3FCVlm63xC5gMsoZjWGwVNXQ/KHij9xzuXdIVvbIdjNRqHRAEK/
Vy3o7z4sXdWVLlBaAsigJ4siluvESbyuY9tlPze228DLGBHiHqvPf5H4+uQhtBMowGn+j6OGgJCn
ZPjHgoL6xVfkQWUEeZUccBrHJ2bIX4Up1PjHGGvhbbRErVQeq/2jBAEZn+APF1x4f+7k/ddvgYcz
p3zho5CwZJTxwTg8kWhyiXtCv8X5yKHlD0xhHG+SSLPZ31+876aoU58MxKPhfL7NxYtzu1656coo
kW/hqkqia0OtC6rrJw4Bo4I2bRqgrE1LprPi3ygrLrRG7lgzylzAy4fGeOsU3FKm1zK8Mxgdq2cP
J0wwmkOnb2t59Fr9lkHSfVeomVZ/z0ceBau8PV0VuMnTRnxfOw5wug1KSXFKDDbgDbP9GgeZSNZJ
BvH9JyRj6+G6H+qL4/XqUOEm3jtX9+JsEGb7Qs3qvTnqnT0u/cW/1NdiKUD/hGYPzelsljlBg9KX
NCTJjF22hWlcVSwlklv4/FhCaVmgPUeFML+kW3RMqhkRXD/5vkOucirzofMU9KFQhroyzTT4flaH
7E0oLe3s2SfDXhRD9wqZah2zy3jnWVEyfdZqwnKefKtkw+ym60H2pupaff+z+qnR+ag9t+ahbzqm
E4T99yBV5WzoAUcpahGzqYxcfoz6XW78TXeOkElhsCgWL1xcvsaVUV6gnHBMB+53IQEsmJKBioL+
E0JPMmKr6oUcnz/LtibH/vA7cCNQGgfutxZjf87nr7Etx1MhZ4Jy0FQZk8otakLZ3JeXy9fWBxGJ
9Fw4u8o3dtxn+aTP2OlJFqFihfDeCXcahMjbHHf4GQXJKLZwzgCNptw07ZtY8ro7yExLh970oCs1
zB8DozVDpkg+rSG5uNZqdWMWKa99aluIVUWjLXXrFLP+im4kqf2lCwfoow3AK4XTTqXKKooW5hKh
10ieesr8Wxxs8g8ci7LYSISjbCvme33NNOr2dilUy5TlDB7oXFsY8hbGuaNe2O7DE51lRAdJyFEl
KgYdocbMIVBI/o+1ReTuc93jqhmO86AevhiPXBUYRgZ3DmVDaEyQoYI0OcFIsjBuhIwMgSG4X/JG
+DGFabz1rZb0Gjakl9tiG+N/AlLWushpRsly4UJDZbZ9jEwAlIymOa4kYTYv/7Vklj3671tWdqj+
IQcxqspDzPPkTHKEgSTP1PDJouBSZhIe/AQo5ROszbSB6qbWTSHUQMBLs4NHltUlqKY3XE9ER9+F
54Uvsv4lEuhv9ligwo0kc/DHgUY+fM6Qy5uFqJklmw2Ut4TOEye5AijzhWpQs3x4KnCLAZRsIGJy
ap0ed1Z/5KeMg67ivW0JukU+5FCUYyAACkfF9QnsjxcsW+EIppG2BCeA9NFCvhhQK3Vgv8uBTDhT
4DaZNcKYnZDFIxr4cMeyGMQXDWtp9RkNZl2EXLxmJB8/ZUIgGj6BbxN0EnFieEbr8sVp3Bn9lTij
Te66GGLhTeyuNhUkHTQceVd2uwKsA6ytq6my7urYlb+rLABfEmEiivtu3fcKud2Ieu1ciF08YTJP
DPwD+Z+znJOq2+WZvWXvd7ndBkvEXslyIXsPNo9EYIUc7gDLXJzc6QOKt2Mclj6P3aMCgAsyX2Bv
F+sZBJY9W6WRxm5w0W5o9bYVk4OnxFvG+kN6dL64id3D3Vh9fjyQQB0hXJU3dXab3p+Ch6ITqZ9C
Uk/Zsn/32vtip5jk0Hw0MfFEkWE4g0VqipD337ppuUyFqnZhz76To+X0rtxlKNdFufLCRPb6MPFj
Nb1CvcROtmtb/FL8O4KoX3dMvDJbw/J/9Jy0UzCaqbUd1+Gd9CjiZ7hsFVdz/GXSEV4QIZPo3+Yo
oe7SqhNib4kFemyiC4EP5vRMomY3eFEFopPiUzu4w3kflx2xT70Z58/fpLa+p/4Cr0W3cq515j/I
HPUgAGb2keyGYJXK27EYDpn1/JLvxSl4aCP5lMLBQLa+AqsvJ9AFjnfNEvR1VLW/BeSjZDyQFZCQ
5qAW+GnBpjucjd+XpRBUYJ7UDpvCLePwRdRqQbLkvsk4G8fWQfOuCjGupYQU0Ok5pBuQk/7EjkIr
ZHgGexzLlB0ooG4P94ia8I5PO59Q8/KYK9FtSF52xCVwYKoFcYPLF2yiCpUoXG8sHLlH8yrhGI9F
F9qUgD7Qe7+vqOtE+RSyNjtI4fgXK6ZDQ4EqoNi4EMATepb7JMZcaUZQ9dFCN2/b+9VwYkZ1rn+r
CDZyjd6ojlM0pgNJS1v+fYMFslpm67akbkirSbbheB89Supq9quPiMkBMvp52oGPeuVxPvW2WGka
E38nMMJ1hkRILCDvBX6LkN3owUGFcWTzg0RN8TgH0ee6R/6lgC2g/GaJssH1W/mflC4bUF5pOKjd
S7t21wlOdb22zNfl7mmVhrr2K3b+WBpcO0V/Q0JEE7saNOagynQCHOoYpTx9pGCi9tpRyhUMx/PK
/k7Xz9Hdk1ImdXPAXES+7Fus8IgH5zDscRSfA+hGmU34S/LJfkgHcu2b9nar7NswyH5vOeFQXgHc
eCnBSRiyGmSW541sF7nNZIlRmEpRgXk0dcP+fTAmkBY2tCmT5VFQ1lsztsfC4Cl7OPhTpnNBwkey
NQyh7/FZOTB45c7k+kJlwsypBHErk65iaXnjMtIQHoC1AC3LOcD3Ydn7xTyvPjVWs6e2dFwvQz9Y
CCZ63cmRtenhfMoIexQOidujCh1DKTQ93e1Id4zed89x/h9awyATpZ+bYB1wWEMciGRGuBKdymI1
WhaAYqZJEbtNPaK7EfnuzMhDY6bR3CHhzTXgC/kIHw7qE/+oJLX5jhP91VVTFxQZWlgVd2NYCxQu
s3DaxFxObteEhiZhvEYE9aZK0zuaQ3S/Gtylo39K506dUYdWatfanGB1ex31Y44kidDpVtYnCmdZ
1Agk6KkRf0nEH9hceg9kH4vcwGKw62dXLwk9vMkh6VFtO7BpQhkFFI6zXm501/5usQaJLKWEK4TE
GvI4YzlxxaStDghQpIrrkBGVtEg8U9a6fTBHgYkJQPGkAek5/8DNoZXMzApzhWI1iskCVEk6AIjt
IuxjRQnOicc3z7i33ISSlg7xjKFjy9tv8b6RRjmKMRR2m6TLipT6ZklhIjhtW2mO961fbvzbC132
7IbRjOII2Zx0pu1RK/XC6yB3YRYgesueMuP0JZr+8aTpR83u7qZwo070OyUwGUjI2UrnFIAShxWj
yyTV3zHcnGzYzz7qF44znnaOnJQqP86YZCnWZcPBX2uWJl6iM3z3tZYKLod8HDyz3+ljoZuO/U/E
UdbEKs5vqYfZXsNd7U5GcTDr4vlJh+jyc4QEzjtkFWZQJcVGwlaF5k7Hns/dNSGL+8RvMW6a308h
JcgGti8BFCMyFPIIRknLVjgddVhbmSiN9G5Ji0zZACw4ywqSgwkkna8tfcZKJ8Rlu1kdKNDYxgaQ
FR9KA8pdBr5k/sVC1lomVI1iSozVdtSd3Ck2T+QKMfL2TYg+h7YHboWq0kMxRf0Ne4x8Ub3z3CoN
/7VBYKfqhmpK+mAVSW2qF2ODE2uGLQEtrArMkGb/+7VFfJSBlHxSdClklEsJdV2H+wX3nrEdX/WI
QI5qql5ndlypgXqMzZ5QvZk7aD3VfJ7kYq4X6kL+PNGoM+vU9w9sS6KtYDaHoiU6C8qUsQKzILIR
hp8Lzb7wxYwQb3SkPuXF8P/47VtgVASXgxut1wwft1B59ji8SDpdUupmLVv2PQ41l3stt4fIOpL+
WmkOnerexOvFgp4eSvsZPZhkVZ/FJ3hl3OSDiDXpSDkdTK/OupTdR/ZxA4ER+cudI9SHQEq6k9+7
yTaPqAFc5Zf2fG2mKM+MHS46xcwGqstsHhEFGZuUjQnPfKKH5rTvnNEi+VSEscH5Miu/EWHYEjxp
fv3nYbJ7Rim/Uz/7RJPSCFmwBA56bqXKGHInS6zWKtHGs9EIkvPHaKiViaf6Mekc4vP2GXC2oVzC
7zK2dYrnWo+MlojaLw8hnpHUQBlAtPHkS2XGIOhA97PjxoCK6HfzrAX6H55GyCWIPdOSC5/V3R79
dwRJV1JRjE/p46SXkd268lesTUhKDMDNLBWIj11E3FULf/5PxEaxRLWPSWN/scJhLsbgWpoUnpvp
cQ3KqQ5YjPrjEXIQmNMYAeLxrEGFbXch279IPz36FyFBNzlR9uRnVzyB4DKh0noxTLIwzhBRp3W4
HvDwL2hHZOYQMJj/g4K2RqJ0BLOuYRTTxiW0ncDzY/8qM7SXnBWc5yZra9BcFnkFWDoB0Or4cmDA
vfSWhO5HX/IiW2Q1TVUHNszAGh8JghU9zH7yCkBaXiJOijd7UgsVQTUk0qCEvwzauK6z80TG8CO2
AmpBNzZ6kHJxIVUsjW5aOuTb0uOmjnRe0BpVuqzQpLexyIaFnexBWlErP7z7+4Ux/Qxxbjac0b+W
1GsmJXFj1WTZ1difOOEbFiYpmGZH20yFhY5XLiuZwOwl91ewaAbvfaZCbZ+OwZCCVDwmkOKXPWvd
XpTuOsYG/GAlynvOBbytEwWS2LZbmg1Fec6Uj5/YJr6PGpWnvCry2T+oT3SJp3YLj7OHn7jTe98B
/7Pcc7fUE6DNrUFm/Bm4ALkITvKICVgpzDOCxzXMW552h6qId/68QsOkJX7yFXdZYIcwMUDOOnaZ
d52qf6AWB10wFMed6q/t87kabRZH62hJRrn2EGxJxw15f0xZ3kRqhQFaZS/mSwRfahamemQ4xf1W
Ul6pnfMJZMPry8rVqmwenJAMeN76k7X/LBpIwVMTfyya1yOADX+WFQj4pyeXWFZteoN8ZdjMY6RR
KCvlxhH5OW5Uz5GuQ2ac0ZSJcdzICm39i1R+2+1DHLXkLvmpwwW1WTVEECzNm+giMpM5C/i5lnXs
Yjd52wsp0bMu5oYfjY2A2kbbZA/7QYzwx3Czpce0Rbu3jp6xCBcK+Pj+knWDZw3dRHG455lE/TFF
Y33efblwxrqUuFE8JyUQv+Wg6cKyBecWbDQoJS/BSlvQoeaV5EOxRW584S4qp7chlBN1yN8s6USI
PdhSBsUHLRLRCDlJdsJBrMqpWtx4v1nRd/cnfd4eqf50AhjhU4b1EiG/haPgI4sbyb4UC1xxSwO/
dWfjsKjM/eXXRkpgEE1Z+vsWWb0WLeaV6RuginoOlVMyW3JAsXQIY5/3usXSnPcX/Ubl7D1LQD34
Kqp8LsCxUOjQxK4hNCU1llhnNSBlEu7k5MPFUFTlpBZbIOo06ORC5iq51Wf2pYtVaC4m4Ojj3J5m
Lh3cdPhuKbCoOl9SnXMu3fEb3YwhzwewnzABdFYl3CLERXoJTOjAmamdkSsPr7wyUVsvlPgG5un/
B3FfdD/WJt39mEwe7RZv1LADxvgiiObhb3dvzRSXgYr6Gtyxsab8wvK62+Etd7NAhShSRWD0rT49
voQjp8DPzObtNXsd32i9WXKp89r06GhfSwxQRn00NFaGDSOhyEiwDDA5LgBDDd6t1WQhHqy7nbQi
7Wzgi/ovkq16+b+IQ1IdnZ8q3EeSPx3e6WfZrUAJ6mROOJUj3wHH7pw23IjlHHdaVXl3ygQ0q0kf
54j9Ke0iNdX9van8no9XrIhjPEg2QAESPuSoyYPQnWNrzkTbRialgeXsGuQjg1HXZt95JZV14ZJD
LEZdnAowqG+zEGxXTD3ul+yPYEMcYcfrWYpXQQhuJPuazWflMbDopw1n4QaqyAEz9fkmSMj2TBw4
+HXQe8XjltNGq4Sy0vDKmidjgjc/zdfn/pJxo3ubCVpFoO4SKMxKMSg18Ln8WD5juCBR7F2vGaSZ
iqRZo5xJ6Y+o+3ur4STWE3gGUHHyMVkXliBCQzbs6KS9RaGb3Hcm/tQPxehDrLwiS7a4z0rar4u0
TZ+npimItCRL/7p6P3EwynLkNgbWE/e80bMwszLZ9X7k8MKwj+99Nkd1xiMVIpkGQLoCju0XRnc6
VKBthkQYrLAIxBAvI4Gpby7zXRCvRyp8YM6lrbRC/FxR9P4EqEGHUcAiqWMgK7issKeSqGlTRPLO
yhAgQGFw78RnZARLDxG2qpWB3VW0a0oOe8wX6i9Z9cPUaB5x9E7Pj6tBsQSAgngrUNzsA1lz17SF
txzcHrB78ip+fHeahFNPeSBYxP8v9MxZA1d7SGlHhnTYZszTLRK/d3UDM/CYHUDTO1iU0fcVdwKp
wXcd6UqVrptAsVeHcEVWRv2i+yJ3SDfj6OBp8WX3KR3eegH5tPODbZXBoBZQkrUFIVocpo4EKH5r
Ad3UBUf4Qy/2h5/w1SbbEcFPHRPzgVqIrohlXS+FZqemhZFhhRXOpAakSYvZgaBCJ5P8nSKmeD7X
Sie2ro5Ka7FUqpMataUoznJEmzq8/jvAAS+ZzLruV3zTkKIF9iIacD77B4aRRT4eQ3teX3EfLSbT
JC4FWDkRtl4ov9wmL2+iODji0EQNEfrkbzCW4DPNaOQaQqWaABIx42Z0PyXSVQasefbCxF8Vytcw
89v0sQTn62FSmpTxPewu2td4mx9DICH//rYoRBUXRnj38uMUUM/pos2lxvJhN094O7mizGaIpGQT
aUswjnYdPdxDkWApUaVsc0CZfYYm8OFaWLY5XIlDLYcKtay371OyA8RUaOHac+JsXksqmxE/S3n5
OunMGS1PZAbV9fQWSjbIKVs/3A9RzrjaQuehDW0rwbN7+pt5jzgwpBMyMQ/ApbaS4qF2jXdR2i+e
Z8Dt65RVncYZvdUyNbC1B5zuXClUPUkf7EmTszeiAk2BLSl70MBWqRdf+E3FtlSRKfuMgYluUDUe
kh9OUqmzsZZgHhlNy4NLe6fp+L8GkgJj/48CPy6tZRSf1i+oscUNz9TgpK6+Ls0pBw7y7IwCW6Tp
m9pzzaHUt72PzpIKjaO5ZxoZC9ySMBibt2iwRdnq3Qb2K6AUjWOpTywXh8Uq3Tj1uKC+BB6CkbKg
EmH7pdu/W0aIAg/A0Mp0QiKmjBtBpwuYdSe7QLQEH1dAI8w3fpqmFsvhTiU/NERsiDC0onKNfNok
YJc9934St+bCewyFyEDuznVz0xY2e13HUKkQsit8U639eKojGkGG8+7/PjRnIMti5T+TjWDe6lYv
oNAa82LhHDKqy4l+2nzy8wzIRFikozMqUhybhuB8MuIpBN0E5gcYfEOWQxPpQhkYkP3KdD8nwC/k
hI3iLT4lUWZvyJcQkb6ntYdbToKpHLxfxoGpvJRm3rJGP82UNKamtfsqgL5fDga16V/pDYatmQ34
MemmCOAJiR9Ohq6nXKnO1CgVmHqgyzMa1Lecciaw85Gvd6FZPIVLhGtHN6dc8E3VjX1MVk4toiLD
kTgav+Vpvji/T44DxKUJvzC1Vit+Isadm7Tonhs2/nDwstnlMfsnZrt6pc3d2i+FYALX6OuImPNS
Mvgp9j6UKC8c4j0u4nQfdkw9Vcv7XOPF0yXS1bTTlNC+KkT/amwKxuQLM8TcXfng4pPvMbZijRbf
lg8/KTOoCTGLMdRwkg+sU4seldR/kf6aTBBq81A4UfZsuF2GEsM4LM7iuZG6uhwfqhLT1QwVm3ZN
c/GbLr1eHB/Gl/EHuS+UMHjqz0vRGFp2l8Kg6o9lc6aiRQ5GN1ncBYW7fm6lL1HWpMVWl6cn8ifQ
k5HVHw3ob7unq0kYK49sobe/ewI6OEHBt/mpRAymvUwE+MtTplK5X/QoNoF2NJwewi1OuukznNJ1
77LvdmLh/I6D/CX80qEWQhMSm08DvT6uPu6IyzbJKzyAB6h+2YIq3VvExFIqpSbXM6rWYt4ng1lX
2RDo51TAetX3XXZ1EEhpS7bhejVSvHoCL4SXo53Nr9fOrSjb8VK5lPsVWYcOjbme6QoZFuI1JwWR
birb6HUhDG2llrujFwZfThgFmfNq2CVk2razi03pIr/+DDQD9lgG7Jn7ArrrQEd3u77J58CZ/8Dg
6oz5ZiZljc1isaqxnvb2x6Qt1W3JolRZffhcUMxsEi/KSIMyI2V4RivU7G2N05x3seEic1vNe1nw
kFnkV3vdRy8teuiWm0w3pOm4sDqXMh5MF6GXKguC/eylj2QjStTMgUmmDN2pwlikjd85V3tg5koH
mjXwv3qWeZnfDe8brrcZsAHd5twOExpFMG3aJTXIQsFEDHCKbZCcxkdLvkfPDFd2FzJIwqfXOlQI
CTTjoS+q055x4PHZwPge2YiR/OXBCMAEslHcu/GrUTB7g+l7nI18akCuqPbtUBTqqCtnxNsTl61S
sBHYUP43ONAAd3vtztgJcOlJCCFLTeobmLy8y2gdXedUadT+ZglLYQTnCJNMlw6c3kz2Q9EpyXcJ
5SVonP6ekUJ4RFhOcK6G5QrSHLxPVAigagCcKvtw0smZ6rmAA6kEF8bEi23zTvPo/qAzf26SLE6o
rWFxiv9/PwCLHi/kZMOPXxNN985HFehFSjv2hH0u6GQaQZqgdEYkayocwGOCy9PhjPeZ7DW6zcpH
wtFC4dYJckUD/2306omjVz+Bzrg2pk/L0lx81E2y7Al6ZtRqedZUcKQIUrQvbcj9AVoAETNoh/Ha
9ON+SkM43i7prsrAsnrbmaAUCkOrhJP22LRIkPSpj/2msdFNWXd143a7qTMv6gCquCIYj71oLLtV
P6bBQhOpbpylHqKpvnipOlrhHRLQefNL4RaZM2Ojxny5up2GH2YutnMdpkcy9OgltJA15Unu5i0o
9rKLK1x72MX5sAvxL6uvO2rR8BOar3lrWxw81Tzn+fS9fycSv/A4xRV2L+Fb6HkozdbDLC5U+5OL
5hesJ8nmc1zS4wN/MTQn6IhxlI/7Wfb/59IBUXhgaFpyhK/qeWP7V9zhNHlGnau4hx1ODwnKgSJ4
JhAladcsmSB+CR2MbvhwFiHxKKagAQiINOotKrN2TS0mCQd2DQd2CxboRetE+B8qn0sVq+vMhHmc
xg9lXzcKJgXc5JyMRIQshnvxmV+ZXgPYRtX5hchk0AmDbWY73tOFTLgj1IFOxT66dHBWCEIWugqk
UclxdTHh9AwRbylG9nJn1Dmexa+eyWGF3DP7gXh9hSF3vY7NBj0aCGZwBp69jHrXq8trW3ITumf5
tLt/l/CmzenvyOrjx+iEGIw/w5PBsCy8uSVR9sf9TiIoXkrlPukYQqoIPdK4Dy7ogUvA4TPJMUn1
55E4AXUrN8+33HXIbZV9BAM5lju+GfuNQp6B6ZDErrLAxTXzTaKpSt2ANQdWOVtOiDt1lbrzzhPu
L5eecXMh7ofucSY5CDm0UFNx3bGxH917/Cn2G+qXTTJ5jb57LJPfCgyTYPP92zzO2+2JjCSxkR6w
hfg9L0in3tRtezvwAu3n97wkAuSrHI68o333EWfL3JE3IIEJMkmWbMJG1xuSV5RPTAcgbAbewSYo
KiQqE+aKFdbuQ7IVORhvMxz2SoDFAuUrpNkGgPp0GlVOtfc87zbRn+aB0xrVbE1H+EoUBTS882At
2GfeTxYUQ+WrbfbZGLWVKFbsv8nFEAWZ8HJPGKG8dvD9cpY63lTVD8ejpUbsEEkRGn67x6aguxlV
UEwJQAZk2LsC2IKC4sFo4XBH68XdzoLx35LGWRFvtrmhXdWyKaq1rBShTcak5hYB+U6rBC94DM5V
HpjLmzUdXmRmgdJnKpfO6UTwkpqW4AVZgcaP3/TxTWc1M2ybpolysMqMhWQ6XFInveH92h/ccbC8
a7CetY5PcoyCm1ZIXDBF0tAL0J10GS1Yc+C3YOeikcGsqANeEP3an8lGh0HMgfidaFtJ7wMKg1Nk
PC681K87GFd4myEFUCQrmtxre0qChbVBFIN4lpD9FOTTVnMySHL3o5U5fLXoVVuxb5LwcHI/S8CF
I1TeDldOoASOnwr3GgnkQ2Ro+rNWGPFGNqaMP/dm3tLBISxCVvJTxxCqJygf38AfpehZOBqIS5w5
p9IfUFR59prDh8B+u842CNbAZRSZGFzLJBNC3cpexDSoZe60TeA4yhn3WEDsBvD8lVPShEgwiWZx
iqKqTuDLu8QuHy67mx8GXQoY4OzEhu8zzmmhMrIiI6LQcz9a1MVPAaPBox9/N5JJkczATauO73Pj
murZY5TBVJCTnPHsT64KF4M+HkzsqWABxg2NZ1oAD1q47zUNyA1UYgBvfUosCrSBLpPbJXAzMG79
O/ieykcSOINv0rwJ9ZE92zvK11zOI3U3FIQAqjMdJwO3RvhdIV8xlVzpss66ZuRaIc0VvzpfReBq
bc2pIk/srqLf61S2YHjyR9mmEO0s6Ljm8dRj3CGagm5OARpSb7nrZrh61VGwV5OwxSGn9C7h27/E
bU9KEUeqxc3e5uEmyhEb1SDKwtV35KQT8HO9AAcg3qKYLyieUqj0jFVSoHqN13Pecrc4mQ8leUqv
4E17aEpu5mthRWISA/r35R8FYbdVnuAGYlfDoqh6tuKCazZal2xPnEaD5jydXRLm5Yf0F93jXv3q
qx3FCOcGDPSj13YqC9crHFqDeERdA+TtY/EvRKAzYHGb6le5Rje5vZ5b+I2kfYXMohA3exTl5kac
BAYU2ne3VhMPQ5x1PoA7prdrSYIHtvU4CeQ2m1LIKCJCVtqPcT3fMRDsxB0YuJjtUsLTgmXMqpFA
KWeYMwOZJZTHWhUCmRx5twchx0nhqkv3slbrB5ke4YtQ06DxNAfEAZKCDmpetC5PHTY5ZE5ffKn2
/yL0uXWiulA3+oDMtdOUOI2c7/qNk0SrW8vaZonNpd+3eSQqFE7ZrI5G+YVhSvF+h5X4nLTucOiZ
AjDGRbIbrC1pG5WesHk5Z2tsJcEI3Vd+iOJN7RBnNnuqWnivzPynJI2InAM1rT62uIczkeTAFZVK
5+FOOLaPMMLVPcTsHG7/a/F6Wa9DO5nEE+3V5uvfmoneuQhpkJnZEIPuVXdoEe3xFDyDfG0/4ajP
0ZG45Kt2EcBw+6PyW5+xZ6anHmnGunhn6/J6aApB/VCFquQPUjQ8i+7f11JOJkYIjoeBu/8NUvzR
9CK6P/MoC/W4CmEgkEB7FAYc8SphGlE/cqn6awsImnmyKfbssCYbwQBxJhx7T8HSYFrk/OHN1E49
+13PIy+KH4AJaglMR2Vj1jB+2Xas7mmFXw+n2YozEIdKHHipY7IsqWyd98Bf/wTnk842H3Uj9Weq
aenAWPSYOkcGJAmMydU/N4Bi9OCnEyJw+GmyDMnuQ5V6AsT1y9cXUTlamNh00prjIDF/KDSECaFW
+G5SfvbefXfODicwEGKAAcm1alQlXyEO9kZoYBI0UVHpLadoMk4AnFaa96B1vF5767uurqGceagX
94Wa6jo3gLQ1+Gkv/KsDtWlRuSu0KKASjF9T3XEgPb7OTjKZF1nqo6PFUjvrZF1lb9Q6ULUjAIJq
a5DwBtMkWuduU/e2jBdV3ryR93DW7LDMkoM0y3BfXZhxWXIMbbfovKD8q1iZ4ZBr6NU+9z2TtRqV
JvJlg6Q+UA4JrZry80+Yc6v9I39ZJXPfssF4zxr+596w05OuLvIHWgiTTbVq3tJyCFMFmN3A9pwI
vFTTX5aRszx0+aF7Uvfb0wI+/+sTUTkFtpJT2Qq/kHHs3aRqyixlaGyTdQmpGvK2QAanHgvidIMz
ZiJdk0Pyh5Z/snHBaESYdzIbh+pSLtAKcQsCG92mJaCrpB5bDbq6VVcnRTS4zUqZIOPzF5dOgsiZ
mYkp49urBUSb2YcDq3mUUnkJSGSnpuyQZi9J/PnHcIysJAmVRdRqcjUCKDcW45cwct4bZqpgYbH6
xlRkTeHl7lSGQHwqThETDiRWufiVZ2h33ags4eNZDAkFSKjIWPggvA7VvYNeEaofps3pO9+O/qbu
4AAQVefq93PSMbRqLbC2+z7InWyLOFVEAo2H0fdQuxnEtnp4/+MXhVnu9sBxzxyczOft40pU+rcf
UdYBYAjDQYLVfAKErqyKRnRqpjTkWnOXxcixzEBOGG7bOQPUydpjLu/SHR2wz73uSvDUJdFsbaka
BCNzaLrAgxCkgqTYOIQ5IlikHb4CgjnaIRFY5EEwKsnR0ZG5zbKcJ2ujz/pbZ827vFpjHjhwmsyy
vQn8nODL7mjtw6s5tydI89uNz9j9t00nsfGAxezqIKIuR89nWJqxyT2wNk8qACAzK5ZqvOo8zSba
qarJu/W+5+DujbAmAPFJaLFHXS2YQxsnjmPj/0lzbyllP2hUU1zbxN1L+9hMbgAVkdUVPmjG5wbj
PdP0RaGpXbBNWz2I/n3FZEfvWwsTxttlrct7sjkLmLTeBD9jAY7xDWgO4BvDKpZUqihgrljvS8fP
C8KfwuWAD+F00qagatx3kt9gQRGo7SwFQUSJhrm3FwUH7suo5GxlD5CMv3AaXE+mH/ED1rvhTa8H
/1CsYeoAbza19AADC7oqp0bTeiaBa3xt76EeDkCkVn88fiUSqDi9nI8B4dKlLtwxX5iW2i4asIbD
dHvsVzkdaY0wsXlG4Vge/0GHxmFZae75JXjK8ED0S3HraSZqCAT3O129JlKubD0RB415bJ0lwv7/
KngeFbFbkD8znTeKsBXugggzieEBz3A+CjvbSKenOgjQpoJVxXGgjPM7Wcxddr7pr8r5hWZnV3Yy
uwghvdu2zOEyC7mxjLWjYrImU5UEA4OuFCioNbbSRfRAHHQHtyqvaHnp9Zyzjga1N9yjgUMeC+lQ
grNvFQpDPsAXclpa8yER8YgIuO7LLZOkF43j5pl0kwL7zAuGCOdhINJrjkJK01NzHYV+ceh8vqed
OQcmy2bspnBVq8qAq70b1P8Upp0n/rdVRjS/FXPra/95/ReqBMfruv2e9y3C/YxLm3AImDwflfNv
iUAQcyNvQJStqpTB9pHpt0CbpuNAg5kegiFt+NSKUt/mvRAPIC3tasGezKPIFOqOSX3qLR7kgHTI
mXYBZlUIkGBzUUFqERQl/sLZF0fJvD97KPB8wPcOzzdj+lXAUKN0+mWIWPIG5dKfMB3DcFUG50Wd
zioxUtYjLqH6dYjvjxpR9Q8kYVwhFP7SzG4dMXYnS82NOHwaOuHII3UiuI4cAiPwHkxNLKuz0/6E
llvKJP8TGSivYWLZDHHBIxVFeTcKv3+KmLQtjLDSWkFnFOTzWJ9XtjEo5QkfOVNr0IY1Co1PVAFf
tjY+tEzoiZd/bS+I+9Cuq7SoYWHWklJOTNjrqv7O/VklO/YYfzKPcuZ5sCjoL+9Tku4mZU4Z2sUR
mTfEJo2dSiyMZrpev5Gw7suehjcGH9gGj0DAkkERW4Ko5FluMtMyN+NVT3j/DY2iLQyLcZ7I5M35
ojXeVtQ6f4O6lrI6DhyUjRG5pUAqNn9BVehFQs2t+u+IoumaTTWUkE/JXb8DUZ9XTUgPwy4273iS
JqceCGjMXcBCHns59b2BrCLSVkdEQOU4nHCGB86oxycBwCQvSZH2XCavCgOmKhJT3u37xaQ1QPzt
+f8GnISCGhZRDTF1fa+k10EJmtTIHvsPP9+zGyzDvBIprlcfqYkNBJsgeX6uQZJVd92yRWQQTtnk
uzH2WKNVemBH2j1QHYYp6qJqZGK7Na76pcKBiFXpe+noIqh9+Hw01fsrjpSRNQpSB9etgoeqBoV3
nobSjfFfaYGDN3mqj6UDVp4BSY8athoj2Z43zE7g3ZV/w66jGlwf7+Pue7dF8QdkbuZK/pw0ftsb
nGgm9QK4vxxdn4Gn9qoxBTW4iKlJ/7Plbw74IDnRCHJ0Tqtm0EbVzZs1sSuJpyvNM/RPqgvFJHDZ
6cJdN47eKlCy9DCEnUfjaaOZbZlYp7GyOJuhL7aRLtbEMKc3v2u+HI2RLjHGjunTi/zdKNx1tbzQ
AK5zogrbjx6CaLHSqiid8CUqUd4gclgNLlOEv4TToBPQpMU7SvnYDjRgP2ps3IC8uS3n+JpSZOqA
32q/K1gvRK4GqyOT8688dqDX9g8i8M4rQT5l5OTLzx23DTPq5+kgB2r+ClY0nwUZxJuF+DTPlnMr
+V/qkSmDWps2NjTdPy1XLOfeADcfswBKGHav7Y4exOwdHrCwm5GDzlA8emDLegtuE9so54swBy4Q
YZpwTDDS5lLBCxfelqN4ervXBGvEnWIPer0qoJrdkZG5PnvKJw8m8RMl8K1F7rNkfWHYFyLBnLEt
Zk6zYVLoY8mtBfkTxLQIT7shNBadT8RV2OSRPaHNVjhFwPCyfxe58uT6zouh8CfLDFSavMrzHCQa
txqXYmw8BYudXhowIbg09r3rCZNPlDkEOFRoGQQsT1g/zsx0ch/Hms0QZPpfPm2Gzh7XohcioBOO
Fcio1B79mq8YMkWGBw5dIipZ5eljruUhy09d+kvaJRMoGn4bHIDXu42yEemlWbChpMW6U9bwW92W
IjDB1Ab8Wxtwkikx/p37/WAh/HNigxwFSEv3CmK06MeeLiGMN2jJiKyt3ox6D1BHMHiUl7dB4svR
rr/3Iw4Zyw4sJnbr3H4hffP68wUINWNWmoCebDUa4VKVMRH2HC/oAZQz6ZjvJNdt1xqmAn0EO1x+
xU54rlypElm2HypIp1/KX/NO93PvWEw+0akNeoMFOOa+S06so2fV/qSBZRhmww+cz2t0CeftswFc
YmVpIDuRvSzAa2W9SpGva1BxurpmX00GOEHqmRSt4i5QNZ25TrvfB/XfF/s/2Q+MbdlJbjh6C1mF
XvrS8iCJDdkbMoqADIjKsMtTbz3iFMizDMxFsv+Ap8s9zZxAnb5P5RoCKHS6r2/z0jQeYBJL2wwC
xB9ggubNgSyAjzSrXMW2S6RcBHAtAsB8++/737QgzSBJeZ6af+FUbDk8cU2apIq+i2axRVhF+Z2B
ddPlVvkJWi83fybofd4oTyDpRd/RdDQn9vtdBibaPOpIHHuLCc37ofMTZuiMG1sFlp7Xamb/QrNA
NCw4ggHhSyh2ilO7Bhy7FsrPuVYSKPXaXiWSIJrFfoUMN6+Nei+80QqXn0Jbr2IsUSBtrRqDDZy4
KRlpN+UOiJh/Twa5D+t7hRJLH7oirWxf5l2uZEQmVyjtGplGpVE+maOgeYXIES+iqNP5JU/HO/zO
DYznhDMtwJstqw8Yl3VK/olApwdTrNGmog48+2wRlNTiuV/CwnBhZRm3gUanV+OmB3Pri79/bsv1
KjSuxZsgJloEmHxHB37qFONlc//J0/iZjF+/gSSDlY9hV+c4vTzhpEgLj4umK9WbUGFOC+4bmxeg
DkYVGd7856YI2+YU19SNSnqeaSlnvFXSVhinUuenZ3Ul7DioNOVsMB4ysspDgPP0hdM4wS0VPQNx
w3X/5sE1INWmwosofDU4FSNCiMxl0sXQMz53QkDPXpJNOI11BMkPEhR6vNEHEa7oKra9nWTJhv+X
saPJ65Onz0u2I/n8MEAaCxVrO7nYwG0usYr4EZuBlSLjbqrL5L3H27mwgJCekvqcYzNGB8D6AE9e
1ZPQ1TaQAk4QC6XqacNHiMQt0nvpHHjFOtj3Wq0e2Xv8kI4zMg7pGsI6IZwFsx7/SVKctpYKwNN9
TTDFKLu1doAhxhsFPZmwj8c1WwbV8V8pw9oXcgaXDVxU2TATQ43k5coKl0151ZtigRLdU+D3IC82
kLt01wv6FWsAJE2rIei0SYDq2RLubUAKWyzci1/UjIdFf31chfmzfoCrJkc1XIOxMSHEdnUD+ANb
BC1l7vsML8g7ObOEZKmL0Qns+IvKmA+e559AvCWEWHu2xqhSBmo2HBHPtLvJvJEgSJoj6VXfdF8G
z71YIhtTkcnW4WiAVlin4ATD1mCZlK4VDeycPZcH/QMMc+eOpN+kGVphC6xFOsxNoI4hyYqrghtZ
tLK/ri2xxeR7QMrQvbrTlEMmIpgKKcgL4gkO/7XOCLzVmjg4mnNaVpV0M0wSTWh/yLbnZgduYiSc
7B5lr5IPIQdITERTDGudmcrouALHGe2M4zg9wUnveBzZYAlVoXaDUqPp4dG2dLNb84/kWdTY+M1Y
Zgi6rbB/dZ3hDhigjppcxBxYGKHrATTSKDaDPVXojPLa05JoNVebZHQ/XPLKI9ovPMgo7qkpvcMK
NfpcCrDI4IN0mAxSisqd6T3Oo6Uwh85zmWMZPAhtriWhyI4AxtMmjcB25vl7vxntYZ/d515WpovU
Y8F3XB40TO19I0FGxbFFh4gR8oWS7oz8yGSbqcUmKWNXFivyhct0vW5f6UdkrFFlJVdX1SmbxEwq
Jbm1DzcvYSCgWAQIBiEZ9ixRejyShQY+7JdYq6NhZVAIgbDc05P+ictvY4jNBBXhdtbRao/PV9qv
yOeVYC5E5HYicmkp2xG49qyVXNjv8PlNtx1FFinXyaxzqrRpTbFVbF9Xy2oT1zVS7Dc26Hwvn9J1
9/5EzGCX0HrE5fuA4AzroK19ssm7+ZMYfhCPHaKjgS64MJxmFEpAi102R+LVglkovBp2MJoaYaUT
KIwO9l2SQ3g2MVjNPF1X+65KxYr/jbeS/o135EEE66mxL75XAWbhMZ4GXRsky9t5nNAmMLwGUpjd
HtoovSnoluC26UOdriVSsgvMMFwwqNRSfVAhBtPSHTMcapL82iPq4uUugsSsD8E1vGwqzRNr5/i7
ksG8Mh9d8iuYAsSvb9A7RsXzBENzIKmlj8T3JcHYI9XYwan8pCI5qVFTm5a/LuVrPItFtk/bd6Hc
uShfFHEdsdJYBrTBZk8j00B8Jj5r5Ga6gqHRF1lLwt1MFzPITZOFDTOm1T8qp73KB2YBs0pQfbW1
qlorzOOCu/BHr0l1XEBf19XdEeMJxJEfetOtOU1GF1V/a7Bjlhauap9ILjsqztqjyGKtt/z6XBy0
VNL4el5I0rOOUKUqhPniMxoCo4gu2He4UiQj0jPOKsZeepqu0LhPC0yLAIfBXIC3soTURWYQgUVA
VOh/iLRfyRD/5GB5GGhK6DPE41CyYjjPvgRhAv/70pi87e1o6vHfbEotje5AQ3W1idwAEVEgsB4i
JO/NqKGePzZQvyjTD4MCNqvPlVQ6j1Iv0DTzB1GKEIg07gXuEHZzQpfC7W+m+ZSSOz5l0XAB/kmr
Sd22jXYsT1t41I9yvXg8BX5Enb3wkiOQ8wwZhlaYbHNS+5uVg91kLZF/Du+end4WmDNW0qwvYYyl
yLO1JsjG7quO6Wk7Wdu6C/u1Nx115DtFb5+MpUdljwi0te3P0cFS4TI04cZo1XBTsmx28gm1IYVU
y+bbjH7gBI1ihuqWlAgcuig4iFOi79/mIG0ms4kgsCyFZEChO6iOcUlEorlvsTgQUAgztjBfGSbL
SdNx7YMntPbsVuZb1WPcJd5J7I+4Z+2Z+FZu2MMjwnW1GwixqFYXDAefEC/bPIEsHrjxYlCFR3Ee
Ns8e/9JMQwG7L8lzMBaZml+t1nyPw76lrXHCwl2kfKnTnHUQM5h4ItQSVvHY4AChFVvOUKgStLFF
KMj6H/p7bEKXOvQQXM0ZsZXh9wJEtlMYsiZtRyEuBD6xhxhiIoUojUhxCOx0Q5A1o2o7Cz6nQBiV
CGRRWhuvwBIWJoXrq1ralK7jBbJMAM+3Iw8+NGcInQVDao6q08TW5Tscgdb3PxRA6sAFrVNwSGn8
GB6L/81qCWhPXLlH+EA1dSfo4Ya9a+x3VKs0/4AJM4aoJ4jgfeOMsDHXOfgfBVU6Xav0ab5O7pMH
i/gBrPYg9HF/ildw7MrsVyucUqErNwils7j8/K6Zimou53pzH177iowlrLiVR1khiN7iGP6FPHwY
4H0Gws2v1BP2bbzpWzn/wWCFWAf7fYpZfCU3XEa2KGUdRp/XMeEiXnBFJ/bfxaEYdkrnLc3dkaNH
ronXjiiQNZkzERAhCMMJS75FMcKJ6omklWEokIuwa9LVA8uYGkuV5NgmotFtj+QDnk/QxFAbqI9H
cLWiC3/lWA886iOOQvLIbteAE37Cq1j1s4Xq99LDF6AgImmWPDS6GA8ofXg2LexwrKSmGlxUVbm3
48M3yrEw9gAV8gAf3t7udflSHu6aPbFSIqF71lZPE55hXhBlEy1DprRCbPJETMlr3RiP1lrNJS8u
HYFjfEmX7ccgVTFpxikl/6pHn6cCqkuwZbdok6PImXNmcGCaUCqv3WfClPKf59QSOeeoFJdP5GIV
wXGuUexE36sykWjW2l6mVyILLUfITzhiuIZlfcWW5XNvxWYPuJvYhxz1fJ8wc+sGzE0SaXfL4Hxb
8abv8Scy1d0NX43gokupM/z7JA7479rdW986YtElO1kvnhoZv+3Q2AEWQsdgwZDmO+kINF3dDTKy
98FTaqsdWylxVS7PHdKFb3HtwFicx7rf7s0MLLi2vwO/XKm80pJcfKmkHcNnqRdrBAVhA2EGThUN
1UFRJoMb8IAkB+9Y3ktNsDaohmrrkooQNahh2qBLqlD8K+fFXNCWFyztLjbOBvWcbyhhbB7q5xKm
WwtKeVAqV6UkatMuEPSkPMpV/YwxKvwXYh9XawskElsy+DmxZ+lM2DzDg+EkNlQNtpBJPZPZ1SuX
UXjPCQoEjcBwM0UxecD4wH/ESFgPoSi+jVE/ps4286oemk+vfyT7AE32Z2CXwnD0h7ZYwPLnFPDu
KtjKXMM1gtQ0KFJr61kYVGagVcO3YFVL5myzbsvO3sCOBBfwVdI+03QRNCB2G/8Y4qREdcwyiuFH
estP5eIx780s/pGTN9efLWg3oAT4/UI6pTdO17H6IVl6Q4xMUrveldvyFJWwvTcEqfmf6RJ2/QvL
To3iY95GcqdCVRyFBLFAyoltYAHRNUPHYI1XLNDLp7JDMk2/f98SD/ny24LrreLDkOAxJ+1TVZr/
BsZZ9JQr7V+3XQ/Ob0F80r6YWhCTvrP+pmpmCdJsXP/H/Z17CPGahmXZFwOsC7ww+FE6V31gpKOo
ZSq64j6B9wHvWP5CAA+fSuULv8wfN/kPAAWZwi9TQy+00Bker/XoBrjGHOwjHSLpPkKdDzzWovfe
Itx4pbHXL1i4xCzzVWt5Dzp1BEOrtK+sNVgxnGOy5cc2U+p3ANozr37/2edAZ8PfURep73gJ+Qcz
sOfd35H76gsghHxDN4Hc1eCZw0giphO5fyhBaV3NkS8XOAxj9XmPa0wOmMyVy37gcdv1uB5rcsu0
Pw+wvQwLE4NJ5MGyUMoYJDO/P24xe7D7OXuMJVxwz8rqfUZrbDmjGiZKqXRVrbi6xq1LgBDGMNVZ
CNKgD6VPIv0fkcUyLw/ifcMV3oEPSmqg1mw1dX3Z715/LNbTmkbUQYVA5jSWxk32wov3iH5Of6rZ
78QD96TOgrVnELoODojlC/b7zvEsnXjH6tA1k9X4V9nja/pKIibScAmIP8SwylKkIEKCt1UKhePq
d7HSf2PAf7Rb1ZcLKAEYWCx9MQTu5+ZB6s58S+0Ra4O6AIWqy92iTSfXm4Wm/gkCxsNe91t1bhRv
DXfzQgdXajD4iGolfXIWxJlvW/rHa29zJnvwbZ0k6psPYmi5M99PmZmpruCcdKr4ft3DpGUwIAeT
iUBHdUUiCreykw3S/mEm8KT/AF+VC19h9/En1oOqiyTRUbsNxYnWt5fV7Qaf1yxarLtvckoBICtQ
LvTB2zaLhqzrvM9DqtlSx24bsDcJkROtg8TWJL/CtsyP99j5MKR5X/uXZKS937lEKQ9HjFQM8OR+
+da5mRZklaiMMFQw68kBcduvTUh2azlezu32Wv6bw6r2jnFVcKoeY3TukN+AV5afBNBlYT8+vOKu
v5KMz6OGKlgazESQkq/oLlf0sSIhnJU4wfUYhqWIujAX12l7UTtL2wdCVe9BLozt26E4RYqTHtWW
Zj3/7JUzimRHbn8Az4StLY+ueVozEDCJXGJEeQi/YumLLoRp85PRIrBch4ZIPP2TTl3JF8YraM42
XemUiru0qPu2LnV+xlED2g7vk8RTJ/bb9aNB1Jzj627iv+gbuljFHcNc8hSWYdt2+/1T19bU0Hd6
3zGpZkx2l1Hp7t9NNQaVZBqTGCMIoHpVsbH+aVZT+xOl9jrwGJJR1yPp/c2PW8QR//BXOhW+POHH
bcVS8ZUkNyzerbuoiXzhEmBA9WbK7JeFMSVY6ZN+InfJTgCryJEBt86Zpw8K6ErcPA/fOEuPt5he
ol3JysZ/cIbqv+r3R1iZbVB9eolrDfDI3Y0Noia82Gfx4IaR04w8onC9MbQanNHNROzuhUSvpjYA
FZmsS6FniLtOpo7mr2Rqu9/DMxgT5agvTyMVA6+LDy2ztcW3oEs8ybeU4twIO41Zdpn9jN7JDy75
KUQAumpDnpCZK6U9VmswTo82Mr1mBxd9kIDth5tUxKPf1nioCBq8oN7ssEJeju7O0UePIfuGksej
9oTQ/GNSdfGeLsOfvxKP315SdgzUt385002Dxii0qLy+Ic1mvH0icQXZGgauqD3hHAVJU+gSPd9u
YfNro4eUpfEVYsT16mtfVXvNPgVLeopNw7ExAdzeg4f3tzP4fgeHtwE8OMZoDibSTsV4+ndks5p8
OxVo322NYRCoAs3f2N5Da6oiZr/HGe5ZH8vJkhZ/w9ZI5G7JWh1yjInOf71rTNjsiOJYrUXiU702
KGS3n88JrFmang4UT3nfA5RuELxyySKmEikCXemiu0O1RqX7E9ve6VAIuSlrK0Cedd0nyMd1oXdT
FI2zKhLQ4TLYLl5YaoTlgj2NkmNWe8cLsLnueLl1zEp/D6ctzkWiVDGJNrICSNAynadHTKdtJzZq
QJVGF2aYe2KozPsVxkq9OCi/OPQBDh7fmbxG05/ljxK6g0TSDht/tR2Ble8MzLXxwFPxfVbB4PJJ
Cvh/3RRCYXfwL7oe3ac9hXh2l1RWAI5IVBCPJxwMI1Q29NPXWLkzx6R6cQvFTyx0yQ/8FbpDn7ws
s8L7p5DrWCyh8FjF3ErgiO6zunQoRxKZiI6EICUFEp/42w9yaPIuqVB2OiyXHrDOaSQNMLYNOXo4
6sFoOfgA+WJpAdgMpKg8iNVYX3e0AiTr1OOlATF2SV5EuO3P4d7DMC5yMOelIp7mz9yrPaA3CcUT
ex0xQ5cl5lbhNj+ZDY30oWr8YzFJgWFesrhZ5LMt1shopg7hBPwxEwrH95xUTfIFaEfSTkpuwwk0
LY4h4ogbUZ8LzIWGxyxpgWLM7qfRab6t37BRo3nq0mVSxpBvhQfrx5z9z7TN7sVFeiWn7eA+aSTu
inq4jn+Zrjib8i9b6z3wELOO2tyVGBvvXHcpBSd4wZYnhJ0J/SjvR0XHKm5vaAJj4KqpuMEz419a
2fvDV+2KKL81Sb96nf1IosgQBHZ7MJmzrpjckO2GAOuWRYhraCA3Z0E+FONqbimIZEKco+gWMuIh
B/4yHGNG7ou6u5Hq8HzJxed/gjZ5ICmO2PZOK1gwcZmx/arG9fC4cZuFghPTNPNzqbeWVvl7idle
YSkM6u+GNRblElkIZuhWYykqvuI+HyJHmuj7RXCqxwoSvctOS8A0RIk52yu2q3z61XB0GKEDFD6B
WO1K8hNW/oIj2DEHXi+7eTDk9XmQ0esEGPiEpJFVZrb5ksiXuiiUVIMlZDCmt5nQX+d2SHEKwcbO
Wj/CqLGB77RZXOE4HGAIPVWT5izEbwHm0JeTzOSv0lISzASD18oDPyMK5sEwfvmnUTWC4F+cox6M
ZfTPPQaXk1yH2viQZ+ZXRD5aXeY/fwuh57rqZ2BlykjrEOpEvHrnagA2m7D0Xejg/dW1CMn5a9L9
BK2hsxSaqQD7PFH24vOihDRDdmj+ODmtA8CDawu+iXebMjzbuf9WaCGrQX8vptdeclQHuvhqWRcG
dDPlkfWuzz7PjGExdJpt194s9/PufVsjGjqtSwEmjDqv0nLi2rKJngmmh51ojD1oYPGwwN2nRSUB
/FknkCjJdYuIHu//BkudpE5esaBazhr5ZEUNDB1rA3zpz8h6wRngm2ahSs1NQspC2NG+h09Dqc/v
ipgWaHReE2pISKUbiS663Q83h/6GnNw5+TukvrWDSJ18HzwPjYBhnyWHL/4DFKL2mCxiFpRcRgW7
lJTH9gw5IRteXWLmLI+yekl0flaia6fHwnHWO+FXsH48OkMPMVp8ZBh+S556BBzW3RldbN6rszdI
37B/UcZPc9xwQdIYDF7hTEQ2MsrHazORPFlWy3L7nJdov7kAMkmsmtFNpECp7TpB61djXdwXwO6W
b1yfIKj6IO8DaTghWhuEDUqfarGjIcPRxZtxGracdTfZCRVppuzUxl7tNVj59uwuf8lyLvDE0qAN
7iHXSGnBnQBSfrXJCbFiSOFQpxXpaxcTpUMUD/4lIyEVL6AfdPOlpc23HL9Ylm2dGMaMF4p5I57S
MbHCdYQDc48q3lolwk95QXqSns+FLwf+q+V0N4UOwn26kngyCFAD59xr7i8OvjZeZ9EomCGtTgub
gu1NOeUsCVhXGaDSaWLvnCIoq84QvGpHpq3Ytuu4cppF8YJkBjajTKxXmo8wMWEJzpqST2oEemjp
9dm5xSBHikdMywGfqsJirI+a7hUAOBEgcoh81AC6LSDaZu7MhWifY4nQzu1DyzB/Mn7IJ2Ij2EbB
R5Om0kvm0rHSVHd2G7dHWc6sCLtHNg5g5Eqe4YLHxSWyfzUbc34faAzHJyvHsbK0jNgL5hUNc8Wh
Zj58m8NyTfHyrbQsXxno8NCNVPjBYYGWrUb8nV8CWUZ1mDjB9P3SVEKHL09c2iuFi9nvcIrkPCTH
8xM06fCnKaRW73ntKI9VUE/CZucQY2DAHE7VLdXOTeEDUq+e4mWvZs8mmtoLTzAjxhB1c05tzqsO
SjYZfP53wIHUVd1XyqU2aQiGqsSCOIxSybeG8BeHiT0f5w8PoljweKjVt5J1SwjvQpZqoJvXDRWS
nui9l0nMEm4pAXi6W+9+CR4LVIf5IPTkQF076jFZ23AAiQULTJ9/itLD8p395bxeQFhlo43Fu7sa
rIV6zTTllCyzpEAmENKt96d/vag2518b1nnSsVd7/AxhE2q8u71+oxrwsTJszf3cHPUut1V1v0lI
cc4HEjQLSxQzIgG0tFSfsEKkGuHUypH6vIsDDON6pjTVxe8weI9ASTSBjV5XeYbcxUjlxTpy3aHF
+e67GF2m5FM2lwwpbkxn4SOBou/eMhbPixj6FKc4Z6ZexyGGoVqbJZwXZgrUYmMX1eiJoNrz2U7n
mZy4nLvX5SmXMfmh8CC1HxtG7TxlRGcklUhqgPzhY5Svy2T3PgTfg+1YmRnndYaG93d6nCNKFgt4
r2Go0bv6+C2ik9KLGntLPh6C5NQzYqgWp3yVohJ/j9XbLSFdwPceLN0ryJ/KYceNZRwpZXXC6w1Y
EGv2H/+TONmOMNvuLDuDZycDQicob43pTqmtRC8bnk6JiqQ13wqmzVZFj1xnt1YLB4X1Ofo0QyH5
8Ekxk6rMSWKLBMLa706OhatP/hXkTC81QnK+jaY6YZTtLnpa0zLGyANrMmjc+awEOZ5Pvkbwu3Cq
dNDFp0lNtHyKhSaDGY9MqxULNuOl+ZHjLECzBgYiVVoi4ISe3vULkIikp71uTFCoioXvv3QaNhpg
GdPzRNjJ7e5F6JXua6baY9ttiMFJGZS2c7AcSTgYashWkDTqE+euicyHQoulQqqSUknadDWLgI1V
R98pDvTppDQVX/6EDsqNsYi/Lqu009USviYQhazkKqJxMhQsaRxunu8XCjY3wHLTS3a4BiWpy62Y
0qqpx/FbQoe+s5GJuEJ81hwlYUokHizuiEQd05NfErbgGUihC/U+KXqIsuAY1+WUiHYN2BqqPKKl
Qi3giPlt0LvTmcQExmSfQunL39hxinaJrkdnz4ePmzEwKgSweBIrCC4XXWFcujNyYgdEpl6GVuVx
g7sjdOvHnUbHxqY3BllmZElSIKSa3ErJWB69K8V5lkpR3s1GAN+yQaVD1ZwQGTQmhqNSWr3Ya/DB
hEXPz9UBaYYunlGxWdu+TOZQzT3UG1YrGGb7D6JDHVPDgTl1d5AEqDLDm59S8eLodIVFSQqDKZd6
Amz6fVUY3fgAO3+j5Ui9/9pCsXR7brSgF2qVcw0ZiZanLEvzF6VEyjY6cBfnjArP82zUd0072hpA
DSGF6J6U2a3e4QPsQK7wxvuutp+r2Wp4+FaKgcEKuyKPzRo+kqdbn75A2rmWxFfiE3bGlZ2VMPLz
rESbhe/bgspwlCbd8CSntIyBbK7scsr/ttw3FXX+Le7nCs+/caUu3GR6GgEz9p2MATD1UbTBsvgu
idl54hFDM8Yg6ZzALQKdwqavjFeXotNCBnKVX571XMo6hMvE1f5LfEDYYpD0qyaskxS5T22uHMZc
JgZKbLuxNmVRgFE1j52H5yOvJmm3R2GmzYvNfrCqAenB7u/ZNri+jPeISL61RWcnAmiH6dl2fKB7
/6qhdQeUItTNivlmIJn4xRQVNfLYUjGq7JL0qM17F/JXt2Bav+XuSWit1nDrQuv7o1EJbkg4yJaH
+at3b+Di+tKaTJw8zZinbsy4qn01ZI4XfWZq1nUquQ5nDWmRpADWzdz/0vXoHZdubk3018qLOlvA
Lv+rO5J82/sRE1wBQLePbxQdOLMwQORRHlrO+SQdE7MIvkK6xUy3TfGxM5bh1QfwchpIHylHRq4D
3fT+Z3wnqj++e4rt8XegCn6/rVaWXjeT8/F1rtKyj7jCx1zHyEame+2NEMej1mOy5s1mVgF47NEr
762AMRppxJ/tBcesm8JA34Ejy8MAH/1op4xR8WLUn3fEs5FJTRCNH3rEnlzPD7IY5NFZpTFvqM5j
WSGWW81CRn5jvaCr+puoK95v3BwdbULV9hoqQ++ewMunLPhbHLJ9nlLFq7/qDyAMJNdBA+t/EM4o
tBoFI3IUuGO1QqUEhGlNs8T5fcDOe2+TaYJtWKgwN0LTJjLr/Dk4KDVgkkhIP+NmiFKi3Esr6Hli
CqY6o3Yc+CwAhQv0YcSydq28R209TugBF5+033SYo2itGssi3DHZU8hyqVQVylxpN27e9sK8kKhS
lxP+xSEF+W7K6fds9AGbuXwOy9ow//ILozhPZxrt6Q/70rmf0FQ8qRF3x6GgJTyvEWFk8lRMDmVg
aK0oA7vHNxZCEcMiUytX9URX/9AvfV+mhHf94q0PDBPz4VNsSWepoR0zq2DTsYtb8jZjA55Tb73A
nSQg/iEAHQMb/lO80Nd6VcedYBVNnvRxLBKFDIaQRaydLB7+v/coNF8iMf6Hth567B+tlsDiujQB
qRJElhu9LrpsOqvSZfGNIQyOxS2Bsev0lOQOlJO96F476tohsubd7nVrIoOQ0Hge8+qihv7xwbwW
T3dYvTc9rnpwPA3srAm/ly/1gMT/EGXFg0nuk7/U7/oGrsM8p+3D19WdBzXaw4bNBqJ54GbUMh7W
TDyAJubTah2ly6QS/7ACBgHLei0GThKIXDa236aS7rJkxkoMPqwSG4Jv9BHmUsMOkrHhQb8PcHw4
q+jK+mRQy2vO3J0MTzXWyueYSA1+J4uIF6QVhvfhuMwAsd92LjtSOS5KWHXvrFU+bPtuPaBN59L2
2odYdaJnGRIloLPLKKRvLiCzqouXAmwztnCcEzenzcg96bGl1AfZ5qYxK7QGNEODVwMTYEpNR0zX
MpkZqzsu4jaj1wzQY58Atk9VlBSKpm7Aj3HlNDef2RPha3+DO6ukpLhUbi2C8LI4OJVpbQkixebT
gmOwVej0vXGmgBEL0rr3nstB6/tnXGS2SGYCqRNVFpJcoonUYBkOY/oWx5DLN4tD6cuUrEKUYdXg
6RBAhxrMCyTfanTnIJFWvns0iVibb/k+ysyENXpwq8bLYGbgjuArV9CZsHq9wZ++B2Y5cCWV3nVw
/kQLiB6WFiBKZlEOppremJIemdGuZOI7z5Ltz7582tuglR4TLhM+E2siY0dz+1gBn7nGu2AF0YRF
CCfRPjklIBgTM1ND1BhIpm5ePOrFMMM4+/BxA2lobiGlkdSeoFUEhreIXpfsiSVv2HuoSsEgvTBo
qqxZwaS9X/tT2RkzfcjpolbQOwpNSw3oKhep6DsXNdVBH5IGujs6KyOdSSaxbhNnK8qN6G19+LXB
PTB/4nXvdTN1F1Ne/Qwo0tZ1Zpbuyin2TKGmF3M+K3TFE54TTZLEMST9PDZQk59GnF4BVaNt4Ncy
FW9rH/XPYvnWZdeK8ZmpI5kp153OK1aq/pWYiElGX1YEOzAR4alSwd0fEJGK0uMyWkEkFVk3KeYH
CEddjewZT+s3zBIB7iqHUEM68RkL7PvcWJQoqK37y2PMG1MeWUYSXv1yXWs3S3JXODoPAT6o85Yu
vqAGkLRkxcL2N+bh1JPmnTX/ioRjouqloAI9NXld5P6bhvTCS34gv7H4jJ7TFnTifuAnvBL9tH2I
HSisNN+0dCeDGe2i+jl9ZqlB6XBMo21FTUZwCGw5nGJGnAadZ/cqdf2YW324PTtVnXXhu1oTsE7d
bxfXszNxIfgJzpBxtiOmMuJlCyTo/7PHQonGxn+gNQA0uDMMZ0LjD+ggGpI8ptkORMiqVPMB8nHM
uRdsB5cAuk9YlHVBE5YFNC6GQB6Wvm3eTidnCr4/8AZwLj+eR24jpiIXm+kofoKx2iKTSQl5MyvD
WDJjkahX9csHUQogZ4UQelS3B3ybXEU1gzwvP0KXPybIXAl3Tu3qdJzy5XXoiuai2vjaEaKhcJyQ
Isz1aKuSkABZJaFcvRdiWyaKE67fa6Fb2MomD5Jfn9WCfPecPz9SDdRzOtHYaNI0lp/g9n8EOpUV
qFE+d7prGX8MQLm1KO3A4fZzGQOOdLgwMV/wJsioqrIfLnL9w06DBwsEHumY20ir2wi4BAI+DN+X
HC8eAq6g2a0xBM1Ih209FZqxDKGhxS/SvWeRcSF/9IHPmpPjWbjQSh2qHyAs5h8OGTkBaK77YTiO
8EKNeO0hU9kN9mBheUg3oxPbKDi6OXOd8Ogb1SbDFhD0JUnmvdF9nqQdH70i7pbcUo2NNNWqvMlt
1muVxXeLMZTEDYtBCKjXPs+Nnp3WNd5om1Ps/yy81k1CiOLv8md3UBLG0RkTcXE/PakMEp7mVfar
rSmpXQVje/3dTEulMB8RGL6dKS3zTHHUqq3TymPAX25JsvSHkDOqBWh7mEvb8xsbDdrM2mvcvwUN
VD06A4+75dkxBeXEycMf0s4SLfjecFwR/PxlfiZv+lecK6EUlVxVJ01pPnsS0kwthUfTVS+ce/XR
9dE3H7xm8ltba5qgDUj2cj/RBvqnJAx/7OyRPi6TLacDBBlx6fNWQmNTGBfdN1zSjpdH+7AOWYNL
vHSLgCxztzO3zp/OeOfOTmPqOzSETik7VMPrnn1uZT2qTMa92An5Iq6Lndsf7sRNYzt+r9p67EbM
Y9117+hv21BuQ7s+/dV5jWAiJif2o82/yIP8w/N7H9boIMyN8GFzSLLAH7rpMERCh8tU+uU+Qawh
oWGbYpglAbKSqTMkY9m3b8fmgw7vze8j0GYsMhxI2WlXis/SKw+P6zBfNWtWUT1yZQg65z3v7bh2
ea/QewbOGVgs3HBzWLQ3MMXfFPFl6Bm5+I0wtt/QYgLTH6zEDEaSQ1/wi0IgqpXuFPYzNoER2CwT
EQ1TjXVuRo7BR0gHFo0AKi2oxf2XdUyb7Ulv3rwnhMxCmA/Cafk0aDDtAgihRkdd4Pn89YTvjDR/
6qE6ir064JHxDzmpPoJEfAKdNjSVgDx+N6WLFdx/oXy++irAftphBdn4HfNSvAnSNA/s1RgwAQZL
mMF7lelfUUUTq5vVMERXuoDpc4OTigFi5PnUldcFf9diSDA8SPJoOOjtq7GJ6o9snMNUpYaCIa7D
CmN4RmAuW6vN/UTxR71BlMjMt/NTGnI6i/iSZXRphWfRCFQ/hji6mAZE5GU2DzH4mAbgpyZsjZ0Z
LbKAGE9zsb6kcEsg9AjxN2KLRGHCiN/zjl/KtxOSF2OmvZl0ykRxdzdfM4LwPyMcScp+6xMBOGK0
8sJ+ZI11wQIxiHyw5WAGRCIgsJQAjmUlEpw8/lUV7Si1W1qZ+9BugzSivdEqRxHKj9oLGUewV1l6
vodW5XJlG2uJlly7QR6jTAkctiw/Jd4WF73PAfphtW1UNFMkml5mW/8Wh0IR8HP5vHkbRPwYhqBT
iyCSqdpy0BRNxAXjnjI1cDDIqXW5G3KYKew68JqpMcPTQ6uGmHvkTAmo6CkbKTcEeTa6MnA0NlDl
oTQ7H41sgeU7fzb9Bx3Qg7fQDyzxJb4ceNgsP6hK018smbwaEr1E0efTDomPNUkIuOf6kcRsnK2B
vy3+7cs+szrk6GNV1MqGKjYnh7v7HPE2CHWr1lB95SbX3nJHuebKbOJYzOmUq+5bZX9N1z3nx/1E
sKgThXU8/vAFzOPlYXTQhN2WEYclFWVBySmOG2iz1A5M95x/hKZ5C0qM45WuoD1YT/avuhZze7gQ
U3Im9Yemj6vMIVQfddr3T5aClZ+J4G+IXoqizISNwK4jCRJ7JFoKwsq4ShZi+FtceUDwSR3k313X
2czzJLn0GVn9Pbq9DmlMexMXST+XUg5lh8gVLUtN4SflMAMQV6vS3k6C0n3xWInTpbPXzPD5Jp1j
HMBozxhp59EK8yaD3d6TzDvtpMtXyh1Lg3sJ0pO/aLHaU62UglYmz2W2w5z9IPzdEqiOeBwqsAhK
GgWIAAIa8URz/+Qv70RbaRPvTyEES1mUEp2uWDxGTNKsBAI5+kIqvEVKBsQ5luWtpyra6JCOmG9V
UkSY3MW6ZiP2zvfmjObJq8ZgSrkTKtvbhj+wHtrB5rt6xzNR4PMq3FHqGYQMR+7ViRGTvYjCe2/H
ud9BjE5NJSZU5446WWN1mZYpcyoJcv8pSnX1GUMCjltddkolOpvqC/XZRGCurpEASj9fCUfFSonV
mnPny3CN4etwYy8XYJGfCsAwU4fje/cUm0cJ1DsiUgNmS24bFoDpfoJq+S735q5xAoIYHrodd93F
bB+usEw1NmU/GgsC47dSd+Q3WfW1Lbe3PJhBZrRYpxYcSRhg8lEJGT8uXM1b2WalASJ9qDEl4ovx
ROVVWnEb6znmoNNEoNPi7NIFoAkVtWvrjGx+UgWmiArSY+kGy5heYTbiLJ/6DtqZa48CNVRJayCf
AAlwr1K3916ln7zAD0+mUIuDpYtX8HLwIuZC0h7PXJ0KX44hXOIhPTWieAZnrRSiHFE+roI557Q+
UwZbQaN6SfwpifjiY24nnRAVDLFKtj1YHCRHKg5wnbE=
`pragma protect end_protected
