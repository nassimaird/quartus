// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qNzEoZ6WFEK7Iy6jvlSM1xPJo7K6frVnsAoF7JqEiY/r9jSsVVUXDz54TCRX/W9H8fsP70lFrNAp
bs9/m7lAX0TPe2avVf+YIC7IMPznDPswe16dPW0RyZXEdQZvWEIKt6qN8EwmdgYbIaOkLzqN8dxJ
9NkeD/J44HWPqlZrou4kdWhVWtosNUB8TjxYr+MZoJazhBf1GthfINblI9e+EqXt9qw4q9+Czb31
GLq6OH6gNCcFn1Rel+xuhzxFsnJ+EiehvAP8ASSzhH56uvKbb+a9yWkzgKXuCPkt+q9bhRoJgXxX
bapDbKVRk4mSoR6fJfD/GQ4FkdiaSe6sofrUZg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7120)
OCrH1KfrhFzCdVQ60Vt4dRFLK5YC5n8Fgs9QxbsbNTC4A9pr2RxhXGi90qHKY4Hfefcwq596k2LT
cbzlyZ4XIg1hnQ2pT0xPdtXvqfFG1G2dxIUlNtf28I//el0jWx7ihf1UQyyBxYiAfiaEt95cqXkv
4Ap4jXgWRkfAkgTLEhcNP+235pCk5e8FD/K5NEG4ksoR/FC786Jscsnn4XLMJWv239M8HcRxGVDb
T9zQAan2bjja5z7aGEadiLdcMiM/mx0AoXF1K8lCThqag0rm+X1si29RTyJV412oHs7Mg83WTE74
/ZL+jMx5f+0pdFzYL769QrFUqJYrx5XCKTIRWWDFkIQHU2TXSN5AbL5p2GLz6WJHftfoGEs5TEOG
Vhc+QLTX61pYT/UMq4u2y3GGd5PddWk7Ng6fQULFqo0Xu69Hthk/mMxUMb66urzo52GCSF18djeS
jcvB5sTsr/E/mdRyruyRSeQq6Q1f/+i8f/8WRTgAgZBS8tA5hQXhT+raUWTPneSr4MQKs13aWBGl
klOlgTxoRlGxkm7ZX6/aRa/qEajQYvVzo+XWMI6egOpOPNhBxHa26TcGxB8Y6jP0VfBq6xZQWyVk
TFdz3rQemrZMV5isQJPvT+uAdqPtaSK7onIkeSqCR0HHoL8GWIpvSC3bmZiMt3QLonkUX+17XCHu
tdvNjmrkGDsvh2uXHzm0/dNxtKi/kNxydaK1Q1Rvc9Fy5Cvz+k7cOKAstE1hQveUH5MYFn1tYvcZ
T4jAkfZn7LaFaJHrmw6OaYaw4Niwd4NlVQMlk5YXsKjoiQTmkLDZn4yVByOtKQyxTRYFjD3kdQY7
VpiOP7D/tpd8IvUeu50j+QaHNTENYyZLNLwmGAXVuUfPNPzkhib7Fr/Qmd1c/NenTu50QHxV3T1e
MFlDNVidmPWO5EjrcdeHwAY8uS2lZhKxKfrOJ1N8bYeq3dJT3f3z4b3VkEJZ2NguGjn9Vc6OvTbI
mtusgcbG8XRCYamGN50UEAsdPVl2YGE/vL1t1eAwhi4IgPt/6jEDctHnyqzOK/3c9qoq+6KCVA0K
QrMbCE2AOA0Yx7xQlueEvm3lHmkJV1jnhSDLF7w7I7Pfm1RxSkL8WWaI1uxYlgV17ZRJ0SIbfzCp
neHtM/d49ypbOxLL6Bzn1p3LagwmPIvJ4ZJt9FFkeot3hUC5Nyua6sp/vE6g3PaQVp8s79I9AorT
VqaV0zSQrdWAeJcvFo3DQyGdc6yLsu72nl7sn5Ok503mu/7qRANSmUm02dVQ25q7R1WMwRVxE1Vv
OFCvr5ONuEV79RYxe6YJbFAHvy7Y6Vln6Rx/FsGUFfOaOV2IL18pbpx2+SyMu548FFOF8Wp/1oh7
epVQiAR3KPeL8PKOeYnyaZJ2PMjDFT7un+/ZHaUGmStCqJB722bPcEJP+TR68OYq83DNgL5WLHkp
EisgFPQxFeceqkek1hM6W7EISM1bGx2+npkM61YmKPdRUmfWHT5V8ViwzLtfpL9R+H9P3Ohd6ry2
N4Y4UUFTuklva6oi16vp3gOqFUHHCVSJGS1boPSITdNz8yZLOQRP2jZfeVTVdC6fb/EL0bJc8V7Y
D9raTVYnT9nDIHcbks2Tadi2ZowbU6k99M5bwYXvga32iv7M2IJgQExIpCh3Xodg+EvZRjgAzRcx
n7m5iuyiTeXZV7/w1f9UMjY38KglV6urudL7A4OXpjkHfMeJLxiXrfr+pbvCiqb2H+kwQvAKGt7x
z+AQ4O8TlSAjHKBzwwwJ4CsnmEGK2w2zexhZM+Bk9Pvg9kz3Gr2/lPjM3fOBmRNN1JlH2HwnzK9U
d7l2bdTBKZjzatMP1OtudUq2vXzHBZbPdrP/myRhd4g//QuIXwEVbBjVyM2R7AEuF5EFpT20zXjv
m0t+MLoLeS3w/Megaey96OM81iAnaZFh60yWplHL59vTNcRqn2jqV2J5NwoRStOqezWWqNFeFY7Z
O4REdfv2rJCFvA5zMiSWWfGDRfOVa9aH8dgiLX0Mubqbt6NePBnAcde1i8ePem+VPcLh7OHXKlAk
SJ9m0bs6dzU2Q9YdT7av33+3pgeb3bmJZZrnpasqVjXWo/fPBatsHkqj8/FjtgfsiZ4ISpiXWqtU
15/BgxM778Iffvmz2KRri0KeBTkPTh3zTdQjgf8kgOS3pke2iVpHQyu2ngKXKEAiIwlaSIj/qGve
xSXkT/ZHOPP1mbOH68U8elbd0Iz8r3wVNf0MsJCiVVkdVVX9b0WKjG81zfMbsofF0AhygrVi3vCn
IuvSltri/SV9KztUTPNaQdOJxdpOPPfiKkGHQ/xActSmW9Df4Y2ea5P+4qbIVnCT7hh/KSAsMwKe
uedjXuZdt56oDbU9XzzHl0asMYx3VO0CWI+5DcrrQX6Nx2zO8qpO4d9Rlg9ysh25UGuTl8DsXHq0
f7WIXjRbhsA7n0hTdxVCBGUHGQOUykc0zUTvqeguV4uKwzIoFsc7pcdaorcYvPaaLhzmWqfpvDP0
2z5Xh7cCenFCpQSZl1G/nYzl/Fw+9baCvR+zQs2k2OzO4VifFjqfY3mDiTwO3Gjgx60C7Xs0gUCm
sAbXtwvvJU2m1Y18ScZjH/bBXAp2FtzC00T6qLACwpePAyOlphJeZPSiFxbNQeikkb5dyhIRjCN7
i4Ld3dREHSRwU7T6DqEwW3U7RPwUdDiDGUbV+ESQ+4eR/swtiD2ijNdl5PdCAbcspMKyLFZd+Gav
52wLSMeLLkm0D+eOhiyrQCEz5Xkcryd92JlSF4g3QIy0rzkHlokszGlPNjP85upJCqP5Y7Usrpm1
RKfhs5W6Gkb96ajr4W4Epf6OJmeT9PxaSodbRR8l7XSLNZdiJwipwCEhHKL+iysPY3Uudz0wreaF
IR4zUxyEoUuwKfSxgnEMvvmqZbEntv9TV+UOcSdqx6LOeDsur5hKzxiBttiuaJdHgtVNDl93dZKe
RRivaoQ30TAVojitmU6mPK7q7QECFSGqbszOOaIDtovYzc/W5+0LiWGBkYUhkTKMsO82DUl5vHSW
cvdRMDVNTFFeYtMbIjst5fM58/P9DYsLK0NhgwQYWqPRuLDxHmOnvbEOekgY7pUNW3BBbyhC2sSP
lcP1WVvONmkgLr/AlyEt2aESg1FbnqcaXVD9Lo+aMUudccmaLfUQGZ8eKj6dw6+UpLKLD/dO6/GS
6k+1nH4YTkfvvJY8dsCQLmzhOKLSAU7gy+tIkYtsIfjpQHxf1PeEk4hH7oMnDgIMrhM2FoFhTH08
C/EUM6Kbc15vVKsp7LsIflHvtW0fjvzA2UIx9sKqVecsZ52enKKKSK7Slk9hNRryoDGCoPyOx9mm
S1pbG/VdTSGi5KTbJ+RId3sjwoBEaSQ5pJNWRPEMQgOMMjXRrZX0/jnDFlfPO79j+NSDZe77az1W
qKx7E+sceToNszewyjZVyUKC9FrQMPlbjZqny5hOZRGuif8tm7paRGM68JEuv6w16oUtUZSgc04x
iq/fRt59QKt4a4NXq7uuMBOWPmaF/FtmPP/QIAxTJu1ZJLYpp9MBQu+ojGPOcv1sAs4SF5IBwReT
o7jw26DIbTlqlcf1nspgWkpcks57X0va7xp3QdNZ3HJStWkNxqbE2W59yGjaqZlAHgSUWg5v2F27
QiHIAiT+MWKwAkPNCO4IJDQNFoc8QR7M6XfPWN5XXhk6GwdjreC0DfCkV9ttTwDTb143HNEk8Znq
9X+LgtPS1Io6jPrXNedpoJJITo+puUHt99dIJPIuRwJ/nWlgY0yPZzljwYM8I/WMrhpmb+dpxDI2
csI+vZkUUFag23q+5MfMbWCRjbeuluoAtNSnvbr6eaqHb5o/+JYL4y726zlIK4reVBg6hSwu8gsl
e08Yto8KtO8/lpsQH2OzHGK+DVWJ45KQw1jjBbmh9uhdLpapvUR+O5xZQxmjqFHkYY/jPOp7wpQl
C19YY/zO8x6Z4u6ZryYtEOrzVo4uVxIVKV8+YJoVr/sG7586DNpclSt7fZIHrvDL1XWlxmQq1iez
02m6pdqVmdDfLZwsSpRzQc1nHRmtJpfyhC5KSfiVeWO9a/ogcB1VHa4D0kKuJrHQtm6WRVGCScPv
q1f/WdbugJQdKrDlPIDvQjzZsCrO5eAGNkuvsC8zi6+y1bYjUMeZrMMYKpmyU7AnU72e8swBJP73
v0uNB2IFtJVXOLpCFMZ+77ecLEeEQrtzP2+2M8FR+2r/YJDcV1zCqNgTrDtZYTDdw01ikebx6OlF
4VEs6co6iCvYfeoXVuoKnR8D4oSbiIN7aCEFiTLvOzp8l/iDPT+8NRJjTsYEtWWru2AjgoPVX3iS
qHuQUSiPdmpOhbUnLnVIJ3ZxuViSUuwXownDZU0/8pFR8vQSQEjmF0PWltm6g/e3EiFlt32HaSn8
GrtWFZ/Iwi7LKi79gl1H1p2FSj3ofTPNWhbLg5/aizxhLlVvvPYO1iANrAq+Dhus+YiuvH8baYm2
tkgmtOmoUvRd7Of9k6XJZRW0GGcSxHCMo5WBCAzKn2OXd6rbYCZngLOSdXq2TG7dK9XTCy7XnNwh
IXqoHaHOtwDQL0EHhqkDvkTPENwyzYpzllaD9iO+/uZAZdXKUBpWjHcd/bZw+o+b3BL2cVHDnHSd
nObBUzQ20HGXahRj0GwWL9FIciyEg+RVPCrcXSf/uKUjbOu5gHkUyLDvV/jj5JnHckBKYzJGbFI3
LyFmjHUn7rd2ERFKT8r43OK7TH0gKKzsZxL/e/01zaPuR0xS6lHQfEepms9AjZ46DJTnlt3hiMWl
uLhLsVb1PmxKpBlx6fqz4MYJABEBjSs+r6bC2+Xxa5qwG/ki30OLM91rqDwVxpKfHUdd/3WLIqUO
FmWGFRn5IxJINiEiwGHipEP1lg3yyXKINb8pKRYjX0iBkZQd+WaGk0VQwSdvRyFF9CgEmEmfQDmI
3/RzxY0HhOZbxB6l2Sp3Urzoz0haxAIVlDxOqGHSB2CrEHf4/of+A3+DH1mRERF89/NRNq/O6sOS
ArzeX8+YqTHiJ7YcthA8xkMvAAr7PKq6/RTWnB+uG+sUJUidXfB/zWhWaVeV/xK74SGZGDa6ZdEP
yECy/raWpzLHFyjwCz11vw2ZkOUQ83mrOjpKlXDUUq15OlPz+In2oxUGUoYHo3s5G5Evs2tFc3Gs
SXSKDso76CFL4mbmcyX6JRJdWn2wq7Z1NI2E2P+kpL7RSD7lg4Dn3PaRFDgdaQQpYre9MaWzmRwS
Dn90Y/58ElHDcE83Np8UA1bZep/299iq3AvCaPasz5yYVp/fafB9XlfEwmftU77utHIy6m4d4MfK
V0W9GWYSHbxVkLmsny/X2njowDU5qn39zYMHfoMcpS8l9+ttR4aHe+YtiHwHt/wAkI6PZ3neAcLc
gS9eBuKMzWmwwQAmPWaV0zt+o+thd2WSaVxHiMsMMRHggOtQskiOfQP1hYzME1T5Fmo7QTPGSGPu
mL9lthFl+lFs/tCk3IpxvxFQ01dd8YisHqiqpZjPr/1YR/vitphT8ggTKUbGxL/TodebuVdMckf3
Y6GzCAmz2xbnzCd9nwXi9YgOatSO6XoorHutfrj4h6/sFoVOPGWBarzZ+1ne8Zc6Ikx6Pjdi0OF2
g7oM50nGFDpEYSasl3ej7VluybieRZgdGRWlvw4moyfTQAJbCurMhixxzJBBkxbnF2noM7DvKGYE
oeAz7fW6QT5U0ZvM4b6zc2OUTMnrvchweqcqcD5ZGek9/oRJhcPtds0WqjaRECygCPaHdr28+n3f
CthGeDz+wfKGj2PU73+2ceILfzbUTOUxFJKOTqJ2oHI+44ceCVOS2UrxjUvKxb/vAEw6EYIHH9C1
23Tyggo9omXEIjR2QPVgEscwrBkOxVr4jl+W0fLgVRjezquZRbaJB9cXvM8WjIRp8tvzXC2lKMat
bQoTNVtRSbX26eYXynoSlC1Flp19txa8iK17Qxs4VRrlnA31JobDFkW4n+aDknYpBUkSgrA19S40
U/s/s3F6KZ9LF6RyoiG8oQrog7KVw5kIuperSa3lTOm5TAvyaXAhlJImbEbHKBPU1WoCpdQos2xH
wqxTayPrjMo2tv5CovAGIqGi4JZDQCYoNFGKGNpGuAVIg8QozEtW/aGw9Pz7uJfRAed1Zw73d8aY
PR39OsT4gLHW+OiCJliBzUIiKTXECGvj7Hn3mTsnLkFO9JlDzJKrnyeM/qZ4GgSyD0mKGbnt0aN6
Qpgdu8euNG2/VyWUSlU03NhEw/QDlxVs2VqSKnoLS5zydXdwWJuOVt5JjODJySY2sjQt3Oanu4eZ
OyKGDqbpk58LpV5wJDNzTHzIK9+bAMD9svKcyO9j/57Y9MiXTwrKfrwVzlF7j7MtcPkob4skAl1Q
XzN5wzYh37isbwWIL3gaPA+ecsolYMGQG9exMuN/CKwFJQg1HeYfTWOXUdlZGhEVnaEETcKEPqD1
ke3dnAShERMDFcH8XLynZNP9ntxzlrX8jzMCbAkqBIQNWu3ETww9N/RgLt2JrBALvBgQKG+qAGVS
loGGQimwiivZTds0UU4owolHbriYtzL+ruqr1KyIjTvpvfeu3zmdnzV9EMOSIHus65/RBQKzEaGp
slf+xGiJoxQ+zVeHaVbq8KRvviI/4ImCtIYdNROBW3lWwtz7JHiFIt4NbsyV+bHDPi2nAkb4vKIn
LNT3G5om09DQDxVEVVnx7YizgmzsiMhv/0tji3CT7+ZlE4RkwPt41FQmkEV2LcqtzPgfi/+JOu+s
ljUqlIdgsLKp0eu6eb4YQyeaT3LCxtX3Gnab9+Jm6RUsHq4dZBtm8sI/averQrNWXcWYa6FK3wRV
YgcoGQtt0OzwfWgUGQ7o1VXFbl9XogNfBYIIxDScMOItI1d74xOWP2JB33lj3sWQ02bbdV1NzZvo
Ic+Zz79R/oJ2a4zX4HTtnfGejl1uxyFga5FWnGnQLBjvFvKhy6/05HdvUANK1fwd2dTKEj3S7Wdg
f5xCPnljGmIzjg56fF1gB+gwUKxI8q5PFneLd1bu8N3ATcyQlw3/BYa7n1+DhebD2r09h7fJ2yXv
R4S5ZZrFpqkzVHIIoPnwVj2ZSN4oS+DRJw79yJ4sKHC+C+vE9hInuHfGvKnHQNp6dkLM3DgaxIie
6A5DI9EQJdQr+1xI+ArmHFCRBjDTYaiENJpab+8oVEiKqiUl6KsczJ912VM04qYlEwNLCMjdZgKX
x/Fq/zoWfWVrwsfUK3zh0NPpaMAjnIM1/Gj7g05UZIHWXu2IOlBx1K8urCimjTWKf+Bi9DirfTta
a31TmlmKOljDkYwnC94XdnQ3TKEnyTbpilmVonGdjNCYAFP0rR0178RxH8mBs/I+4k/EdiXzBlft
IHfc0r4uAlEZdu1x4zj3Svd2qRQtQh9ykVB5tr7igZiF4o734qkL3AazOa8RytoXDpEg71T7R51S
8gL/oZOhxvKSSD4gM4aED5UA7CB8J0laocaLV1VhFAMKoEiEsSkyVtZgdkbbI0j72Xd7YUiPq7dl
fr+8e0/6q+oEr3Xf0GqE3l8fhNhdfPIPLpz8/A6bRSQgiVzjVm2Fj8nlIay5BcfuTeyDhvqfay6+
6WagR+TH5xL4PQCujCR3rMppUh3ruTLoelJP6ltASN1cVK3VF9SoQJLE02iwl9W/Vrc67OdB6cJ5
sXhnCmAIL4GZV+oAmQqaSXp3V3olA5AQNXTOWWxjDiyMqI+L/iG8D+brpTmf++oHbRV9uIyDYOyE
gtbwzeKEDjVfe4OX/ZgRxdbW1bBfTa64M4B2CtXSmGxh8Akf0k0cnN91BINeP8T62RiGp0EcULww
M3EPikbWVt3FOQ4UiyNqCfaZQ6E7sg0o4PgnJrybYHOyO9Td0kvddO3Q3wd38V0NrSycss/mmM7g
fYuI9xH+BbpvSGPOnOdH8iPVNVQtnlLcmyKrsppr0/0VyfjGkxbM2YMI9eSiAFncw9p1fkypoFCQ
2m05aU3pVGljZGjfwxMUhkpvs9kG8ohlxkVwTsjmo8OhUSL0T0ZHp7MkQy/EBGa9LKjQXX7Wh0d+
r69CE65TpcWSMocBStW2MsvZfLZJCP9lWO5sIMdlW9Ki8L4x3KCh5zaoOlR7GZZ0MatWfoYYcdGf
mTPp0KEscAW0Ur6YmbMDxgwrQAw42+5Hj9B3zpyKtLUNYlMnFhQXvj5dH7q5KkeINDg4w+6KbBAU
7N7q1xZ51RsMI7JyYLK2VudLBfIg1nRKC6I8SGb3N3tKCziqXTujkTXFOfOmcuRYWSc/8pUOLAyu
YAIf2XdGNiLsDxURmUeK4RBGmIknrFc9SXscv6JSqvmVvl5oJIDym4O6H5e1J0+kvl32LytSq7NZ
GpivJ8ruCyyVE5S4NNbzaBoJilWnOEslHf6MFZ187VAQKCtcCkP5juddPvL6YMmA98p0ftE49PXE
W2Z0+3K0NyWgx6j3cVC0JdP8k1QNlQQqoEJijzizxK/asjyxpV3V/El3DkdHlB/OrOEyOvMHXagF
u6UuuP9EOrIFmkRe4K4m56SQxFDFUpe2F6fHkSqWeH7UZpKQnNy5WnxsQ1ZSDTpmAcdHHFClt5wS
sGjAA01ZOTz4GymGLyVh7+m5RXeyTTcDifKRCKglvm3dlH3YqQIJ7FBqEjt90b3CZFKzDklNCNMY
g/yRN4Af7JebzTPOLpwsJUgKFIcIxylq5bczC2K/RUwKuV2Y63sNBBU36lov4Ta1hZLB4bWc8Kd2
QY/+nnTq8Cm2kygg8ltS/BZ7Pl4zcApiKexowgyqK9Rhk60ZwRtPX7ZlZhZxBZAtbKYvF6t+XDHB
qTHNM5NVqkDNofa8HM0U7lZi3PMGYG+dDx38NwX9R9KFCr6GOyK47OGDSbSd73PAj5EkqCU1EtJW
/XFE3mwMOJFS+80Ssu7OFQdML0nQelnVUblyajo/0D2onGwlD+kBfGQFkgVKRgsRJOE++Ghm2ra3
V2E6K7rSaVUT2tN6dkilnwqt986az441772eYlFKrSrtuJen76MvTMA9kSlPHhF7PpsJ2rkHkL+F
rLk0hWdrIFTm0EWUDZuTy6jQgUaEInc0kFSRCsrUEqST89oM+pXKIk04VDJ8oOZb2vVXjdt0xCXM
4Yn9XpJ+bfSdhv/QA70t1I1gys0FiVR0xMxRAS79A+NB+yx/q5FGqqz98BMsJsMIrua2CXhOlXmb
KtxvIT/6eNU2QJke8ehGBj8GOnmrqOMs3aL1UNlaSRuXky//kmi/v4zEHtq2OAmaJpSBts0V28B8
vNXm0/56FOfeZ7p3xwykl6qS5IDYwE3hCl7UEMGDJn0YpXO/YukYh4FT6+0yGkoAnjkFIaXF6Xmn
AEVzI5lWjBZjQn24TZ7n48IEy9mkrCxsfZ2GsWoAkDLjQW21KKoAuFmaB2unK8+0mR6kwXT5nYqz
78i9gMpPDER0d/2UbSALlKF+xoGzUcZEcNbkOE9CdXzZwWSfN1awi93Xl9NJCR8spRTfVQ==
`pragma protect end_protected
