// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
j6v/Pm5sUwVqlweYBxtOx6okFp95HVOFhYR5P7tQvf9lzKlrRUqrfWhDfvNKNj2rUhN4ReCObc2I
XT6dcnPc931Opa2MiIQfxMXW9vgGskQIFyXunwNWz7hH3MGjNJEQntetgpLIyf/ymbls+k245BCY
LrBspKOLt0/79/b+E7SAut5kY+ZpdUe7PpWgJV2lkA+mK1nk5fKaQD9KUJ5/3X813nYxVBu9+BRD
jFiVxd3a9RZ56Jcu8ymtRIpQLoBA6Cfc2Ht1nORhaj2XWQjJlT1VptTu8um18BdcUN85Z+lKn7Nv
wyoY22MPcxxUVXlnFeO5csd9pvfFLK0p3Bn4zw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5808)
SvuI3LaX3ydD82WBdR7vEYcpI/Z1ATHyNRiHv+tqtf0IReJS1Zx6qvt3HvGbSuwZfja4GdQDjCyK
ibXnIq05dT/GLK3DM7GkLH77JCPnuhYfEgwL+3DyDy0YqM1glo4QnVXjhCE94qsDWNlRJz71+yWW
EHOtUJlCTtI9WRaCoNbGkJh45bod091o4eBoPA107px2l/CvI7qDAU54+OyowIlYH0OiCeO9oIHe
CRW+sKRt/HlFfWriEZ7Kc5Sr3/S+c3o62Iiw6fsgKfSmfJtZ4glkxAXIc/x+yoWOnVw1mnJhZg9d
Tqj3ThdpOKoJLhrAfjUUUBfZwSQMXqAMR53r8TuX9kvTnuTWlIakQlZJ05YpVoCYzBbRuWbnxedp
9moYBXh7pNErKr4XPeXswSEEcHTTHysMeB2huDV0drLxmaz2z2tvVH6K+hQJ36JrIVftm41mjysZ
6/x2Th48AbiS3S42WvDZoWZY9CvEz6ssp40/9BiWolxf1VWxcWh2AXXojL0q9EXSn1MgAeSeYFfD
j1VEfxb7Dq2KMBWQsKdcu+DSAyg4Au4l8y4Vx1DKQX0bvnCFBLXBcRXNzD3eRVEfsHUmwHohdQPe
/dsVyzN43Lkjx/RpIKpaFCeu+uA9DW3UOseeG3OpNpb608HJsoAm2okBFj3DVUR7JcokvrFd9NXf
3K8bZiJsP5bzybo39sLnUtEqFVnINOYLGfgTDfyiffyHX8uK6FiMYTl9J6ioTnA4J6s6GEw6qEZS
L4Nb3S8w3o2arajuHHVAYNBiebWk/3Zu6rlz1HEsB9USG6bIhsaGVdmTbyNCUEVtKQBVxlAL5bZI
SjR1OsUZpC4nTfIpUvv7Q8GIXEUaGBr3nJizjWV43VIzOzaxsja9o+jcPckUJuFEASlHoRBb7/D6
fbsYSVbPmLwPFzHQshGaWFaqVOIitr2KE271C6nubcwXRoja3DBSRLN4HlY2X5kTfeAZX0AdmTkq
MTzEfRZhqMWvg4ZfIJG4UikKZ16rsP8/GH9rCyL16R/6pB1hUof+0yT+lEhD2WNjF17aQxIrASPl
AeisgZQ+60LEjbz5ILRDkRtOBV8LkTssvsI+kQNMY1ZJGfmQdn2V2YVl2VLAfginmA17ktssx02Y
yyY7mHQ2Yg1TgWija0Jeld3VO1miJE9gGiz9sB6rC1ktEH/IwuOtl5lxs8Fh45dy+C3CxdawdU4g
7MqXl33P//B5l01M11WQJ7xcGth5hzOXkJlWo37EiK5KqEgiFmAeYrxo4NoW77Mk285yyodXQByB
n7Rh+nvNLvzkmY34LevQKjXrLwwf8HmDe+8GYhuaYt/YFf+7EIwUaFmLcHidqjuNggScg+ziJCQP
ZFDxLC/can14x5Q18SgziCd5fQmTPnqB4lTBrYt7XWMDrKvj+b6LAcJ2nhbiiu4Imt2lmbcffAAq
eVR2mS86ZeCr0iYs1TQ/Gr5fDt6gswT/0Cnht3x7v4qWOSPj8ZHRMTxsjgGNYNZjWAmPn+GHgv7r
tbs4QEF4zwUKMgXhDpc4zIYM0S3qSaWhRLc1pMpeg+GwSBtGtOtbvwMGQ/fn1Q/rUIARJfvlc7q0
94NFOx9pKnQ2d3QsKzYLBEWb/1OYjBZUbsyRf81SGBtLy4rwDszEPhA6LNcu9REhiPXPwUCWvUqu
t/7gwG5PnjJRp3obrVrT5ntjEF711sLhp6tIpSQxnaPZ+YYKMagq61wEhX/iRLbmwg3xc8vf25u4
JxxVPC3FPe9VjmrvzPkrm/JjG6A4Lc8LnskmuEXFc1BI6AITkTm0ZSBrsaHAcqgmip2JWIS5ghTa
bllGEIweIDmVz7oe71r3z7DnVg+PuztBBci4Y4MENOY9Tci0MoQ54o8PlnYmgUw6OBPIZGoC6XdP
OahhJtv+p6OtrvimWtNzIfKAWh4NseTpxgTRv5WiGF3BRJaZ1b8z8LIt7oqRyEqGRB3cljZY77Sa
haQL0bCyRf0wquUWGTFc/SyIdw3PbW88WgTZOghxUc+eKqOXUyyL8ESefQiZ3XtkMExc85fKINWz
LR2TBrx6nQIFcrR8avrDnPG6Y7xEqO1mcwmt1dkx62yWrETokWmRkdBVDfx4ETktN+9kgbHC1w9Q
+RryM7wPgy18WCvJBGs0UUv6En4nAg2u3+UT+n6alz5B3nPFTtOg8GMvF0eDfGNhMDaMymeW5TT0
VeImdZgOV3CRBFBM62IFjgZ2xjR9PMr+iWE8b09PjrzvCSd4C5xM3hln3QJPs6tMmRXcauMeimnr
IZz8DJRqumCmGQ6d3k3KENzk6k6DiO7Yt/mDFpTxtlXY9eYjL+XWHNewAcOybx+KIV+URpLVaxe9
XLa2eiz9biKHf64m5lRwERsw+7GoTTsuFjHFv0U63nknZcinqvz+mCMFIs4sG8S+jPRdLmq0e94W
zf52taLMfv6mLHtuF19fahdWhps83S8kztkwaJmdJunm0CCfrHGUwYr1qIpME98Vzv/4HKtz7vGb
m75MSfDSABbjPrmSgnU4KikFZAtfpUUsoAAP6VZSYVwwDCq+SedyX2TdtHqfJkDlKcarQ8tWCXi2
nEJQfgK59e+S/zEIOH2t1giEX9ClKKbQcRXP4v1BgupKusYzRUX0FDJEjvmHrS/FAhyiweB3pTf2
RVuxXdr7WjQTBETIg3qkIzWJlXi53fi5IzdmZJ2gjDnSYqfiML/vRKhKe1zQzSsS8NLFKnyVztZY
px8EVrypRpvIquiAlOaZt9luypvxxgGqQAZWvWaxyvabwLXFaIRxM8A8EPggLflmemVi50yyJLMl
fIoBgE7UPU+LGaYjH1jNvmVwmkkvtViyj26PvqeHbCZcR/8gd3YMWYg+O313QqW8f3VD2Q779Am5
/Yut8wgjcIgfcloj2esWLGGmFi4OmUlIGbpq/8mHddpJxhx6XXv3YZNHoxJQ8rouPQpYz+Oni4xM
4jz3+5qhbUT7MSjX+MtzwkOyTM7ZBTWUC3UFMHKSrZD0cRBhfVh/iuSkHW5QcinMedMJgrIlmscl
WhFQ0YSS7BZl7/q2zDra+xsA+EFx2lf+19xRbxzVTZhzpNeP9kaGqqfrkRDXIdDgJDuY/7a/qDmj
Qc4N0gZUabugaqalTn/k1hhtKT/fWPEd2G34WsHyVQxRYRIMqJNod9CJLC2Hf7/qj5omvXvy8Ys9
4kFBeaSCK7SHFWqlfGNJ8/P8eAhx4T0uImzCjOmGNMy+od9M56oPoy6sD4dIAGzezYx6VD29IXOX
nLmNuQXkn7Wo47pmPZvy4EbmLoRD9IFeDjBrTABxGFGPZhXTeB8+u/XtlMSPalqAbWLVZi7KQe1g
6vm7NsIXlam78eGFI+tcEw44aQU2YJK8P+VVmvGpI2fGAs8ltsO8vo5TNW4YryoFtL180g+mAfZO
FnbM5BZQK1Yub0TKVCoaSoohiPTF6vlcI8SKf0B32FU6V1n+mwVx2d87mnRvtSO+kKTcyv6BMl07
U8Y/nwIYLQHtsgD1LjsAVODo1GjwBpItIKYHo3fM7pM9urYfu2cYScmBfJFYhw18cRhVVPZXYtpU
lymBYqbNYfGgiU1BxbkIuCjhXpCQIWKYCH5r6iQ8rPV8AB/qYnJYI3t6vziVLa/sNb/9PN4/oZaQ
jsD7f1M/VTQi1sVKOS5BLH0ZiRFTTq7OVU2zED8uI5f/YyUNi+TZxwtd9HeKei5e7Y5L3MLc8WFT
KXbE50EIse6uwyCvK5YazACc4BdPSEszWJcN5v+0TDGQxjmOhmGkW+Xaw7RNLnrQ9i6IvroyY0/M
ZmsdNc4GctaZTDjZjV7b8A8+xmatNgblYOzTsr1XxkEHKhrNAnyG01uY5TXA0NJGtD9FsaY+dRcs
N0wL1pb2w9MZlcQOe3b8lHOWo3JQIGiKXmcJh7e76nmxpt+Ts5wS4eDUACt9goRU9u7sHx2k1MmP
N3uggHb0aEme2v8dtFc1qnAgt++GVYAmgYQNgUN5w72g4/CiGOijGSfVixvKI7HBswaV23ypXzPz
8pyJ8sDj5puU4SshypvsVF59T0JgziCcTpg4S/iq8xwVHXzwyORhaQPr4RAF0C8y/EnZvwj1AHPe
BCZQU/mOlWjg8fz8WJr1XPSgtybayV401MTUMemROi2/DOhw9Yu8QIHenbydKxTZp4z/BxADNxMl
zjd8Nz6fGKAGjcVWeDK6YcuDO8tFFqq8mHfB2spoHBkYnawB8UHbK6TK/D0ZiOJ6061wcpNJ/7iG
eRCmU4ixuanhZeUggeQ/1rYGO5V7GPZZNLrxH2SQCoFdu0I3VacIBLxsTPa2WZgGsGoVkv4bmq+B
0BKX0O/SKfvdEGBs9c/t3lVfV7hofDpHILglOIRc1r89z1Sydjb0PUdOjQ/8v3VbHeyXbiiN73Bf
0CyiqjFYnTQGTHBQtvB2vCHFHq6cHNsjKp4t16wZRF1b00aVacBKX7uYdy1iE4Fdpj18Pv/03VAc
PP0RKrbvSsGTPQYV3xReM6I1xsZdmYJlO1KeBcUZQH+KDbj/Fhq1zpr+5rz+W8x/h72hX8HtTeDH
1eL7eoLADsjQYlqMIcdoaW8GCO2kNz89Beu0P2UZI94uuptVanvH2tM8ZCN0SH8/j0z44d8ipKbT
IdF5hbquR0kVVqcKqA9mnVmLsSC2wHjYpgIP59pTvu5V+xYgPrjlTI5yc5ZQgs1wgslVq9snPoUp
NB4f6qmt9g1vzujfckB5zOQNNZ6GaeZT24RbH1moyv1CZRgrswy9uso0xkZiUu/wIr/pVQPjy22i
ACG9jqvsaJExvXxj3YQLZUzcrhIZgaddZL6AtFKM9ZXgYfY5XT5DO1C7u3yzcLTGfYcL55GRaEA0
AXYTV4K7J878GkTmPrTj5PlN9gfomcsbvymW4daoyIGp9cZ3nyfktXWOsDtTMbIVhsE4mW3XNaFj
hHD6YTGdHbcAWz3gzYyZO93sZ1YTI9Pl9Sl3g2zVelZPBoDjZ3Mkn59qSURe/9FyJdmJdCRA4b6C
y91AfHXbAKE+7FoJ5xTIDdmmZI01V61NryljrzqU24MWmwmDYuFC3hgHAk/Ee66CNcVFE5/IHw2X
bg2nmUXMH0vfXtipeFaz9IGBl7MPa3tblZ+YqB+LxabjbiwEH0V+P7ygomnLkoKoTar0VlJCS79R
4BcxnDdLu2wrxB7vT4+xNL1QGZyMp5mpECe0AFcCHeEfGETdIf7fFY5esTN2OPuEebtT/2s9G3HC
x8FKOrn1106myiIwht7D5ziNOHH9t1gSVWNkbEvG/GW4LZ6KLw4tWZvNKRiUq+y7GwjgRLqs+l1H
HXE8KmiaRH0lT9/J0rAI/ZcZfkKYSUCKWmOWJkoi+WovZGTke/V/V6psG2Wx21tmjOhUGT2fH3dw
iye3XYj2O6+LtzKpUE9NcfhJ1WfNawo/uZKACKx7EXJMUdRQwvl+WMAUozcPNAdhzk0bOU7r9Bsb
bSA2R/FOAAgbgvCX53z4Vr1iJeDviOvF+bL7OHH8FjJ0ZgXSkIdUkQnWJZRbnckAa8/XtlXSo9Fd
i6IEyXVf6/T6MSkfINGJpAJ2HxmsNX1R/cpJww6/8DKF2xDMgGa1XTYxDL2PGJn7zUuh0+huhOxx
KLKhOD9pEQx+2q7eeErsWRA4cbwF3F3EzoU8XYsJAOcvrqfXTIqIA6H3JwemnhYZRCQjdbPAoL7W
c++SCgxSsTZTtXpiEg9MNABw8yJ7tCLkmXFlH30YG/xbu2uZkDXgy5IoB2vsamCX0CKCpejVVITd
u7Cbqzsy2cHjfUf7bcSV7y+2wpDEc2zUBSXU6UkjNaLIgdzr905pFxr31yJHxHCuu01U46cjzKYc
Iumtg4fm6393OIRNqpwcZWbBRpg7+irFa6lxlAizuCdoP7QGYaYzOKIxw8ZAExJ7J5WXK+cAKNd1
OXKDVofAeHRMuBNJXllk4bdB1wZZIxZnMjK1iSr6AG4KhrkP6GDbqMzG6craxvdI4j+gH0h0iZ9J
60EVaI9rO3wE87KGJQCV+OYp4hoT6hiwEILDvsutr5z8CyCGnucWlghayr2b9+yyTmliPR/gtpuw
G23HKHo30DkzUU9LrjK0zkBR9BFCp6fAAicmimk6OXaVSDJBdjm5S9FB7YswOzp9wxnLhX6nuZXG
vyO+RU0GACVg48bF+sEEOuXAZVrttLXUrVTEsV2SVAWblaQAzHEY4VGknq8CptXJdTGRtx2Tnc31
YhCv4uGINoxyj+V+6JyPZbaMaXl0jt8NlXdN/s6lgYGQvlWM0Za0GM4mWjX7JU0VutmTdcBhpgWL
EzfoIpCdtjLsibqOaxloDG5Mf0knc7TFzfTowXvXF9ny+7k+SvHqd/+Ty4E50QPFhl2spLkPA35M
FYP2WESanbA8cPlOoC+/fqlANhL+Hj82bDzFJ/67fcG66IDJt+nXBOdmu2HxZ3QXOycMsg4533/x
UZ7904YTQAaIDzE4S+YopXjUus4aDPYQauSvzjifZBTETCgJCeDqrBvaQlqb6kxHQpbN0DtrsinR
o34qjEDHQ+WtU8xFJK5tWosBNYuIMk1uGKnNOoAU4bR1EeP938Fog0Tt8x0EPNv6W6DQCXRWhJsB
VrPfBLTgI0ebmC2d/d4+L0IaAsm97LE5vvir107mATuUEcnpnm4TFkwKL+KegIKLg8CULCOey99g
NMwjuxwwltvtJW6XQ0AiYM7n8XjhPU+dtNVwZniLYMXU9p0LQZdsFANq7QfTHMFNB/o77a7Elezt
cOZUPdSko62iZ4vKtBmn8rz05ybza17LwvQeB2MacVknsQkkbBuk1eVFszXgu7sjurM4fhBdSjKE
ChlnYPL9lgFD4zmrx+zPGmKbmYBvu7b/yiD4C8hr0O9eSvRGRTnUfQaPqmHFt0JQhpGxdlZ00J6M
VQkA7FWQxAqFibIxzO5guUdtLuk1w0jGUcSIwbFLIJpLRnr4cSsIgbiI26znD1NT+MJ54Nj2BSYs
uoDVslwvs/Ua5R2PAaBJoqc0y7quoLJBegmTeSrCOoP1sW3Jhkyc+zPDxsyBFKLB7bsCh+GvKEfr
cavKuxVhz7nXRl0tXGXTx9WK+jJ77JKlQwE9b2rvOICVFKLdc+k9Gh6pI+mAF2CQn40zrNjNhokz
0xWe6zXpPsSywU4phjKDUH9+cFS9ZnX9OpvuZ3DalcbV3FlLUJLL3Kw5W0OPwzx2KWM8f6q/7bq8
2UspV/KzDQzeP1AkolciHphjqsaj2RA3sgIPcpUH7bKPfo9tcqxCkMsjXdhqcxupo2KlT6E3cmbS
98N0womQ5oZ+ke+sLUA/0t2aeYzeNue4h0xCSnJ8B6O+4LfQSvkSTaO1zfdassys3QTBZSNbrblx
oxIWckgCLRwZvEYVw2Io3X2UFrrZX1ezOMa+/B/M7tq+gRlC6gzzT0erJ2W2V51EneGs7RE2acpd
dWPoYpYG1Ke3qRsIfLKOBmjvqXyStPXkZQqeaYul2NdsUJXZfKhrofLkmi4Pma7FV3vC26TScoze
Hwl/RDc2CLjIQNGB7gC0DbLOLgclpWTzaLG8OqB9gnwU1zcEggX0mVV0QlTG7fGeOB6gMPzLBI9+
YKI+CdiZhGHe5Jei7xITB0ccjjnQnepTerTIy1kn7B8BZhP7xMsaQ4hU4+xakDb5Wk1tqu5PXCue
jLv7qU9YJP0QyBRq9ZCVGn8XyOXr5xX70OGzmYPMgGh5XpnVwjOey2A/DCUTzmlR279C
`pragma protect end_protected
