// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qj6FKk/3V36h8ZKuz7w/hRvdOrBbT2r+LmwbOJrvxOwm8qxApX9vI19Ks/6t4vAKCMxhPGNyKMJi
EqNjwmoHWj7bYj+T7Sx93E7hCgI9jOeVppFUGedeny+wJdkv43f2tm8ROQHqK8aTVZizsK9TAf3w
oW9umdFZ6D1LYm+Uv1xID5dEVjfH64TACL28AVg3ZCmSzG0K7hpjCRbGgHhjaqkq78yBfbZYMexN
hDtmaLAmxVS2/adNQovVSntEqa425CPQiyGklHtD/pHxzQvi27PUVZmBhaac7b8PGMIwQVsgwMRl
DFpoXC5njKygSzsyk2XFjoqsB+bwp3kWW4U24A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11136)
PzCUdczo2HhtbyHtiwYAXI+uihM00Zy6cTLbbWmDm0UBeyEjcxljgc4E1nKJZQof/UOwlWXoWW4h
zpKjToDlHuGgK17TbMF9nuK648f/wCdzdmsjW4409wi6uHEpcwe/lxqlT+gybiHf37UszGX9wFnR
4FfalT9N2UNoFgatRtdid2+LYurxa//ozoCPqfyfKDqFpNuPISedmDRdaO168d8KCTnmjvJcgZVk
k8BxXM0ddAS0OFd65CBiDdiwvKczDIcf58blZ3qPgbCR8jgA8HLPspmqJlf8eNBopCCm6vwfv7TN
A+IzheqCQwUZWtybkG4qx4stOb2iUEESfMJFjMWKREeRAv66Ew4oWMh/tmu07juC0xQhj+WVF7ZN
w3ipyDk99BXgO9p/0B4FLfLKe4VFVY+57Ctdi4pZ8aHUfCd05ePmq7Jxj/4kpqKMzprpSG2WwpRz
NjT0W58kuq+huT7DSOTJlx/A+1ni4J1Ugj8PX3Q+8MAfTF1QEcyDFGoM/JAtnvgRQWyShTZHkbYo
CAQ9HDvzDnyW7/ccYCPxIkdtJIjWvwmtOea2HeGjMKGrsumyiF2EvEk5o/OPmwcXoClyzcsYUD3u
pFB2bIXmZTI6ekXG5h6puMF4nRH7MXKuimWDr+GhAZJv1HHtv92Ikm+xUaaSNbuTu+nDwZIh2AWv
b0AGNxhhgpUvvWwNfN9EiRyp9V0PBOF8dLozLSHOiJTqwh0VvuK14mo/Yjc90220zHvxMbH1Q18l
BG33MVSjfqo6K++28QAVZfY3BgP1N54qZ0Mi8bFw+U+p8vLHwF4e1lAcq3g7F/lI7Zzt+O9+dBKg
dJMqLB0G/CUtTcTHZlKvGd2pMRRPdMDbRN7F0OrvK+UCvTsXiyXuUUBcoPCeCd5r9a9NdMwcXnmx
9+Ww8e/ez4NOdaY9zNv9Wnq/XLvEa/pfJAw3HPy29c+JD+bgsOFeMpfTEA6AWeYOdnEEtCj/qpeH
37SrisCCeM30UnqlP/z5TZGEMHD/2ifEJamQDaClJLYTVaQrDBCNrcoV1AQYGCTfr7wMfy7sbRQa
VYRLewWqeVPUR0LsruLjol8NBcn+Qz8QMR3jlrp+LmZr/CQ4El8QoXGEAXd0sqNUU9yXvNSjQjDN
Yo8KhIWMEaHjgBWZwet4Xy/4ICwo8/aU9X6PGJtBlKO0e7M2QdsJVf7jsmcvE+JKEX5/RXm/fqPu
b6H/wjz9YR9mHaAxC8tpJziYBt+SGvKdxcYmD12QIn8padeJopuXAVydYdgmcdvS2CjrC/p7gE2t
dWQ6Pouf3D05HT0x9FtSwJ2ER8tnqIXS7Yg9T6BU2KIUi48Cvuh5gvpasS+FPncBQBbDMnVQ6zlc
ar2m7IwLCWIb4hUhb1D0fkQmtC7HdiWf1ayJNAEBT36mXq4MB12rGk5eHXdw3w/DUzBFA4vSaJuZ
ypUlMr56N4pcYEZFcQMHrRx4d1EjzEzaZhia2TuwPOFUMhJL0yGR9ql29mZ1qC8aDucRbkOjEuE9
k0NVGDnBecJsYVwya5NnWmh8S15Ak+iL+a4pvGE+suM60k6tlcZTAcgebhnVnnG+EQe9ltekDL5/
8I7oBtdt9OM7fRbdm54Dw1wAJ/Cvu4p/5sujwBQHyCxvwD705qX6xZl4lWliBGaIlEKwfUACj+Fy
oVO8JWTgOnWUywoDwozxiSW/H5qA2i5vryru0GDgHeDYLKoCu3H2BTRmEgH6bo3h3gyUhDITmYDq
kXzf8PIz3ZTO71PS+cobGbwSAHlP913cvntgR+2OMVDGPTs58OAjkjEim1wHKfCCE3vvThiv0lw9
/wlg+EvmZKnTp8TLXEKvcYdrdrzaM62Vo584HXEexdEmxNmGkdS4n23Ddc2J8PtNPgf2ky/M130k
e4ZYmAoK0W2RXh9jbbG94knolAZY1FSvibs+YlfLycnxcy06GDLBJ39QK1PbBLlVOQFKQBQEKoEv
C/9wcoa4ctiBmk4dV3N3Nht+uqT5XIUAW2Gy5D+nRrCVK0Y4CO6ec/zhGNZOJ45b98ALREqPZLCf
C47AH3Wlj17hfrWs1ggL8k42UEVCg+ISMUyN4/Z0anv+5BMQakw/LrnkXRqYGr9NR9syJMNLP58G
mrScSDQtgiw8oDK3K5ObsvD2dYJQ+NYpjw4ZQZEaDllMfOiK4aCONSHDEYfy0hr1xuKCX4feTh7J
G8d2g53hhMz107vCRwL/jTONEeV0IaA4jA1xqBiob0btCDGZAtoxOgBg1l+M6jn21u6p5IOZCibl
klZiU6mwcj49q1XFAZb0KxrOB7/cBhgN09rdbI/q8nEF6kG5qvsMPjYPzKKU1OMtGkcfWaMUpczo
rk5PfoZXUUADrGGXFGByFITWkv6g3SJEIRLCGi751cLFbN/UH60MtZBt2x3SjjKzpgHsN0pIUTdB
rXhkAEUeMtoqCyCHRxBIjBEUdaHCFNea5UgHnKL+wEk+x62RChgK/mg6WITzoKhXn1ueidBmm/3g
mZuBDW1rb52vjW93fs207R6/VcFbZGIYxFsEmtkeYtYveyiLq5FArozZSfOtRG2OBy5NGKBITO6e
UWfS+oHFvXSL+aJYymg8TuP7YWyg2hFkS1bM4On38BIBOi7Kpbj6tlmJa1Fi/80cwkUMSPw+TRp4
MmWeXaiobMoUWr6+4oKQfHiUmAGWOJQ4USotQmoE0TC+UmeEI517XVpuJqqEapvsB8bfeNCtISlD
pBWQRpkbKeRxQqYd/yiaX/T5o14Khsbi3wToAv4SL4pbJ8joYB+0TCtkBCgtE/VXiVJKeT8YDjKy
YMyQfEFq6sJOGfwHl2p5DDGt4rXPKW45Df+TmcXoNAxltq+gY10s09Bwf9UPWJQ7xHmbDdAjBOms
AesGw3RHO/ag16M8GcZ+dt0Xkej3YcLqVZp8G+dAIkCOYYKula4a2OApYn7zZcMQ+XkMOK5DZw1G
eTwZRiqwjeNIKu0ae6b2+QLc4fHvNAk/jDGs7c5ERMgYSfPKtNydO22uDIB+CDk9FNytHncYnMIk
VDfRNjEYNb2QAvMdUdroj9Z3+vqktBU0D0SnUmSYfph1VmAx8XfqnRFw7xJ9iivgYdaOP6dTESUi
MCe63FICL8/0Y6bZxI6sLt1FCh1bSd4zLLnYAFBxe0SSiUHibt5w+b2Fv72122qjIh+bA60D7GVo
j2JiL3tzgfLE24kQ5bW9UtgVDC4YDT08rLcDciqlaX9mDJ1YC2tzgmnDUgs97vX4iP7Qe78eA8Ls
CfOPkdxkwOjZMgf4PT+WNudrw7E+twZlc+yL/BhAVj1EPjpgfmC+9GOXZXICpZLKaqeF4UFvYLDk
HDJT3kNP5jR+3kzzfKzCyZ7pRb/xuUNT4KS88/qYBDluPbZnlDseafZAzDBus6YQzxZco8c4Nl5z
AGNT0GrvzdoFGBdtb5uTa3MpAIQi3GomYSH/8X9EnHmF3Uq67GPBvog+oiZQezJXM/T8Ms3aWPq3
AyYybKu4emmRybssF8zJNsJuDTaZuvQnt+w9fjfZD76n2POHtGxQ6vbuvqYHH6XY44Qlz7Nk8kiv
9xDTImIXD+WzYZN9FDI7c9b4PmfJZmTsa4peskhZYA5U1umAsqYcffDOxehmWOKT8SSfIkVHRCmA
7Tv+pdrUhF9WxYOmJ3Qj9n3BWFpHz9/4LDm9aDG2pPSyVuPUmTMt5xisGfuoXrNb7mzsDaRfSAGz
bEr4fK4SkSey+IazbFUdmflKwlJIF2ydhe1zoW976ENJYH5dJuDT0b1Q5DpzCQtyZ/VgTusd8UnQ
khEIgRRWya1wRSDRjcpmk2zI7ueFag9eWQgItPhT0nG4OyLBOtIx7Q7jOPijOO6++KHnM1AZ5Fwm
NKwGQzAqtA+Y0CXJ90cKLKFojPMxi8n4yam25aIjZC8iatLU0hN7k3xxR5Rft4RYPbhSw4fkmnzO
6NjFBOMS6By0DIKZXzAZrh5sX5aZ27s7LYjmQDpe8mkOmHKjOoNwrZDb13rqYMxiT9SaT+wiR+w3
5eVhVPcc9GilDJ43Ct5bC/T1FfxF9TjE+L9bWInxW7NZIzaUHMFz++HguRdvHNim7N77urBtGkvH
+q1p5RzuUQ6bgO7O5a+5jQxco7Miye466NAGClinpDECl95qxF2Pv+xPig6+cq0s+p4pj5g6vore
097Zp+aXsW8wJl2U5osng+a8/3XPCJRiD7D8GmC9cRuqrcgCAiMVoRwZrt3PXAeejtR/7Q4kLInD
q1S/LbXlL0Hryib/La95B/TtowvBfK6fuXFoU7PnZL3hZr2ymbFF9v5C9wQA9HY3FJOswucz36io
MlixQrPLsYXEeYQEl3r3/P/LJ6N+s0PQRRLZ7DloWjhwLOEDXbNspks2iuCdSX6GvNpxq5PXfo9X
DZbBsGG8pEBo4y0vHmj9ixh8Qy+8S696AvfiCLCDyISMbopjyIeBzfw42MlXOlK0t6BvuAGnDA1N
xgAoIzJTfTI8yC0Uz+c4lbI3o4qcu1JGqEMeLXjYj4OzNIsEGMr2AZnnoY6oVO4ApjBPDh4Mvrrb
BlM6A30UtfeaWpwSL1/SSzEOR4XY50GFaFK33vtpO4ysSlm25NQe7nNOQ9wo8LkmkNEsXtvE1/q6
HaRt5qzbgJap69TNz7DA7K362xIrffegMiWQMdxNJLye31C+DLvU5V1RStOHGUw0BB587y+HYCka
KP8GHl9m3HcIUvNJUXaB1BaIZlvosVtuEAfZEiQDzYLleHlq9aezq+JqUuFr3b21uycwBTQrGEQ6
DO1EHhEioDVI0Am4iNjeAE5ZBLvezdJls5kJOAaSsFGNsAhi1ICpMb4MclHhhRaDlBdG2Ml4a7U1
7QnPW6uH7wcgCtbFzs+m6evd4kqBRzwSb4Mk4Q7qxJn4kCCBAbHwA0OCjCQGNbEjtpLa5+hIGZkx
lIv3i5nCf1g2EkpBlU8bV4/rcWmmwgtk8wnxVkGZqZVcYvLqO/soVSabQrmQv8eDOMlLC5c/b8aJ
k4KmRTpI6uXt3+dZBHlpk8XOrf5pPt0hh6TQ336X+X+gycES3FmhdUgtKkemeoGoLvxSPnqFvRqf
3HRSxzUS+qksYUR3STmVUCIo8QifxatQECkuAP1Z8YNyCY1PspW5JTEAgHXPrOWMJjFQmtIJTiGD
IVQEFysj+4Bql+qqQkCwJPfB1NOqVIiKD7gv5w5OAcU/AuEshdtyk01nfpFGGauNSIie6vwnXqTL
8OV/meHnjXEy4BkUmd9qHeVRrGq+6QXj6bDw1+lZDHa2jFlgIiCuorK9IksN99PnpX6iJWRkRS0+
RKYRNs9cwyc+FvDUGSjb2s2VPOfMfOUmItjNyYK/hcaSJfM8hQp9skCJFwIIu73uBdY3p6jVr0Vw
LFiHk9oXFn3u5DSPn0vV7DjyMPSRVERtPq0y74O/fILZrRmAbCNDvHpR7OczmM+0FogIoAk5AreU
DxuFrPNvEhiwq7Pe2NUh7dPcw1BoFtcZmtI+CzEqBnqagvwBvNNLR7Lw+xN3eSB2UbopsjuBBEtZ
Am3f+fUDsTl/pW3s+yOU4hO4LxghbjqKGbfShoDBHXtC9Cr6T/9eqGanehwXWLUYtrcqHRUhdJL6
CQUpwY7rTdf18MjewwvX1hdcbq2eHqeuhT9ysJK4OWeW+uPpa7A1+Y3pcqHY7/eNIPi7pxXQvfD4
NVn9pl3skayGK9qacid8WURvPlIq1AKHSpE2y5a+O6s4ssjc0k1IwWvWwowBD0bowwl+9QxSAcX8
FpkglseIMZNmXjivtCgGb7eSmpC+nW3plppVdix96PxOaz1W2W+tNqwggeo8xY82GwfnsekdnJAd
73nwzQj2ai+ZzNcm1sIh2izid8wTDLs+eriU+o9AJZEtbP+2lV9ddqb5s5hBGm6rdU+7NBz8NPDJ
zep37wBeM8yKkBqiRoIccyLm2ILPJVO2skaoyLQvZu1EerjT4LgHhzmgdpZt8Qs6Ayi7nebfQBQX
OkGSwM40q5jBcK/ZaWvwpmKA/TpJ4mJKnySYnPllkFkh394XQHNu+ntrUA9LkwTBi05phmFIjfdH
aQ4EL2MyaeYIsIHblwuC9dnmMRJauZ7V99fX2i/Co0TsHMOFKzL8XXvfDsE22RwIbZ5EL3Hcp6w/
S1z9bWL1aj6Z87dqbNS5YYUo8ffMfyZho1vzaJEg5dzc15nnhKTlj2M34k3zN1pn3JnruNFH+H+v
TreAWG0ZiRfG18WNFmHCn4HvzuRgjRHpRXOr7FrxjXIhM35bEM34tk6la45GgX78yaWVwspfYWx6
vB9boWbvnXkgeygDlit5IBFk1SJ47SpgTydeegeSmKLYE4ihOtpimo8XkRbj9lELQYZCblgaoUV3
y2A90+eC7QnwqtY93qMWj0D9FbIg29QOk9Libudrfksf5ifRw6KKNg+Lrf/k/hw63DD99udJldN3
6qy9IsCGUAy85E8h/R3HpO9eFLD8ubrdFs1Z9vrfQxG/3/QwxF71cRgqBcOf/KoLsO5V8Ys9SfXk
KnOynoA5Fb2D+im0wDaDJyVmFz58piFgi6NUNJxGAkU31JvVf4icCV1hdHDK831sMe79s6cHvtSD
7vg4r1z1yk2ef1CgCtyFFfpYZwy6Zh8cBvRzSu8Er3G7U9e89S7RG8uj+3gSn7WEuBrpmaiVnZ6f
FNsQ8XsTaoAAQ3XeHJo6OxpxYuglOfoElI0ZZLte9rkpX2IdU3cosDliOS/kgC5PyWIQ0ZhgC3wv
CIURMhQjzVh7ZQdo8f4eelQbQaBZaqrQ+atmTyobSjxxA/i5JHjsORwlj+bXpFW4l09LWVlFx58H
EfNbpS6TyfRL/BXAs65BLa6cP36osnOd/MzbFA2qrxbs3vDtsLBmmoEwoGPubsjbr4BCTPAVI/Tu
hWgL8smLDIulFL+ezQ/1C5s+dpO7I+CNC9OWS9r6J2136QimZ2/3UrjoA0EbR1l0SpPZDEBDv0V7
APMIPIQy6qdMQLBxqjyjlBYM/t8AOwaRJooGOYdW3nySfBgkTq24vN//b5F3nk+duvqx/sRxR8ca
3WjmNwGy0xA4AQi3ZHx7Z2U1Ier6YfAxT4bsVK+gXy11rIxCkkQmTuwXhtoMt2rfwupcnTG2M7Lh
qg0FIe7N8iM8nOxjnVoHotioDEGDitKPW2Wb1NafASP2W4SHfEo/0KHsiKMA+qcX7XOUt+WLPR4a
bQWVoN3W092xnscOCX4Fx149FToHJ1QaRVhfCe3ydlM0BFUSo8P9OJsvCeyLoQsBNX2qH61pHd9X
IJ/kHq77N2XfQiPS8KZ2gHGquShvpNZgjfU5WVpjVtBRuD7GIHfoFOwjIQFdjO0CXHucPHvo3Osr
R9d9eROcIbxAGID71YuWH+3EVYpVlgeuiAaeLYC+PcdkeGsT43AnXC4oKSB3Wih/YqxbffqsjLQq
lVo42ZKbGAqD81uXtVKcsDmnHTP3k4q6GOJZQ89QIhgypdA/TEiVTPaU8tnXkTowmw2+A47CIh5N
e9EGUGmJPyAdl5CMxUJFJxDvoQB0MPuhxD8r27K8fAyLcMI2OvpYUa3A2OVCgl0QOFZLibezlSQc
iLtpcF6cvEeSmO9q9D4XFR/15HfPSRuPoEpq04ujJfWCIa3medVqDVJ5QHI0Do4LUcvae1Gv0di+
UAZw/7WKZ4LOB7cqqWWOgivpCxx17AdOiSnEN7HpJRJYwF0QHFW4rp+r0BM8h50ahrXGhaUb8Yx0
GHqg54OFiYmE/k91RelIoakgPzA6AssLSCpABpuxdpphNNDkjh+1zHI/prRDtoS8V2rxsvNfGd0j
ujkUiHW7BSyRP4aBKYKQ3J7bigSjFLnOCk6tkrBFDcI31a+tq1USV8WhJ1GPlJrWWehP4Oj3wIlJ
k7DLi0RKHaawDrw9hJ7YPzLHDQPSHK6u65KD8MK3FVYMp34CM7hOOVKrvBbN2d82hjNunUbXiQ7b
r4OX3i7kUOQW/AQlq+mW62bfMDOG/NcRD1NMoSwnV5PpfGjeaF/kGsIAJfQua8I8Fs1ygfD/EOQx
0sTpeSZYF+CqpPWlOzrUZJmZC2zkH55TKvSqe55eUbWontA99XWJGC48k6/xNynZfgHIZumc8FrE
0ZeT/LWYUuzbebLTNZs9jzGvLn+/iVOeqNr94BJsl7OnY373gcGvp1NlZII4DQlP4x16fUXmAz6u
LbakzyDfueyeHd6sot6iRyR9ceE8vL1oxTDElXWk2hUVIyELTtp4WebiiMsHyb1E6FZILZuaxLyj
90kXx0HAd1A+BHwsCzGdIgfNL9DJ+/IeTBFAEkE8l7dYM341KXD1dQ4ljwRKwfzvdixMT2BcDiL4
YMWVFmLUvZ3tjcgAE5PyXVnbg0PObi3MeNNZ0T93cxjJbts5E7fCiWdHc9VfxI5yGUKnnWutlpxY
ZyIoZF86a0sLbj4JcZs3LkIf5zJXLHt6+BiP9/x8rndcSPLuP75cNQNN+dQjp2+yyWk4LeoAqEfA
O+bNbwxgv2qZQuYAwBKXPdC9CexAPF90Fx4v4UrrnNrpzRz5Ctcvz/sy3ZL3jPKlQRQh5Ks9JD+F
SOJJs92dSD5ttEsaKXD7JUoEsPG8Q+xHE7jC8R5elQR+v6EZCWXr+b0lEGc4PSKzG8VBzbjtAkk4
7V3D44kyzfJ6yzMVpe6pgVvFq+pzVuTfDNHzCf0SZbpyDiRVlYdWjHq5ZY+C+JvnPitwZwCEoJMi
9E/PYwf/Wza8NVGyVvfduUVkGtHo+5oqQceHpuRPo/MsteDWXtxvqs8+a8JhUU9DNtiXXwF94S9U
NHLCVi/z/ZFB5IQY3/0ZN+5/yLMuRRiviRRasLqNNyt8YRoWyqlLvyqicWoFAgJXE91OUlhz3mcl
ujB51Z9x0GLL7nR9Vifg83WcyNVfuD5tnNfGYoCELJis7eXg/UXjQv/dFlG2IJw4uBxdvOnmpiM8
qOWSoBqZHN0axyifLLohNiEHF8vBur4PTMeaUu5S+iuW/O7rJJvNBRqEGYbjJZvNhWfb0LyYPjZh
JpsGRp0muNWT5ew+hEYeNOpCZV3jksI+js6fTTeMe146zHeOxvWA70/fWPrc2vdukXMkcc5m1nNQ
5scdhISswEZ7SrtNMksRNGzjWiYqM77HtQRlOdsv7JBCKmTK/hsJFmtcYY2FJrMJbSSuMwE4ZTzz
MFclziFr/tMAmUAEAbXspvJqTMhOAqM7+vkMwEQpmcMBJI+brITrVMicokGMpxY3WNBuThwVRwC3
r+Dr3nkDGLAnMvwpGqLO+RLVUAUJLGDJHDqQMRlO4HRwOvpshEWh/wGDH5gXsoA7nZzKv0/b56v8
FQU6ITNyJ4NtWGpx3aBfJpx81IzSkFweeky9VfMnTAXE7LnW1UT79GsVSw5V5gH0kHSOlX/VVf9R
kYwnvIo4HqUWUh9GceamRuPK3GMvrnXT6Ukj+1+hHOisYeQ2Fw/df1/uUJ484vwH/qVXPH+Wd4J0
HXXQCMCiIIPXcKu/rS/fYNzn2Yh46XDKBOaLk+69+q6B28La02PTLR9xgaTx8tvN2Vkf0latBaZE
KNGqZSs59UDFB61Pub23yt2RgiTYPRpan0BQ9IvqS7DMzYhE5OGCVofWHuNKwpJ9RMysoYfDaeat
7afEP/4HJvfWol+j6YOsVM9osOm1BgAozBRUR5stKHLS1HcDzbIs8ktH9E9RvY2Um1w/19SjWvJR
7/g8/OUt+EW16DOZMRZmZ7ui8H5E9U1dokfeFhevq2CV4mDbeqXGhWQPD7qeZgwg3OLUDyg47W0t
YsShZcwAsnrg7042e/+NC0yGwi8nL3fGCFQx44mHK3NkmEIj3jk05H16tR1ePk8rlOrJZqNQlV6R
88+v7jJ/ZDGiqSRV/TGs9wLIdHGnKeDRgdNoGysUagurubqTxZcZagrROybX1yidXmSrqTEBse7p
oUkrbi3JL7hrukGl63NUwqTL/MvICC038uxwWPoGLT6vbeoL56J8RI2NtSv1aMDJKW2pemI+E8rn
NyQ9qBDsSL1Myw5nRuZmNFRNjCb/267eedgPvqejQwSXDb8K56dD1/X6LP5e099xt7ndg84LtyPr
Ye70javlOAhBFlEpKdkOZJPLUvQIVD+CYa8zJXZ5eb4eZuR2dGYCKDzzWKpGTDDGRf4Ggr/wD6CH
pxPYy74HaDoAh85DsgTYlnIi2rTUwggnhJ24ZFeurqWC9y7F6Z06QaLUJnW1E0LODcDQNbaVc4yB
9fFueDSKyutki32ewrsYNooPczBxrc9AF2eiYoovyL1VV/SU8pdtPXPVQKPLVL5XTWOKw7vTX+XY
l3b8SmtVFExxFrGmJCEyFLe63KDNSIq9ksQqCNJ4V+RoER432H+7WwDOtaiwPXXARgKVGNsDeggQ
/QkLWV4Div8fIBL2mYTpyoYOnMALifumCizBdOOv3abj5mK7gmf0Ivoowo4++Bh0B3T8cwUOwhQt
Hf2sB0PA1937dil6Os9X7wdF7nFWNJ57CV1uNFY7EeMnalpdQryQDPQlQnQRRYy/eeJ2YwJJaaT9
x4kBu6cwKEAhn75Kz5y5AOOvmeAUoGcWxKELF4GU12XXpPeppooT8j0eYR4Yb/VBY8qTlV8aNSL4
hTBIo9jBd1rP0foPi3SV0niWAViCYJLQWTcZDHqX8qW4THMFjrClUoMJzoxM5Jjo7szQtp6N6Mzp
7oAEef27nHZMLBOh9t3RZyiLCoOzUZEsbob+3SAv3URR9oAA0KummpsobLaQG1oqs2iGvgSCRCKh
TH2fmbiGFugDnG65ITTtJtNJ84X6hi+szPqYrNUT1f9g61EMpvcqG1Fx4MbP8tsNz9dPm9mrUMCn
kwmhfc+g0a7L3ldoePgGOaZAdwopB2M8vdMjug1Zc3vN4Z0Mg4jPxb+67QHzlvnSiJrrRBUf79Ok
JOVTr2tTQo4LFq46AwP5haPqo8i40xsQQAtBanHQ9Km1RrM6ej31ZwQR/oR88QHgpCXUqg8e4Rv1
8C76sv6nPOINrNY6Txh/yCNrd7+kGTk6gdIrKvgE+ZCc/Y1F8THOmvQRCqCMXxMV+6u40+NXmheG
EllDFrZCeHhQmxB98LDP51D6UWhgdOCpgcJOjq9IUaOmNK+sarhMvmWjoJLRI7He5Iw6YZFw7qt9
mElLXcZYTzdSHSxutmP0SwvZrLjNL1HQAnTVc1vHpaAqEFMxQafvRCpE38k4g9pvdfuVyE4Kq/xC
L5qUrVenLovJ5/fl+tIaEKFdK+L5yFM9rV6UNyyAbMn9G9X0WmnLykQXn3lbwYkqOg5D/xaKDpDN
qwVq+NF35UkZhaQXGpHxMMeWmtEnDw67PAjaAEJnPzPZwSw+UlZz6GPc4iLjArfbdlmN6Tb4R6dE
cSaR7egpcJrXx4i8AP0cfVAAX/VO3trS+3cb0ciNeOz2Yq2b/ZhQhZpc1wXR+BFKHVP9Y+/tWvkn
acBnopZXANnapz596KXLWiruSDfk0sxLtPEKBoVm1aT7XjVwfO/I3uRPUA27bcj6ztIKDrnvANNa
hHbe/pBFesIkWyGkGOxCUNHy9ZROgPDClyNdCAuBkioiDV+qxdcBsPuJHjjztMssSZVKbF29eowN
HSvhXC99HTUaagufYtDBVSdxc+yuPb0j/1VadTvnzpg9wAARNf+WbXZez8H6SN0akhXennCB6tiy
CIYqstnT1+Sjny9LHYGWZc7YYBLlByRUJgI/T8KcS4yH4HYvP0YhKfRmny6lTbb+zZjQuMQdfGdU
/6CXi5Yud7rJCtFXDNTLJFw2UiD9c4QafyQkziPje3mxKxFno8SmZ++pJVKorP7X13aKN8/bfDph
oCps8bbg/I7yfDo9uBhV5BmARwvw9Wtzv5TKoeSoI/NsD/UeG89POUBHtsQttCPErjDd2ysGRvaA
CNQkbYt0nYcGJP5dfUVXYSnowr+PWzPvgDBlRHTB6k+OMvRIKyCdPhDWhzkOXUmoWuTNuRqFSgxr
Mwg8pONlTOnx+jaIS67d2TI+ejhpjDTTy+0oEKW16TpRnFKkeoYT3cGwdIWWsMgYqB93UjQI0BFj
jtdHKEAtMwhQvS03BG1nNfgUsdoIxpRk2CXECuqYlZkv0i9ItQl4yeGb/tTaw+1QVMqE7U87pLcf
eYMgikP2jS1u3NfSqaUfH0UFCUf1b3lIjCLxHkhvXlIceUrHI3jY1msJvGVQY+NROTnNDVpDjmWM
04Edwg9nK13BDNHtTIW5cgZ2Ys26GYX17seWXcdTMjN2R3DPdv0or1SYykrN0LW2u+RYSPQnSaOE
ErG92YgR1q0/Ew+kL/KHhS7FTgMTRmrPr4v/pSjKCSQzIn5o66FQ7n3nub8lvWsk68QRTj1PHrii
iRVhByeR9y9N1I0OjKFX0KoisB6mZakLCVr3Rt4Is//DtwsIgrFo7ulIEMWc/vBJMdLejP4DkkmW
uXb07AJ22rxrLYYr+QJEP+glg4rfuIUkfdvssmtpUw7QkMY+7KM0oHdxe6npzuLa0hENYTX18ete
2yoF0VLbUKOCSLSCaAWy3IkUZ4KiAaxrrZF9iE8zDtflQNngTRd5SLfOE/bT6mccQsWkEU3zOU+L
MgJehuTa0WDmXjKRP18KbJXjnFCFQJdcgScJI02YkfD++A/NM7c83ZUSW2UmljBgiah6bUnZpWmz
fxluLJoeyyB9PkY+x5Bmpay6UKdJKi79o138lNxcYxG1xB4wVh0P/uDxZczMDjlk1ftRhAxytmk7
TcKqmxMPiNLKMaOeXAM6h/NjhPSo//Qpob1B1L/2IzMr3Xh3a5nm/u6dtmMna2A0pjoLZSb1RW8M
QYVTYjALvU+sNE3ElLFX5JZxFBSlN2kSUNZRIcm6cPI0m16uoxI+TTQAy72S8py6/qW3Pzq1Hm9Q
fBsfFtFXBwn315pkXiS/V3tnmC8InxonbSm/Zmw+57F6fRgk3xNJK/jmAMoGvexFpYP8E8+v1y5M
3T/hObC7o/5AOE0IN2ch+F0ls/0Hj/igfbpuPSv1izTCXfM/UPRgMJYpYk3j058tSyuVNKp+jFM1
YYGHrdilN1h6sStKgtCLVKUo7InIsv+sgxUaBoygGTE1kpcLowWrILcf7F2tKyhpS6AE0mPNCcPe
w1EfgVAp19xL7s0pEgi42Mm2FnbThOwXf/ns+WakWiF4XGuvI8cPHMDWN9PV+xl/tOPhy3CwssXf
sQXmT0zujbRpggDsM3GwhCW2j77gwJIZ9U04k8RKRF2/wQKslHLFP/BBDQCyifoKzmmVO4QpMFot
Tdl+o7etGsIUSxTG6BIOcE6Xw5DFYsJSyq6KF1083lLzrer2/QdKUOA8/Wfe0+/oiMBSRofxnENr
Nr31mH0S5T+JXZ/RCY2Ebr1WJH9GhvhCHV3freUb/KEmHTbSDhmL9QZ96ZFIfyfHWGTMZKaej1Rr
19FCl/Bhl9kl5HXoO1M2e2pfl+gBjEFwKSDf2oHIlMbW68+a2qGpqtppFeLLuwegfjicLSHNpXHM
wUde1poqS6LcHsm5zQTiDYdadwcoVLFoxy8KuIqb9xkOvk9w5Go927cQ6boPTrgrLsfk13yMfWG4
E3xoKQdJw8VXklDbx3CKVOGhU+lu8GtPK0fwNyXPaBHtNdPcfPxzgXRD8+n+o+jYg3Z5kPWzzJd3
gG51lszicv1E77TKQbz6ll+jMW3tn1P+hiFD06nbODZFFU5NQiQUld3/D9enJasOOWPZ0tM4Iu3r
p4EQAilCQFMrpAoR4sFChdTJOWpZ0sIbX6x2PmDr1haEn3/530l4GaQf6WafxiCCJg4I2s9ALX68
JYXtTonIYzik5G6LTY7K8IE4jFrDivWgrIsAnteq7NvBIbW3mE9BZoW/datqRh86NODD3zGGuSaf
MFRKYuDSHr5UAzmQaoB+oVcwuaGceCgnNAmRKYOeKCdHDPzuBtyKL9YxxbQZ4eBBD5zI7ue83g4h
uT/AicqJ3qMvqmtwjCOpZ98R2SnrQ9Ct7galGzobYgP9cudhsX66RYbbiccKvBWUMBZU8i6l7QHw
T84T22gxUyyUv+ALWy18sFbKauo3Hkx3Bi0W7V6OwNbCz8Ax5rc6OukBjBD+dK5v99FYX3Rj7Ywe
rLD2rpq/znCB3MjGTcLoyytmAT+mncwT3v6w5/ZO4RtqAxLJM+WYn+oeNJHqhC+JC7jRHplmexpX
GuM2m/SQ5eJI90oZpBD5hjA8JMKk4ONCMxbisloI1gWRzjB615FwMNaIv1rV5z0l2StRsKdtHCKE
8HLrEQM4QMRwRy3hUjfZ5pqedReESTaZwWnGzqjY59GYUKeRZrIMi2AEdeHXu+2UysM1R1lZsuVg
c2dd8XYK5q4mCViMAJm6fGfx5ZUpixPEZh54jmPvMYu22yix6G0HJTvogiVVcXu1nXaIyA84x+gc
uqmpqvViOru9yajEV3Rb2NVik2W1ieGhGiN6mGii2UFZt4yxTPtuP4Z6xI0nt1Of707tMDsvHgEk
0kOJ4pA2NQme6rbUefbM5nC6cJiThneyJ51q0SK4f2GfXjf/282CWa0Dv9MRgUQDmvZqdFwYnWgx
jNA2dqMmxJkDvRzUUwqyvy3HLavxACHRTKAX9k01WFtiTADq+FMKuC2z9358ixVuaPI3UpNDUffD
9NuqmVqpEE/6RgKrXKpRuw7alLjCye1tluyEKftcULkDEVwRMyaX9hqhPlczXYikdNJb3InnHn3e
q56Xjs57ESomXFzsqyzpqtdl3cqBbyaf1NQoYLJep+34mqKiYGjQ8kFUe1B11pEWVBjQ0o48UTRE
TieUymQDfPGONnMV3698afY3rBCB
`pragma protect end_protected
