// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
frPk+i0HTdipTIuNQgw+D77UEAMraxVZkU16wma5bpb0HYIA2XAe53jr9UhScfk4cCPz8UTNVPu+
9moNFSyvhKHDi9V3CyOQRsTxXeWsxYOKvp810lbB4NGSTONY450qyQhIt3UZJwNKAd+jInDXvl7Q
Y5I4YzIlcKDsKlLcM86uy7NbgSD8jSjb7j39S9kO6TkSKP0W2bi8qDiIdi8ksxz59WIIP5hw/nTm
rMDI35yXmtIGY4yZTAKfaZ/rmZt0NE7qcoF1HFcn4ISSUqvb0TLzgdKz7zdhRrVhSgtXxDBk34xw
MbvIHz5M7Gljs1sXeMSoO89kMl0QqFTTycu0lw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7600)
4pMBIofqxm67PLaPGipaCElwlZOeOgRygOV34hCDgZILQ8dyT6/fy0jSKPWAsur2qTQ5QfhWBi+G
opNPK43G4BnIhDrcL78wLh9qntdXJaP7zE5XuSNkVi6GqXvIkLCK+UwHtqXoNDrBEyRxAQo7REoB
8pQPTU8hq9/4sNgTiJyj1pwtrAOkCcRZfpz1j40ADPyWkKp2h6OE+AMbPWpbmP+KqJOVOzy2PcJ+
JyaZizrBqudoXpsZIBJ1bcBLBTXQJMT4XkfEQkiJyKg7c9JkJ/mA6tqpR1QYjF8Dpe0KuRO7mR4A
d7+R9ukAnuUQWZJ7DJTMxeF2GLkdaDt+OXuphRii9bSRgQZMq0n2yLyyFZp53rQxF8PsNyQ38E0O
Z4vewf3S4lhMWxP3riLWjQtekr4Y9D8tp1GabMEwwFN/VBlVccxEFU2MB/fqemQFmG0quSjpPEg6
ILQiwb1KWoyVyVGXIqp0gQehaWVQ6B8wWFHaqLXyDHUcJRrar12Y519DQB2TWPhoCSn8RDwySKrq
9koRnIAXO7uyjhhaS2EuifmeYnjDNiBIRI3DZn8/TQnXDucE0Hle7P2XgjqxsOtrM+oAt4NPdtY/
pzejWBP4Oxq0fyznLc8khy+jFSH0gfReRH03DDyf8L/NWE0q/tmu21kcBhOCyHsnJLsmUp/AzAID
eZiaZfcEDLMwD/nv3J1frSsoQ8zuxUJXj76M8rw4nlTYlXtcFc5GC0K0W0QKQ1liQoQPPDfLKkX9
PTlxKn6ksHaWIu0V3TIWe3CLQLPgGMi9eTGgY7V7g2BCEURIGnAXJqfuIAWAOicAVUYPSIL0ImuD
jjTI1q8LoaQqQ/9F+FuWhGwTM4EntkAi0Loz4mKL5YE3/fZdK3ZEmSSPNr0hSPNI0pkPwKPE3hsp
T4nZ49O3HGIt1AgWhH82posl9bGpJaeejuh+p94mnfduaVAS4qNZH9fO9MVr0HocwbSc9LNME8I7
TXzbE6mXbzxdsNO1a9X6y2Sj9dT7EX7Mt2yaJGl4m4LqS85QZ4Qdp7TywJMRzbkIGR6jyabK0ZW2
0qqEdN3OfNylcQy7KmCQw5BQ29qud95xXz2lV5Ci4OJ5HExUIl58WFYDcaPZ8B9t/iSceAH27eH7
yCJL/TxZUDvQM4WR3/+448xAs6V+YAO0tr1SrGB7NQ2wvpOJMVnULTIYenApI1DKwKskW4IK9RAK
2QYjnDpo2Npz2LMQCyrIKRDAvATGVsjrB7x1ymA88DLhEGCbj0MHj8GkDYLNmkSqcbmNpD49diJE
O3su4sX5s+ftwmPJE04Z8cyG3d2vwhwtMDbcDZ3GcGgBmupAr2WomVpVIsJTU3pLepDzZcTxB2Ii
3Pe1IU9sauZAmTk0fu2fNKoDaMAzWIAyDwwLonZANMoiVLY8RTSn1VShPJPoZbtsfylXh6wMjqo8
BsHBKQRFRAVfAatx/yNTVArajIX/EzWF/II4OkF4MSdSX6bTrOsF4o7tUBj+BQNffmXG+tp/wM03
hVnaeGmA9CnjgqtCYxJ9ZLqAX1SEUQMRpIPjCWFsgNG/8qtcEfLrMi6c5FXOcK9vzlaq9BbssI47
sGfP6eQlDKiDBlmtFWpKo3RbHWlOXpP99lwa59XJraGpyaNmpF0gVEZMb5j6ZeIxNjyPncY9KXky
Y9AgAVEbXxHIiFG7TUV8ZxMJAXtCZNZQPYc7hYa2eNduXAYYOQU84J4kYfIaD1SDGx+Fxto/Okke
MXbHEOvfjSCl5gtpBYx+o783OlQtV7/VdNqJTThFnFuGLqBc/h38sFrwp37JvmRfDprHKco1B9/S
zXbEvEznVSyICVgXRuo0O9qaQcwuqBS2R68FdkhFXtaCV04CBf6f9Dx8PdBQw1R2qOuig6No8Hzq
rmDuEyBb1md/m39D9V19ANXljKiuZICDX7QQn0dIDbmMaH/hnOkX5/0mbIkDInznRO8u5R4l/ufl
GCifoeKOO6WzUzrSWwkG4Kel4w+pV1CrVxx7LRdX5M3jid0NY8g8OQGQYX7zMHfKCzwXKIoaN73T
sQSIgiwnageijGAfzbF97f9hIDVG8SfijvhjFpev1ClZhCktlpya/ekP8N5dMlk34q4nRI0qU0Wn
Dh2Z+975aFWQBq6oiI8UwZgfXOFe1m8vcgy63yMLqwKETMNRx/KJn9AyLU6NRlvXEpqON5ajCBhU
RtlEPAi+BkK0qZPk4ELE1Kw3WFJYaOs/bFEFdX+O3GXC8G87tu9MhdCrKYjApaREoh/KjmiLR1gB
lhRBhsV3Mmo5SEeSKV/tyWD11hxu0vUS7ud3/FbDy1FTGOzt+ie6UyIfTtwC38TIietUNKei0SDR
6jwb7Ig+ei9h1QSHeRJkCpGgTpvyOghuTz2dVzTp1v8wzGRww5ZE9/XaISiVuGIhpNZAFhpTQe/6
C73fLAJh3MG1i4INozE7NYrXXYdos4uWPZ8p+wtDaMJZ4han1ZnlDWxu5BGMau/qgOTjEFVRzw1e
DxWBwjFC08c4DvGk3F0VAYI5jqR/rxWiQvz/B/hj8wNYEitPAt892/ucyIFnSsU27mE1FDz9xZrM
+Nk/8rtLKTIDqSt8+6xAte8DJJl1+YTomgxlTZn1/jvumabVxhUNCGJEKgI0q7ZJiiZhhMKGRfnR
20qcChHFMcKTWNZSQrbxwPTWB0XDJrc8551gZhb9f6Y8wMAZ7upcd/mINO622naXs7/rUZLB1pWn
toLFUdPlwR5mhdTy80HV09Ka3eIv2oAiduymVkNZKLF9fb/AtvijR18ZeQbGJSoLuC8EqNUCoCct
AcIM0/z7WS9IhR8m5H3s/0yKIzCdRQmaQpwhBGHcHQoT0oJM3bWElDF0d0s+dzCXXpdNyx+Zkyrj
+c7oUComnocCcujyPQZotqP3QFoyAlaEd50RtJG4kNpFdtGIxPCVkxMGI/9G0b5igBX9Ter0FofW
/x7UnJLgkP9SzR5TuDL1YtW0HAMXDLDPa4Udzw0Ho/H2bc2gzepXrkM3k5FywJ9to5oqOZBtOMN+
GcLSUiTi/1gJOEUcD/mlycJXFX0xWTGmsQt7Cj0ZKKJO+hIG2ZEWxmZkmS+8Et38EpZlFeCDiJTm
s8onBw8Uh2oNK0nkIN/288yDO4Kpgqn92coH63V3VfFDjjZ3MZgp1Q6gLJ1QQekZ8SCENkAvscNi
VO4fyqeLS3N2jByXdmrdqgMAcZMJYnfWJOjtVFHRA/K1+0Fp9hFf4K3o8SPKLxKiEy21rjukpurK
gPv3TKFhVwtwD1e4/cmQv0A2bJN1JLMD1xxPylJo0PZ+Pb0IKpUnb/MXrv/dc8krC5k8AMEhC5a/
56yM87fSfZPq53A50G/nNA2Uz47Mw6DXQ+RLRIh3/KUXRN2ZGP17iyz3U6vIixVHnwpyLjK16131
SWrONq+qw1LdzGEphx1p3O6BkmtrySVP+q7qw7N1chr/qAAsw3QJYtZr2UL645UNXLTDULU1+AdJ
Ndj1QcEb8CHfhBHHAnOwqop28tmz1Yu0Iz2seFirMY7y3ksMBhVikTC0QqEKEoIBnncVUrhZuQKL
F1xNt3WesiGs33DSrGGBaa14Awrv2g8m1Ucog5ManCajnJQqGVVK5kXT2Rg0ePuNg2YN+5/15zWh
M/yGhVF+FwgKmUqXeg6INeU5EZTiHE4lS9Rf6LhclMPsG9q6/hisa3vdgrZvLIl3t7elV03W8JoZ
CWpjQOevk/Gho03K3v2EnQG4L5vYSc6zBVBiFpHa3+W4gB7hQVcmMQF/RnYGaaJUg5w/HHlD4v0z
30eJYhusp62hKB/sYXGllxbow4xKSqEsD2gEcJfn4zdyidVKMw6ng9Lmz+NVz4RnXfVZxuvHhd50
KmdRTtKmmS0Jx8Ab6vVuDlinBZjBW5QV7oBiDsCVFhY3ygmnPzQKAfKQ8LYR6VGfr1JyqFYCUAe/
0D/BA90o+qJAgsviQ/jSVh7U2aTIDKUnE0yEyLJp0fFv6dfaXBZQUKCMdbIt0l//Em+NxUwH7EZ6
KbGLTPKqSeYLCjXCbQDTovilFlXNn6acQkU+Ugq1dPk91uQmuF6M4PXujRIzzj+HddpqdnY7/fyt
CtWb699VdryQPVJXz8rDmrPqfrozgeENCdpIqrDQpiX6Jw3vC4uzcerJxcjeknT55S8i2RhfVTgn
fNCsJCAtvpId1Cve4SuliwKEN81fzwZ4+yZ6e8VB6MizxVVh7ZSZbabWNcfc5MeFRB2uK+I68tER
URgLpGzxfkaYDb/v87BAMQYB/5159Icn1clgKtDkhyzsAw/e4EDaeIUqTE+KbKb/cLidEHl1qDsQ
bZAGYpvFaXTw1O8m+O4ElzxFWa0dicGooXgwbUtlX3GVkfcdJbqHK1xfEkq/nIk0EFe+cm3dym/g
R1YsateMHnATM6xrhRNXUyA22BMXGICtPMcmOHvjbTN9rPEfdXH9+/aTxcgPrQDtEtrSXkHCNJrV
ulV4gVH9LLGsWJzr9AC0XCKsCmYPlctZGflqdyV7NYQw8un6Pz9IIiwaiYUBRR+l9jYAcMoPe6Dd
eQieYLfBlTFVKp1/zF1R4wv4nrZTdyKmCS36FM1HT/NMP7R+KBSomJggPeBxo672mHESGiaFsL3o
9rEZsI98P2QY/7+WSF5/k+xBI1uiftQgMZWaihxow3wjWcv9/2r99sZ81nVVc+pIeme4XOg9C37r
24XGLkwgE/ZbYuLAhLBEjMGa+6bd9KZ++nBiLHvQHtLVlKL3BwVd8sPYNXtESuQHpC4u86HXKskh
yyug9CtoGB5k69JtNKX5VvxAUrbBAY7rC85MKQfs167RJxKh8JvzE4iReE+LmAEIsd4qbekQ6+FM
E1NX9mhaRcpMslBwmB6vyuruznPgWNcgJmRNFtAHxvtU3BNR4Y6sTSHszWoVOQ12FB95331+0Ije
JRDcQBKAXtfMW0A9t4ZrzGA2mZY31svGFF/ni1icl17A3qAQvoGbH9WfsjtRmd7Jdc7p3uV8sv/k
zKMZ8ZYUFIBMKmcMSTzcrUL1LoC19qLjHtkaNp5UTZnm8UeYcoAk1Hu+1AjU3IJcXYHIQqdBGD0c
HXUEoi7ot1T/RD4OYeu9LCHG7SsU35CCytt/dsd/q2IHB+/QGS1jEZFK8Lj62A2/BV1RydmbfUjS
v8nQizjJipM67dg6Q7Pime24e/kxm+OMpY323NP2I/JBC9VwjO3xHuDhXBjM4uewZadPjF+IaRcr
xtGyqenb6tsTechqYGRuVBK+WYwQFqm5PsJDFlGElaiY49S6uMl7+s6VQgYb4iC013if2wnZekaA
rPx78huiEGITqwbZtYtte0K/Yi1PQ6x6R7woT21k1HWiAB36H1pXTsEjz3nVIrGcB9YGTMCtJk+C
EMS9FrRPD/BFfnt47+Dh5bxEt5FKMvNyiXUtJnf27sNeEYslcx4F06zfVE++YIGuSY2AZXHtFvbO
Iqx6lC9nQqu8n1+f3gM8G5g2o30nY06hlDo32SOP6B/4XUgFMfCN81IsATKEDXjDtCq8YFu4ZQPR
ob23z/IP3yLQcUL30zdK+StUAf9PByoTtFLoLhMYH3S/SfC/aDot/VcCGx1vpLayEzLiCChYXEys
pnpqdmHxrQT1yDzW/b4vjxfIz1A4nHH3WZ90leJB2kudU1hpcb+0gDu5UhPTgH5FY8SwwH0s4i38
lKjHH43gtE4uqlY1afd7+Bo2M3dZB4bt8/vtqHihTVWYoAnxV5OB5UuStfDEXwiNr3fsjJmucVUm
pJWUqgIpxL6Xaelb+sky7TOjUDIrwMsHMlU50bbgE4FT7XcxUKdoPdArU6AMkV22F06XcORkE3aq
bmFVYXFQUQVsYxWEjtBLTamzZqidE8Osxug7I0B+JlwslsONeeaYc2DpLqtfpgWgi/KYN4eA8t5/
mYUloFGGu6lw9MUUFIZk9iJ/fHpk2lJpVzc12fPNERb1wgye0738YrWFcfINoNURIFRs2tmdxeJA
bPom52Rzp2zxwnErtVGQvZE0w75uNoFGL/erw2WU6Z0R/oCJethzzqWXnKR471zcZeNfSuc0E+wY
EOm4a/fiawQFpU0S1FjrFB4CXATw/OMu7Qp6HOS5jEYhelUVwPPaZsrA2MJUylY5QYPsJrXtmg7y
QVNHktLcEgyGPKrP/PX6UdwCsn8ztJjqWlfAxH3Ro2oLomLyLqHKH6QgL7WcOMTAAs0/5SFCfRB6
hmvycfgwnQhHim3uXJAk6hEvk3cQy6ovhBKd8TpUtt59BuH11C4I0zdasteSHrWYZbGv6eTgCUAd
EU1BrXNBadr55ZBZLWpRCAGjadf+rZw3qieNeb0t68sx4JlUmH4ktK4nDGsBzUNNtcYti1ssPupZ
0FqFgoYP/odXc5vN4VwcALvKrkyBSqlGSLQCGw5BJc/00NRlqM0FJhmYH8M49rYN8S9iaUgAwCXS
Y1WwoNl7P8lOScgiT4j9q4QewTCYfrhUPlD/sSvnAOua+LceEY84noMWuy5HEV4BpByeABuUw5fo
xMqEgVewArOaZW3rZ1AndNPes4MOWJHfQYmBnrDfS/TYJ/0dzWLrtstPWjuavIEWSJwil2Z+Xy2w
IOvykmVQMUWIBq1fc9s6n60hLuV2a4jTvdQhiBFN/oAK5zm1kNhXMlmV0iYX655zxuAiCkOM2vfC
65U01WWglxoyTj7XS2V08jispZPuPf9zVrUkrW28pvifeyjIK45R3r0cIodGSxxO1VzcMmTrlFwZ
fAp24BHdKJXAort1EKayv8pxjV0SWsp9SkzVaXve2njcUdUkherFoyFzcPosnNLrMZUhNHSN8/Mh
gw0YldlkGvTNJaiEiD1ZmAOvRIqHRPVjab8Sb/Zo70yO+k2GDW1KQ3vk22dy01bUzU30Jz/706EJ
+5f2uVl2GQsx9RDMZOgdTQdcu+rOR9jUnDIgUFWQAQgh/uTzozfejAxgLLqMVKZQFmPVv93ceY3p
aguiQ2xc9qn+LujliCoohPSNhlkGiY48rl7PbiChHd/Guz4Km1G44Q2uXEBSZIYKFnYajjUmGEHE
Fx2ncOsU4x0v8DTOKK7lOL6mzpbkifoUEBcBJ2FJf/IkXVQF/NVg0NtPUDYrSjQUawZv7W6bT2+R
ipHzCXA7QW9Nr+HByEtXJpBMPWH0Bq2+QvHdwPmTmnhnqnrb1seocZzXRnpf47Xb0oQa8jaOdyta
p0N/W6l7LhxuJlLW5hXfyW2e3M7iqUQVlbwm82942wwjahWU/SFCD4uQFUmCsCyeU4NJZNZaSBEe
3679TaIEFIBv7SKAAVNfON/CjS++2qXCh3DNGtuQLxOdzXs2njnFDNRrsZcBAU+14IbnGe3kzZtT
o/DYgbBVvMqb8Mb9p686RQOr7KQj7M+ysU7Cq4UC3OqZ5C4QddyHm2EItjDVtN8AKxwiD5rWEibm
77loG8jmxwCjkQ7vOIF+IPKzd1KZdn9vArzZPdKjMDudRJbIau0bYUHH2HpAGLHA8Ch2esJJV6fv
3Kw8itBIr6eO6txdh70cNsa2h9uzrfP1woOeZdIqBGvhF+LQE+9zVRbUoo1xhTb41DUGvJV4t+vH
t2NXPdZEVEe7HIh/hjUcIJhY+pqPhkKkjgsdy5TgjSKe7btcCGCxtWW3pkYVQtPQgro2JFZV50Zz
aZ1bPHvauKZlMDm4toDSR6zPlZJyfFwrxmQVyCDtvLab5wIy/oKWambmCzbZZZXlTzbOXvl6sxd5
NZtl7DQ9nyduf0PKdqWxguEf7omOoB0LGwDZONiDmax7hGzm2KPWGTNtY2gk6PJ7cdxpP1/4XiSW
7x8ZT5LqgafZStCSleBWUQmZzYbd0ZaeMYSuipFMoJMjTKYqNPsvTMMBWGnZyYLCGn9z45V2OTUU
kzJ4eZGe58dxKym64VU5QwSz6K+sRsBxDkcc84CE8TXJEUijn2GFw3qBClSYbovcONkTkzyNdy3D
rosNLWLP6xbiZN/QCwcs4+himqSNsw4vHHVWeVmeT2FyXfylEekswL8fqZAuljKPk71uGKH1H2XN
MWy4b3mp0/AsS8tUJKdieidzvgCIIFZlpGab8UAbE5PBup4ZJOzsarRep/KqVXGdcM6Fm1SyC3rv
3lyhV/Kp84DSGbQNyAYVv0uPuK7GRJcHuecxvKeD4YkviWscggxqKJBaHAc2zOMacJOSsaYgj5Rd
faqnvB7sXOMVkiBTqUAwcsH/HCNFzzBr4HV0BhesDL48E653hFfk9z6zKoWYlvu+c/GL6AYYNryn
hxrNzEjbS0MOaIOwvzOhG/lObPAttgUpsUsEiIIsayJp9DxeIxmrdDUaUS886Wgs5uT8nweprnGR
x6eJkL0REZLU/TduwOAOU7BgeQDh8qDchFsQZug+IGM5MzxyJwbVBQbj0Zsjyl880VhjnbOPMQPW
0CxrRdhgaz2qlfQRg7GzF/+L3v+LOhvpf4SZBDyI893E5kNZi401qHQaJC/+mhsh6wbQ6dYZRVFQ
QMspMigbtSDJpLDGRiEejQa65Ey66xgclfovxOKI52IRPaDrgSXP2gA/EVs+ciDFjugAwbXzDxkl
dpruFMOjxSqt9Wx5cLBv3/vbKsRaegAZsAAlVFLpHxgxVWNgYyox5jGhzHUAKhAh8cBoMV1rd+8G
6cssWUoTQ4o2k0vlPonPqp7o3DhkuNrhVSLmVknK14Dpl+cgv/xa5SuGYNwakFaCnM80N3OHU6Ew
BwTqhxc9ZMtRpE/oQYUGSLFEqZWf9kC1xTeLXCEoyDcrJMmU8JOesFiqyTysCU8qbocCyEuFYo+k
JqOWUGo9cC1PxZaIhnJRDwP3rmqJCN4H7RA1s0FVR+m1kYGa6bOvbh0GVKxrvP/UeYCRBjSODEyW
K7Yw3G/qYsxtMP8tTVJkBtZOPqCt/XtKasIZSRcY6eS+9uHkVaVZP5z2tssgvpXjceZWDR6RkJMe
S3riCC0TGQbG0tk8j5NRrzO18N895qYwFUog1SR/yUwy5PRtjUIbgeRKlhF1TMOTmKZDjBE+xnjr
IW12b8nxCzDGJxincuj7MW3227NcPShNwVUhP+4uOXASt3L5mighyMp0BhQXZPeO4y6OWKgrW4vl
abnFSnRr5OTLUV1VuFHuMvoBhzjc3ZI0nMyHdlcfBGeKUENQJXtjINm34ljyeSVJdsAmTHB6vybD
jq9RRSSwUTUathALaPD/BHZU0na0I0yHx8MGl3Sqt3kObPF/BFZo4dpe0xf48DPAP9y8ecubq8O7
0ch721BDBnGnA55FizrdGsH4uuw6wg7+X7J3qYJaCMolLLlmBu3GjIY7SUjLD9RqjU8Q39lP10FN
ALWGTStD4ldQuCkEMcBviMgwjFjta0XZJRw7CGBMXbuY3on7hx3CSpHXyidAJ9tSXQCnR2x1WBQK
ics2eX6h1J3ZMvUQIQ0c+6dId1w67w4fUiuwcn8w2a5nYPR7D1I6iJmFyu1JncfUrWDj0RKZoZys
v+Va+Af35nVIVQ/3G5mazm1TyhQ8FQY7R2p/KxYqTmqV2+FApYMo5AJXvmVfFIxhhz6l5v7Jh1qL
BNtRcQ1STqGlVMpQtqRSj1RfwlbMC1aHgyxCutsc3NLTlY4RIL0/rzH2zf8IIpzAqUNL3ymrLp49
YP/b+STu9Al3X1kGc6jTHo874qjrLhTNJ8Goq4lxKLE25XW131ngp89+nOtQRPl8o05SgMtVATej
s36+CT7TO2M0k6Z5lr2aUE0/1Wuk/9yt+27SOek/c6ZN+AtqHVMiHDXTWfdhbLL0CPNkUXvtdGmc
sxQi1ka1KD1f0tmc3GJ8K7uq75C6UNSfrGDCsW6UlhI6T3oBElIJI0UVRmJ3mTVKEcuag23kUUr0
gXb3+sOGbN9TXfswOiyMdvLrgqBCUwb+Z82IjXDbyA1ytA+S3QmMzKCB1cG3ARvYn7brPDCkQdwa
nyi6/bneG1BqJhZjFGB7KUFb2A8GHa5dfilFU0d1G1QCjMWL/+qOT0imKxtLmGIs2U8+YQi3AGIr
4f5jXDySRAb7Ebs4isxbs/H2sLohPH5JZ26aT+GD2X+Lm2JNFIiKpCDjYDD2aixK6h8mRjZfuc89
gypMgOrTIYpVE0aQDkxk7NsLAw==
`pragma protect end_protected
