`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
elVsPjR40hk8mJDfwhlTLj+vOgVe0E3uomir6A6iA5I8vONO0d0ZCeNNGOGuaem2
0oGlvJ9MRSeabIfhuQk62jjteR/DiRbArwMC47NVWegyKkAz2d1uSw+a81TmMW0+
MEY6VDmCcGCw9nj8Fgfx+itrwIcUZ4xcRcCM2H87Zl8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 67664)
osKzQBBIelca75R++GdbvZ6PrhDWmhqCtQ1q3ws+nSl8V87lA2/o7Cm7ZxROB4mA
yMuHrxI3PYj80aPspxUhzAEsV4VS17xJqXkQ9V+76UACwH6yoqz3G6yuS4845ORP
ObHWzLRWVF0GMop0W+JOvm4BjIs/LVL2zXZEH3Svm6E+nAXEHBNuo08KqWBZ1FP2
M7HFqZtWByrHyMmYxoWmzXq1mpKyXjFpROj377/8gZbZItkU67ncW67qiIl8RN/t
laID2hdMbI1Bj8LaogdmyUNMjMKQNuLo9W36NdcNii8Pu5tZ4FedUNiiewzBo7iM
JB8AUFvvQe9nv0NKiEkBLfxZifgttQ0ZSNPW2JasRu8r6pKtM9NGxxSQuCnnpwzk
aZlEqJPdgrfLYJ5CKsny3EpWlDbpLT50c5+Qr2c4vsl0HCq/Bf+GnGCHM0cT9sit
KXj2PKNGUdEh9gIeXVQmotkPFtSpZKiqHCp5b0fb/pTouvR/jqiTWMeudpkcpt/Q
oXUpvb5NVpaiQCVBqzgfGU6QHSiAg5orSdDF5brpU0SE7DOOYGuvp3F3sbnpklE5
tB/qPBaRr4rS6Mcvuh6fkSD/DT36Bv1XIdU0khQxcZvFmw83p0jRhoLmWzBfuGWx
Te+LH822pHCbVLEXZea46Ts2zdnmU7iMDT6ns47TV9kO3NA6oTXLVzf6Pj+Zpjd2
QbGghEJJeC4WwW2WogGASKkJWD38ObJQDk463DyT7iRpzhDzGXIgVsMcLqu63/qe
9N+L/txMlSWS9fqNJKtUMdUd+dMdo4CpxMe6lq4aVSf9oXFDpP7mhVKa0FeXsoU7
PyaZrjYG01arF7OkmXHo2QcClUnBHBQ3ax+HnZBG3ClpKW6KFLt4HfExP6Zx42Og
fIOtmrs4TNZAg5fB5NfKbigotU68OTgjkJSTQCmDJsgWqfKPzzfp2i3EyyVUs+2t
BfnPwNgZtREJ5v++67tRGNdhywhoHF4njinujJJDBww5Cy0QSmW9iGE0CP5Hd+Cq
7OG4GrgoP7kb+wD65Zt3+Vj2i4vksCpxWO3iyZjc6+j7wAAaFAa+R4jRcAKABbJ4
yAZgBkmHPizVov5Y5nLDRJN5EthFRd4iz+wKsZxm6qFhFKD4izyGiTcvJcGhQYsv
JickXuM+tkz99blFubOY5hgN5FmzBfGiBviJ+1mlBgWgUpWTBir8tTXDDmMYi61d
M4JisE5tT5A3s4uDtygvj+U89SceT/PWKcY35pnMkhXUFFIOBcOAllat0T4zX6Ez
0DPfkG5wWmDIOuurW5G/3fnF2TxBm0a5nlbpULAvVQlRn4g3b/DM1+w1W21lB7Ok
6mfwALa/R2nahEumvvcN9bMPv1taHqjlw3zW029madKd0xm6iG2MrIvHg1yLZOeC
LuSQOlGUdKCBHhuYq2XPE/SWbdhkt8jN3r7OVCAY18oStWvngb/0C6U8db1QZgpj
cr1W5X+WBkOcGPjd3mpzcNhWnFcART/7qNn3cPjqlCocRT+/E6dQrsM9dYNL9cFU
coV7Y+bfXaiCyf2p3vZDf7b/r6uLQeZvZUfJN89IFFxQsQB+koBD0YDONwCDRa6G
Agl1F1tFBR2KEegbWnZ5hBvKppxx16LmUX2+W17kxGhUpg0qYPxv9ZNHlOdz6din
iAq7q9PGR+XjPE+/8R/YZlSCstJF4uDoXOPdN8PGsVxKmPlj2F8V8Dm1TjF+2JSt
JTJ+R9M40pe9FfB5L3gAd7B4OTMHQa0a/4N/l6WZNwZYDWAsW6wNPPwZPRLKbjuL
3VE9w0wHj8YEBrxyncgvi59WP8pkmq90YrPu7sLLkhJduaQujQEckXSLeLmn9RSl
VRGzOwix81wbkHoXVI+SemndAhm1MFKg4s0HtQe0p4t9YLU8kL6fcYpOykVPM2aa
F59TSEC/4DR+0mEm91vvnKZZ4A7eqq9kyfwErhOzH3lpA2QhrXnWPF6P+rHxMdCm
TFJunkHtQ6Ns/uJgWea2tmPGx7ivKvjexgRAxj/xJ12s9puLRno3EEXRHVEJOVCS
I2iseultfdBj0l7cVClgqGt8bK3AyvacD5WlCtgyDcSuLD9hKyYyFTrTuKkxnOyF
W5OlsidLWxo/QMrN6VejFMCYTXtGtq9yXE9VzMmCt5jcqBLl1GHUy6wmdbKZFIVp
s+nPYDmv/EChNlX7PAPSgZ/4ISAjhoAf2nzLCz/EhB6Fh3Md/AB/mfmqud5UJbVp
jXEI3cOFN5ibsRs0XwHIfXSotMGBhBfQLHKEoa5PKx5C6yuNyseOgCmUZeEtc0WU
m4oIsbcBrGc6hdGd9YMahRzv7UZ/dNFKUfqtX9cq3XWObXhKPSS4xy/WH8OaCEGi
InqvX8G1y9M4lCcF8bYreIlIa8rXrhojlBuQ3EWVf5YFICblaDo1c6kcQn4wIKcX
UmIrD76ldsfZag3Hoq40n7HpI/5034ljkpTMgI7nuS8T1nfeFA7aj/S6boFu3h6s
gCADg/AqN3XRoILGiCvO4WGheTsttLUX3tLVZ2ibODZM1GZsjxwsfnHVWkk1jGec
9pmOUryjlAETaK8MI0gUeIioDVJMm6TCp5rgXkQ4kAHlU8UbasQLE/Vm6C+LQNeI
XAkcC6bMoBOut82FeqsbHRmYxS7RcjqddF/9JRcyloe9hBARZsf87Y+lrGZMZZgT
Ml2A4Arqq/MJCq6dJWIpolNt4bZEgaketIu9MgEF5TrkQYh+C1QTUtlRAMyZfZzY
ZQXtUXMh0L0OcvaNDhDQyDIvfMwNAWmZZlHumGnBC22eha2+9haL19ULNm4kM27/
AIQLMPKOwRjsGwC3oI/menjV6MAJSYliOhSrHtCi2n4ryPlsoG8iqn+g1hmDHh7j
NgviohMr58qNjtBbcgiC9NnYWrjnxt6jFp2xGRraY3faBXxYeCu6s5xusUY5c2Ex
zMyRcnCaGARmUyKk9viMgOXPtcNYlLWoUVQh+YWGAeZym/M1c97ngk1KbfDK3eBE
PpEG8GZKi9yxNPz3JtR3xxtKNSqyRDkbc/iSucRrOMDIgWwecqcinkqgUSs+O5WU
FLlCBQTPmSpUpwejHEl5Jkw1npJf5FIEjVD6QKV57+PwqOIx39028GQAbkw8RLBk
4dERp5++p/GQa5UpKFvId/mfHQjx0e/8/bd0n27tLj9safpSlhRfVfvumY0d8AaP
ajhSLf4xyVfPmTXf0GNigCfis2yJ2zAAFlY6hXfaktLsv62zm8NsqWoixFnye6hJ
XgS7qScVs3e2XKkbsllobB2q0aO0iEfw0g9Yd33YyFit4qLppQO0hRi6JOEe4SbZ
Hy5LiKn1PJKKKBQXFElUI9rlK6Vq8WznVv5uJovXuOHUmwdnkGVM+9x4ioHRx5tK
pp/Q9QYbfey65QT+Og3jTxq8ZRTKZ1hKiWLcL+VxH0n76dFD4gKQZHNSZ4PVPfrS
KUfJJfUOpPJoj5z2PGhkYIuzTGYFs8vdbiEepdB9nIQxZ5WqyIScG0dhyagSQ2Kn
ATAxXcOt4NJY8k9xjMrIHAGz00+bjmoOH0dpmn0ptcPlhuy9cyzqamLGHpkrH6RJ
arcmRdW6++14EfcLJX84QA1qIBCX1gGERq7Dw5ifBBwV2MWtQDRK/+X3VTuhqjKD
xyEUHAwn0K1HlTNOJnhDUVdaiSSUInxFGL2va6kp1p8JL2MFwPCXY6Ob5qgMOB9y
rnUELxS9+Pq4KDipp3yCIiwvWYwBaz2KGWckuioH/fhFaDI+GE6kYHvQjYKMuPTn
a0vDT2a4g0HkUOx+Ys3bz1vO3WUx+ydqFdyekQwTjEpge7iV3ZOyYUdI4kLgCdjD
1qn69ndSOemUZYbWE4d9zfqFkKFX3uLJ5w99uEgPOI3EdiaEu1QUwtHjrDYkepyZ
5f76UgTfzW17B4sfi2UNtnR9HvpURcLVBdDFTgeHyON4LQhgy0+ZJtFKvcYkLbe1
wxRqkJ7rMH36WSCBBytqOH5IiemHt6hnb+utObW+trTFcnOCteZ5fwGc+xKPTp+m
diG/nJba4NKe3GZVfH2BkqUUk/uqpG3mcL4JFMOfUZeZ3NZADPsJ1XMIBXwfeD6C
QFgMxH0Z6UQn0QrP1hYLrLwR6BWpZ8oYMRKYrH13+FR7FUw1cwiSzroYlJ3EG2NG
9wXI5/190d2u6wbi8l5BspMZrAmYLF7FKAdzJTs/xKRHE3Hy9IAZICfjTlnMARoP
PfnAUJcVOBRE/Ml4U+ZLArjcPT/AHnmRO2QiVPnWLHAPpY7teF1eps/j+4Xr4Lwn
hboKIiOpWZP+F6l/nX/qX7HRpg00wJ4mgLZX9UKICMpRYBRy0r+5FVgJk19h3emU
ovkn1ErrTlTe7XoTOkDHsIONl0MSIfYexvpR46w1FljrhGr4nkwEJSDEkKIF0+re
fzNRhzjoDyJdXJQPAevjeCKEhKIiMuPvrZSsZ+sRJ7+BrIf8j03AIHSzub4M3WGT
n66TX2LHHREnE/+9SaFrRS8wyGTJIB90kWF0nSYQECGJjp+K7k9SjddoSkJodPil
1W1HFN6YUmXQdTRSDNBGb/0V+VswWUwEj3DoAO/BISNsKGl7RH4eTFEeR4gZrjIr
pAJzmiNnvVIwJWI6J7KlKL+JBjtcjeMsetNEn1348NIkGsM9rLXFUmvzUyMZ7Y6U
oF6uqFT5AkVn9vCxL+wr9zxN+lmmWCWbdjNpKLPMoUVOnRA5j9yIAdoLStpf8cg4
S0nA2ytkf4ztlnsjITj8lFBdc7W8zYuxP3ciiNUoU7MWdey4qXAKLmzhmuIw1GwI
03KNLMBfjQIrAB68Cd+2QUylEgQwCwqJpXGt/3cyp2uqMgh5t9r9KxdM2ABvELnX
63HnGNuXpirka0oOerGqUMw2UsEcjoVeksVx10OuKfd+LTHEBhP0/N+iFxnzfOi1
f0nNO3iTgISTWNd7WdsVujrkHcyEaX25s3Mv7z1iPEWJ93SYfQZ036eoCpLvn+hr
cT3jpT2hF6G7VAyWmhsOBmpQJm2bcckPdTCfoMlqCBtcMvS1TzwpgvrFRUtZIgF8
msaPGRYJuijKlhS7UhFNeIgr/LIT6XZc0n8Jttl//zJt2R451VpQu//SgEA22+b9
tQaAgfkQKtqYXVE4o6JYGHEaztxvmJOr2Yc3A3V5S/0M//Oo6Ui2+IbvSx54ZQsC
CtYUcSlME/54ue6/lQBcD0W8H7Agyb4C1IRVUKdSuq3c/0po72++gmg2tQk4+Gag
TKws/s2BAk4Rbj0nLfsl/NTg8Ifn0u+/2ejGB12lYXP5XuuH3vS5GOmWITJQOfN/
jEUuYaPuDK/gdjxfUBidAa6lfxqN78ZrfLyVe8gBYFGXz5vEwGcnN2Vcd/Okd5WR
4m7HSNDbVImY3wIpoEJ5vBXT/njLT7/IN5RZwYRoL3zu5VavODifUT18QZ3gK+DR
vjf6gY9Nkc/SZBabGMrMqnYfztOG9tx06hJpDJAa6wtD9CBjkSMLv3U80ScVZcaa
16bCVhVAGHR+lJ2HrR3ldmT2rT9wlbv3kZbXpg89BFCFQU+ThKwSFRFZtdd5bSNR
yI1l1mtxjYslRoPscwi/PNf0dyY+MeOHVs7G/OehO49oEjMTUULD1o1ogbfXP3S3
8x7TPeyGWsrhgKFx1uZbt9mNredneH4QSwt3rr+PnDyKcFlpcJSmw2UWR7n6uZW2
KfWsNl/ElGkDmSOwbqDBP7HHrx3Y3rjQhL4qAlrkBLzJnmp6M8Xc24aBcks4jXgh
/Wj1dWytbDaGlWmH9bLAJC+QcFBj0VPu95vOn2FA8HNP1AN0+RsDoyvGlCNt2xVm
EmDhnJcSBNLaXo2EfS/3TcluMz9toyQzZOZkuhHC2n4PIxmo+Q74HnWfit11cHdG
7bxXkRL6w5Yr4cdSEUOjqgIEt1IAhPNFWAOBCrJygfveOJwCH2cvudtWqfq/oLr7
MmoUhN5HSsN0TbS9gWHpCAUmoFbsz71jGe8DAasm4jOFKxOwSENY4ngZwMpNP9hN
iQEAZCo7PCea8ev8IzJK3GA5qUdfgoj16pVQYnxN/c5ipvLTLe4PHBs8DU+JcMzr
a3JCKWrAeL0Dvn2R0Zu1ru1z1LPajL2AsL4LLSpbyq5j91+LNHDDKQs2Cr8JqVkQ
pv94mpsY5TPxvjSNuogQPYnXfkNlvPixWF3pVwjWSBzckpYiUbcaXlyD3aWwRk+/
j0/jcXzhJwjAvlR1o6uHvlszz4BPMf0dxTw+9s5LKGagTAnoeeJoGDZgEmK209xz
QTH1F564izCzwkdodWWbtg2W6iiKw2hyIxLY+N+uvsAqbm/OHDOzETyMgp6rxVCt
Y8OrXoI9If3lVavHYylxfjnxy7VVgbvKEDADj5TWsxs8vl944op0xsSKwyC/Qgux
P0VKjT56Yrtv7Na+niDpPCdUqLX77OetLDxZOwhKT/4BZZHeGyC5txSnorsLxg5X
/f5TIiAcqmO9BYJ93Da6zBu4wHviVLa3RYfQ++MSLscKBq4RJDS0w+gcjPq5Ntzi
ZkPSGo3OAjqXjYnBd37P34E2YL01JCmzVGIljhzLpZ2eOqyN4HiyVUParm/j3MAp
pOXKWYspwiLFRSerybv3T9Hxse2qAJqg3e4oEZD/O7qSMf/F7AbK03pBpjWhb/Eb
KHjzvqykLfod6MNw9xNUCXgZqyc7nLih7ALjzo9/uD4FP052wyz27o+gY2x4ikfM
e34bNKqD/q1OBOFmIj07OPFbz7Hs9FpV1p84RBsGqFoYqeEpPOF7XumY61TFA7lF
FcKp+o3R8MyY3MG4PV/t9xpQL7Rjzt26wLTI6YK9etjDPR9DLaQ7k0DOVHk7LLMV
cg48Hm67wPGs+/XsQDwHtgMYle1j/uFbYb5O/Do6u/jMYZeFn2f8DuQxtlALjdbi
nrbkq4egbKK/cmIL8Sl8EYcaKk0eBmREqOPFi/+JcH5ifEc7MLPgCXLfzC/KPjAB
mh/tk6fQkjwLeDu8xbkGtk6zhrKFGvB8rCG/wK68Q/2CHgRKmOfTwaGc7CxKjPyA
sLdHrFWN8ZGZm8CKnS67vEn2J4iOetxgCtkV0QcEZDKCJiWy56duu8++pzRHkRR/
COxQzbzl4KjZalfCOBILl2VcDsASj+D6a3vGhyx3ot60hqWjJu4fFU6sXDoH6BZx
ShRR6oNOt/NYcRKIF8kvl8VWHafH5+OaWxDZsAlAMu9A7DOz1rzFuWhI1N5bJ1g/
66dj7TF3UyX7eSTQ2Ej1jm1iqmIf1i3wNQoFMr7wz7STVN5yy5aFhjY9W/+QNODl
QZgwAojXnTfxO7bDCmm7zCQysR9IXcZRX5cKNn8Xj8lPIchgYqZYXruEs8jXphZm
Tx9OLMBVXwKAM5L1R8eTMVr5WPxdQCDFiuEGjDj1375L4ZSUfRJAf8OtLnurdnpG
V5pUtVIQ/AQlQY67wO038pDayiYw86W61FzUju7yAU0TIY+deTPx9BZhX4dk8fld
Rwy0omNKo8qwhL2Rbg2eL6l5hgwYeOYP2FpQ/LQ/uFN0V8hHKzaPa0tCx8R86QDr
a9CVCkV6B7+OLDLE/jv0L4z6PAls20jLqCyNUXVn0Un9WqlIUxg7P3CyMz4Yf0p3
pJ/YTl9/HThTtO1U63mB9BpV0Ij6Ylyp8FNmOpJnYaCJVx0t+mqqQlBwpnLtJW+w
+DE2YHIe50x2q29/48F3dD2gIO3j2fC/uAcBN09lw17jQowPlTu1gQSd0kDV3mZQ
YBXxnIVysCjx9+7BsJihJvfrYj7ze49c9I0Mx7pfLNlCY2KOqmve9Iu+tN0Oj8OU
f+XHNScubV9zXYIaNgfDdDmpcSYzlcE7CH/XnhYSBVG7M2Hz8IquO2mp9kyE/dOm
D7jsI2sIJBFeVTE+z/vfAUNO/7LR2kRAqHLZ/mxlgMrObdI+8kgDJl1qgGpdEqvi
RP8xiWA4fznMlHIMhQm9Cd/zN3jKHOjz07GJSmcb/+/FvqpChv3cNYhelkzkg6AO
DdC/w7PTcJtIE2tZGBibEvki5SZNJjvKALisCHCQMrqu+N3LtKb8xpeIdkMnedVt
oQAFY0UG3EDRq7sDU/G3q+ucKBapbzMKaxknRyirx7MqiO8zvRr4s2MMNugdzEi1
fIjRxyJm4a2HMWoa5HViE3dIlkgKRGc0Y8VPsfqJ5tHaSWjkvPKMRy2emenLW3/R
mOqfpr4b1te36S1r3dDW28paupsf6Irm3ndUSwESnsKRW2ZZabS0j5avv3t5fO2r
kotkv/K5BL805YT8EF4C0CE4ufvwMng7WKCMt8nXssMvw9NeBaaiGHGvKWjlPjkv
MN0+1vmbUEELdYQwURkWhZUJ3Y/9NhT4n2M5yZto/tVrINLhn8r0snETOL01ZqJe
nayJoXNAHAfNAJhBw2xRqKumdkkITwAsGVKGPIkkrm2sttWnHYXx3wueH1U7TUIu
QYv8SdE4zll1hGCcGgigseJIuNJS8/mAFKRn8Yf+geZ2rxJTj/6qW1qBjlHoJJLy
KiXPOmqF23jLX/m2fNftppRtOV+RzqD4smVP3YEjqsEG2DW8iFXaihr/Z9a0z70g
6GB4YA+mog66xcTLspZg6ldRQW4ym4NcefoJw5+I712L1KWO9Ep1MAuVVHVsKlqd
ei3u36m/uYtcyJAhzQcPnjwznCXXiS49UzSeijdyrhnkikSDcJHc+27MmKr4RCX5
/o3t9ZrI6kVCn2cfigS1OABQJp++NvBNq8Cm1flgRjU3OaD7bzgCbL5T3fx260gL
Pdf0dPcj8TSTUUyeVfQJDWQvJ4ISPuZlOlviijDj0YOEYNycreD4Nri6EPLEzNqA
syKMSuW91oo8gBhpC05od9m1y+VNoQgylS7xTSIyBzsHmOuugvXzqAcdOdi/Jtoz
cyalxHGx2YclsExA5KhEJRPT5OAXtvuX59KN/VbIGTTOb0sz5+9mKIoG/icPLsI1
y9cj0gU4AbcErFcCI8YtKGUls9QeJ0H0z1YGNXpUVYcn+JjhGnmPRMt4U3B6kUe/
pZMINEyZ4xaTjWa7O7ZjBCBpbnVgrKn5iZZQMKMxrJiqqz1PBr2oVJkV9+uuC82j
F7D0TKsdkBG/JLcwJ0wcALyvaP+u6Kv5ZcI/oMs6rQtHscvTuR4WAchLX8YZ5sB5
aF9+/ftSAq7vNVTEkl6YmwJ45NH45hjL6cYD6mcB0gmCUOAvOuIAyR+efg4npVX+
ZcKMXzmLRWK6ggSCm1/qJRBi3yPQoZ0/oSmyfV/4LoFUTcuLT8ds6ArWSM1Gbujo
ilaO8Y0m2+mz2DjZZFYOItK5ywyqGk63TsacTRWxf+0tURc1bY6Qv+RpRGk1bFi8
4O+0XTlZsik14zSbSwUgFUYaKLdSorz8vH2ZJN+i90t8h4eY/W3scAHEBX/lsgu5
dxmkZSdYLYWua3Z3kYncrPgc8DfOPDFCv7iCLeCS7MimBTh3RajOObfoTwD/vR2C
mZ0BZXbCxbYDfklp3vWPRlhj+MWP9Q5aW+/4zPc2viFg/3QdNe12OyN7vTVKbHrF
EAHhVGsWK5OPPoo12qvYGydxJskfh4Ye1HOZqZYrVKWvpr9MjnXeeqFswfix8hbb
xCOOxAI/+i6JcjbOx1V+jdeGyxBwhLA2ENi4fBQ1GDLDkV/68DQiwen7cCIEex5V
As7uJl0lyaKbdZzG2hRK3uyVqCzEt1BIvI9elli9Qy2YiOof3kk3mJpoZcr6zRmD
uOvdrmKh/kfriKBUxmdaot4VTkY7KMOJFItCsuHsaKAE5pQDJZbNra/dh+9ADRQW
quehq/pjs+KmvbAef8Auw8pbmQrvqZNuOJbfbSPA6+H4EsSYbKgjUUoFdHqUKSR5
TdufQTHpcB4HhxpQtaR5joIqKpWbtcVlqdkf9Y1HEZqr0Bz26ck5G/l4Csa30vc7
M7TpxHrg1L3dMkAndHAk9PEEFyU7x7M+pvk28YfwDUKSVa6kRqd9emQyS8EaLCOK
8jPec+qXCIDlHWrcrCapOOC+2E7bKfigzTlws0RCHHUmU8FepXB+XaPvw0nXsKAt
7SqQvFgwIB48nHYNutabpEf8LzANQqdTMA/0O3/IfLkgV4yUXiOtQd+FWMQljsrt
6voxAv3sgjpchlvdPGXXWEkY6vnZO1mrSRRA6dWCatG0Bo7WO6jXhRLDeadJ5p3W
QwtlOHwkgtlvJ7mLUu2xPBA3ESyokvhFNRCD9AXS1SFVR/hDqzvjGNatJ+cmtIVu
O0EDZdKIlJyNn1ZpMj2pg1Ak1HjRyVwmk6Q0YM0EaQIEoijtYXc/PFc7h+hCWdY8
UTUoHC5kDUGpkYSTXi48fi4Cskck4ws0dE9+7VKSYqFwaVi0yVYvqRkE1oOo9oDD
OT1BYCa4hrNS5dN8A7ST6ahWWFaLdjBUfrTuIJnUdtn23BYfaO+qD58gj+s/NB1q
WxgBUQZjnU4tc7rJYeG5Xr/v52d4pR1hZU5NrTHpwtwmkHwpDvoFyxl1xCFmUikE
kk1vlF5VLoCp3BxFRkeVAMsHGXHGNqgdkhCKZYYoNT4E9oLw/HzDWxaObftgZHKz
1UGrrbqZruUHgbE8jEflLZz+oCbbnsqazgWAaFfdB4uIfEEMIofWwdVYppAZiHVX
jMXJbOxJJ9qY39czLr6PLySaho6J6jZJmujNDnBXOYwpWtMAOr/wx4h2lvzQsbQ7
umzBI9Xb9sb5FSM1m6qx89YGkcuUxoj2UzxC3f01lzop0ihePhS9A84o+wzTNhNI
SNfMNC03h1cZQVJ55AcmPEd0mksE7CEQ4rOjQDnNEI3aiswDNI/UY8s7dZA9qRhQ
wJ0qKtHci/NXhFwdZCPxmDyoed78kvAPNHgrK7Q7xu0NkMqFHxEI92eHh6UcXGJa
juf6jzKDWbwrqnogxUdKTbqNH9PqhrlSKFQodavBVWtrj6BqQ+iAI/Xy/LdBp/uo
/V7Ul5oMpJ6Xn82rpI4Lj0DHIyA1Ula3r4VH8TwbIPcfeV0s52nyHiQ2TfV6qJeh
Oillb2NoVvv43qxLUlbrNxm1Wa3AnB3R1Cbpf7VZ8ahHa3Cudf3MwTUAgyDSuo3e
GBX+SXZHryXgCyDU52VmrYAgPwnfx2qr5Gfz6FPQ/RQ4JjA9NM/pHm+DPplHWW1p
LgALzRVmo5P/ywQdeG0DwI6MlaA7OOI1r1xTYEuQt6bbyBiMtZTIWB+1Rmi4wnKx
m9QlgjJywhpbTkqHly4nWGEaNar7Xg+ehTWTBCZo4+sC6TXvO0BvppAmQI6Qtzjl
V44nr9wQMCoT3ONUT5GN1yD3iH78MlyhewetE09XXXj0lzrxYEgzVjWFNv5jXUcV
zCK395YC8i+MW6FBeJ53XBsdOKr3jE5n5f6qwpnHanGN49bzjhfBIZ9RGFnnan9e
TR7g8GYVYfPzpuncTY12qrFRi3076icVSurtk1pcn/5vXCGPYKtoQS4ni5rf4EQg
svSaTNUZ5T+0S2ufLTb7tVW9bzNxW3LEW7LmF4HyqUbhNEgD3JWgCOkV/YhFvOfs
kOgDksv7ANAEJhn/orgrschEzf//JY/Aikekponf30Lb308+svbcsbd7lLc7x9Gd
NXmI3VWQhjYL6jSq1lUdR1p4zmYykC003vOU9OQP+ePNsqNtAHpbHQn0ylYnPwxv
V+xmo3DmBqxQ5TQ9eYVO6Y396RO4vpdB5EfmjgAAjBZ6ad6QmFOdioxPubzFECmb
zu4LIqZxnQ/ll5d9j+hontXfeJPCBN7CrEfOnnLJQR9YEeuyQMO2xD60jie2haix
w4Z61VZBZIeD32vC9GDBzj2la8Zrv6Z7IfEdFPweyI5FmHQErA7dF/fNOtpIY4nd
PrzlyE16MOlF6czJYobKsI754gqKnAJmrzCArqfUMdXO/C8AB17VGnfHvj6zjKAS
ES9nZ/PZGz1y5EODH9gkOLpkdv2BVQ8RpIy7wRIB99/4FohO15bmYTeOP/0VJuWS
ha1dQraAHWoVN1QfOBUOx7RJwCU9ytSRB8FvPJCfFCfEl5SE6CMPjzFNkhIEyl3g
b4Mb8OdCl/jBjtjhjTb7WXgH65OqQuxOw4WvPEdw4NbPOFm23XjcooMht70iYzTE
fiOl/n5uKJaHSUxvZQZ+sZg174GunabShUbXtIp2vn3QVr/rrd5Dg54TqGQMyVTC
+driA+Vxy+okOr39j0tP9FoVDqGlcx7PFXywJZjcW2RtYU8jMJSuNnSnhzDBcHTo
UwuhaBCj5PoiCCdZzwt5faTB9vFVuWhd89UpQqOt2A4/2OTlMWkXbY7ETdeBQDiQ
ha6/XoRdmmQ6xVCPpq1FzQ9MzaGdELrs8J6v+HRCsGRSINH/bL+565dExRQXcOYT
k8uz2Ygfmycvxat3rOYfk0QfglZeUKNbyNhpp2E5GO1ouCC56aBCGA/zRGp3F3OM
TPnjNTCQAiBCGvym/n5XVgNEpmco5RiMrWAxjgQENxtEuGbq0dLIcA9DyF3R9po8
xwMSjA9poLGrauIQO1T37eapkDX6dnqIhRN6gn+fHgJu1gRZzYD4W0MGGeRuhqr2
sh2M1Q9hLWtkjoh5hgwlMT3mJD8qMBuhzB0sCZqPcHSaMfld93z21+tzZLrwajCE
gdQ6c8TTz1KXptyhRRZSV94VEK8se+IIf0j5QIOD62FUX93r0rzhdviWNHt5vB8J
7XDtjgc7yV0yFtnn+pe1szYht4dgfQrfpQDrgNtXRd1DZlPAKdJjpRcccZTo5IwC
sHnxE/h2QXjtyDRPFhyXx74Q1XZFrMfjoxwmKHXu5F22TQfHgYh6FIQUSdiri4XY
qgDvpDIIkaIDFNs2orlcTMt4speQxqImuBZyPmKK5Y+9UA/UGT30wpTtA7bvLLmh
tsxujbE9lAoNNHEWQKLDUgZ24tIENJXHm0jqcZCuP1gHseVEUl/CVMJOGAPg6cSi
TwMdB397TwCIYAbLBjbyZbp6OpHUG0vW+IrwFa5NFf5xuzzKAFwQGXulYlTFi6Bd
XyYk4JdI46l3BjaSipLnch2yt8N/rviBHK3/8XU9bVK63ycSFy+6aTlRI6DZhxNv
5yGF6MHDeH9mjwiYw0q1NoJZcc4ih/qmhipWOQnM9Nnqt+dATuX67UwM9OY/mpdV
/cC+xIAvOuJF0vBUnwCaLxrVkZK7R6MwNJms7xjuu81qwQJZh3BOTY4EL7igkv+E
PH70q5cmwQDcBq5KNSeV24Pve982MLdPmR822A2Sh1zvndGJA58/+dKhLI5yL8yL
1VkH9MFFBMz9rm2xh5rT30PywKN9Nc37ISUDGYgkPj1dh3Hz5ig3XSfOij7T+0Uo
N6EbzEueAeHgDi2jKODc26/lrg0SISbtRnyXsMdTqNGrfts3dIoujuRCvyOkolNC
ENwd3LjqqkVByMTCEQtO9ky+zP9M9m/9H8XoZvk8k3jJAX1rh+S8+pu59kgU6WnA
CcbyQKXqIhNliR603of7S0B8o9zbGWXcNEqcQELh9oiergNtNoFTZRcSwLZaIeDb
UX6OQCZocgcrEMozQXOVacYZXk9r9c4j/Tjf7ME59IaTI1QECKyyIE3sBdMUmQl4
JT7HPkEA5BL4fY4cL6bxqJibDmbRssaaATFtVvog9NJENH4qI3Nx62/rAWf+J98V
QkJx9opA6/K0nRI45UpT1v6X2gyYogVXZx48AVEuzlKMxkADatKGCcZ3yL3AKWoa
PJORfkR784TaPIfxm2YAEGKRG0cVnZLmBuuqlm72pRZSNGn9XPsH7wEMkTwvmFOl
TOehMG14tMDzcSEFLhYikEE9IKX+3qTyhibNEZQ2mtuyc88SvhIB6ClmLvKGrW1c
sdinm16kWbYok2g0JeBHq/iVby2BR1Sr1PiPi8lUYNhCcTw9bZ4LV6GP8dxDWNVk
b8d+bR1POpa34qp+08CWXQ6WlXKS4WEvy4u8iSJJBgzudfDGHr+CUs/vb+N5934c
l6vemetljSN8k/6F+xH7OBhSkCnenNMZ/3lnlVAjBQuzpqdV36wI0gD5i+/JPyvv
KKm7tpgSQipoRyWPuZml7oQ3jpq+lpawnQVQJSp39+uu6HrQErXljf6Cai3b1Kzo
aSHYWrfYafAmLoGSh36c7RsiLq3nnW8ODJDKZjP+vL1SSxZRQcBirJHmRIb1tkAw
ZUJ/Qb+RrNp1rIzSC8bb/op6AtaIB2fI382YNRzB6qaWT4yEAyYr+9qI7YU3+xGb
1/FAmbuNGmjT4seA417zZs+Lfr4XV/YgMSCNuyAlbOa5m1hkRHjUd/6BR8tz8KJa
Z7z9TV1ByLnv3U4JbtEXMDtX17CHYiXugylMxCDUdrlNMJyRLPCUVHhrq/IMSaud
/LkJBkC9mJwgmc4INrpq7M9J/x9Jzzz4OWxAHjOsmbr6BuCA80whpv30uObZFV4q
Bo+2SjD4IPcxOYEK73OfcG9u5UQEFCxSSIADLvoMYQk8J+g9Cvq8fsV9SNv404aG
QF8iMIT6fZjB0kyIjqzxhTX3W7hnS0ET/yvsh1f2CWvVeZQD+ex4VIOCjsTOm+Gb
bYB4KXTKjyATyRm5579fLW6BYz8gsHMPDXBGA4SWQpo07lEXPUP9d0M8R/1sfd9c
uhTNYvut7l9nS9NbePPhbxe8z9s+nzDe5T/rosYHdBIabsq/HNPNT5WEm4FzW1SE
SYGwSHTj+ARrCEf10YZXvdzxKmqO9UmeDNtlEmt7zXzeJgqfJjL1AW3/VfcwIuTP
tgLamB4DfvEDdUMGaobZJV/4vf4qqPHBCaSG9SOf5YdYVl2JlSlc9QtM6uasRS5r
SqgUEE46k4dGZViM5d3fIvDroeSlYmtPTyhZfv5FtjoPXCLw791buxfqT3oeheg5
k01zVQm6h5yxLnWn302vAPlYVzwU9AEsnavpsgR/5LexPwCnY9hSvAEWOE22G7xS
o9MHpuYMbKx5X2jQJscVcqRFqtPF7VdnCRyADBqS4KdNCRu8y+0oxNcKrNT/W9VZ
MELY36EddWeerAYqCjEO6pfKuDJid/gW1IOtjDN85txRADPwPehDr8PkmdyuOJ0k
2aqeb+le9gkHNCcUi+zgwkmgR0CYcJFwg/IPwrYvYU7AR2tbnSZlKTDOAMd6DO/P
bXMq5DbHd1UQGR/R3QCO/as20ZnFudy4edFf/13NGyE9olQOqoili3nUWqm2aLfH
+fEMkC8LbLGvJ55c+RebRuA6f8aBkwbJ26wG+6MLWR6Q+I+0k4ce/x8GFHnoe/Ej
PFcRokx2helMdnv7plZKdE8On1E7RSqi/6pM7tM88AryHuxEKauCxDPq+TxG3R3U
yETY1IuefGxenWykA73FXD0IYsBJe39zgzOoReI2mXyMFd2bfVjvVzfF3NZFTezc
XbQ/RkIuwm0MKpJV1naOqfnqGznXhBVae7yCjW3vZTX9xrjWAWf+ynmw8D6K6pQ3
YUKhqXTQKVXBqrKP4Y+34jkwhXzjuAYlCIqM8QO6Q0+A1f/5kFgb724yTLYjkMXh
t8LzDSetbYgJ+jJKVjAKIQ0zBdILrPerjXIxKvoPUdet3BeK8bC4GKGcq3CE83/o
HWBkdQmK/8YcB1ZMCZCAS73juKFAMKegem9seT/9ozY95RXnlQNQA0LrHso7nUKZ
ybmrREu5/oAvfrxNLMLGC5ZChu3Ny7TUNhHn/+DiCOepqNIMwXZpCUvvfLAX01I5
WdJ+k40AYG/iHmuRniUYQ/2a3xRUiLAaIomnfuiJGrVPVzrBnnl+D26ORNyLlwVV
M1bQFZdJzWi3h7nfbHfb+ZJ1s6ucBrKGQ+18iEXCDFRwRUvpbkQ+XHuQ2DOu9GVp
GX9yBzfzLlbUqFI7gjvsmp4fhIQNl2O9ZBfB9znhg+FrkksJbKgXGe9QXLqZckdT
30n37CQaLkmKz9rdixK3HqY2cS565XZQNF1h/chPkM/GtOWWQnGaT4xKDUAFBq5i
janT9INzxDh0OLV8KxdBGb2cpKts9FupTAl3KpHAl7IA8TZAOGMh+gYGhs8eFGon
xsfTnxjkCkO3mI4h1EQwqQ4sCjJU/lYktWJV4MwX+mK+n4W40NsiEF8KISYQzImN
bB4L1GtG9ZeydOha2EZ1RWCi3hz+FIgqMyvfkVmWUtnm5T4ckOPQXluauvgtM3ON
NyHPCDpDT87xMsbnt+5/mtAvVPyvlxmzq1oB75NHmBpa7Z+O9S9uCjTX2HCnL4t+
GhzyuUnaM5CWESbOOaWD0vNNRDpszXT0n9Ij+zpdynBMNgbBj8LQvLC9U3RIRohc
8nEbxusYkIio8ssNlhtAt+ek4Hd5pBKHX5Kk+hL3PpGtIXodlY8+GH3ywyKhyIgR
7zyqaTGDxMnMjvk+n9/mGafN36DSN0SzEfNy7wIZit4xZQyVxiMNNxjNcMnqOXE3
Hs6wHLvFVBj5E08SBAESkudpZcYax/QfsknXex56C3VcPEeGnEGLVUf8R5Z0qOXE
y+Esfwk32TDKxQ/4hkcJkLjPwC1k3z1MEwyW1yukYaXUk+IMJLEZcIOGuUPBKDNg
JkU+ia8Z0c39Q/XUz7jyrJ0awjsH6LutNdctlAacZ5AaqyaXRQym2h3Xtt343nUp
aVnkNxMV3dIElBtVT8UtBkyNl5xa+I0XVrPn/y3+7j6YyYY6NrspNB87snVh9F74
W8rBmquJa3tjJq/+7CIrgTFrX0RVRl/hho4EqDehyMcofqRX0BqF4cjnH+uNridr
jtxlhy30x0akYgEa3WrkQCwFyann/uBlWREzMHbki+0iDdbobaM2naWsfJnZnEDR
QRiZ1rzcgPrVAF2HQNMDDY10B9ZrIRtpkLA4fAJte7+5Nup3r4qBRwAU/4aw+7ZM
gA0Pi9Z4ROTWrRV3xh1VN2aDR5p/UoLWZGZvCcFgN73ZOovewPOZP2NNcGlK1iZG
HcqxiSvIVPKCaKSyXnNxt++Rms3uX85w0rpeaO4ad6hpnw1SyrDAzaYcUdTE4SDh
1ukv7gS39+dfWjnKZDbnz1Jck95v+eJi/oAIl0xmhPoK44n5zUE801wYi8aConkz
oQ+8Hq+IrdWVXVXchxB2NKvWhbsM8ozko1upd4BSY9ke4QN4gMLJ7hcSd3G0ebFG
QQL9tWv/cGFQJODTRT2NrFeTTkxGvdMQRPj4SYxMoJfF7FwHIbeRuBvQNae5RlxN
pfrMNmw2CInBXZZfYNddp+YmHb1jf7Ej7/vYtG77oKiZvuDdzLGi5Xb7QIzzixYH
bEW8QXqMTEtQTrkIGJzQlRUPY7pDib5qR9Bn25jKK9lXy1g4KfwlpPQoAdwQbBEW
v1BjpinmiE6MiCTlEEidP6BO5NzWk84QfQwxBY2xkfJtt/UrniJuAWsHiUJeS3hY
63Xqs7w2Ck16koCayITlYSleGc8ZfzLPO5J5l0x3uo9ZFCLkY1vM0yHVWr7BK/de
CG2br968RnTEPdnPiFhAZbgj58vRh/iDAt22saOTSzwqAu+ybJ/5/AU1cdWoTH2D
lWL8LyGbIHwK/9P9xcwxWfvQeJqy813IcQJi3zKoyq9vC0r6iIm8T/8LmNHrmvSm
SwiVxCNrCFvXgKumBFGQu2pmFjhUPxBZ8Hoi4kTSE/I0XzFstOI01BJk4xHcWF7k
K04kEAF+D01VYSM8PImaE4JeKhIUFTcpmXGyYloSdfeD7dAbxnjlAvNqbmf/uuM4
RJK+3uWvBlSxDGmdZYDE8vlqgvaVQipAnydo05DqBXXj0fjs57kuvv/dQ1yEjnRZ
FG66peHtCRY9bfOacr7eE309HO0KcA/M3l/D91rtXCTmK17AJcDrY3RgMhUsjOZY
DA0obwXH14190PUB+fJqIsQTD293Dk+VnSJBMGGDMHLJ781Wb/ogGe+rNNBiBl6B
k/URyLkHXtewkMCppIcXow61m53vlwOWzvJvdjyzrCjNSCTbr1NMhAGvlMw7mG4u
Gq1XXuRjlgvb0CRW8NkO1Kri14j7NWyA+tGdS0SGMUEsE+uGEKqszA+/r2XqCIVN
lwWK7vman7uq3UBFOZ46Z3A75gv6aXEFIVNAI49ndDD3lRK9sUfJRLaSyK1keIRe
JFxvzbXo6dBVGm2vbqD57ypPZfMEH11nUSad2sW44f1XxnWyplNfIgDxql7gsW87
vAnaGbGt2BHE7uLA4hHVVgo9p1wKtz6kH9ys+m74ciu1SdozE2wKOmbY82DEoEJ2
RJR61kmR9XBFn0Y+LySxUQr2j9/usngDoejCwfA1FGJeIkXO6tjwQOypU7bE48i6
qOL3Zr3GK/GS3Bc1QiKZ86lsTQfwOFVo4V4xUqMNBkd1UXJ7AadR12/6LTCt2JMT
eAnZeCT9oZakwwRmfj0B5XkNQ/EoY1Y936GfRw2TuvIFdyugmOEWwTbSQDD9f5eU
Hm+/yhdZsLuzWMypIeDG97aERZuskF/jJR4B9CscyOMAO+nim+/PXnmM4XU7/Z9U
taEuwBDDsS6KGvpPFVaBNs9JEHeK1QhiTPPL8V/B+TEkbqFkgANs8KwhpshYc8wG
HViiWHbqJveHPW1kGZ6qjoRiyXLTvpnWu0R1zRPZ5BHg2YAockW0VtYvjj2cP7AU
+wLbBxLZKWVwvjdBfoQStTRoMC9yyxH2QGeUGWuOYzzHShl7OPN1pwY/oj8e8csG
GEfFuTXWg7ycrp6k7SJhcFL25K3C0UwPHEeiB50OpQdFWWQk10D+mFYEdhvTSV3z
rdR8H2JJkKBwY8wgoDCNXXkUQkqIGAeR4YBJbgqOedWW+mQtdXOD3lvLjg4rsLtS
H5Tea2w0UGcI94KaDzSanmkXmFGehK8fAUI4cd+F9RfkHY03E5ybUXBqBl0m5+14
dp1MKgsTs3cWYcSt8tkYXncSEFssrWoiF8bCgZzPy+z1NcXCPg51WP/JqJzsyizu
aXXnRDWnNUICCop4pCFUJtFMalznmtLb3eqVLFcfKbovze+kDD2Eg3S85opgtuAO
yWqNzhPYNRtsdnqMRCj/WndpZOtaJmiv5xmzQFVCS+xsmydasxrqyZ+fh470ckRt
TaEr0lDcVfD+ZTiJ6QZx4WQXUIQYm7Eng2Nkv57jW5tuVhfRsJ+twzGWHvToXAhA
zQ+XUFpVMbdHxa6gNzj33yewzsO0Bco+pSYg1ZzGyoZAu8/SRSFxlrlmgpQY9Ova
xs2u8YQdN12pLgFwPV6CfyEARYOjklPXjzBl3+GCN4jCod5STkSzFqf9o/Rxo8Rs
AbJjOOB+IMYTouOQRopN3N1AS2m2yJpeWKuUmN44gE7LNc7WVP2F31fpTBxQU75b
0qnmyZzPmWp2BAsSXcy/WA7PVVQsd+RXeC3hD4RCgfp3nL5qgKiAtXXWMt5btQwt
imJg5zufVoZfsjCWWtSbbGpajbau1sosfTWJIm48LTPtsTSLHjeXrCvUxOvrijSB
6VKbythwQ0hPZQ497ohXvT7cKo+wFt5Na5+V6/6jjfj2Zq/svnNI8kaFt0zXQZqH
+Wwe3QZVovoskvXMMgGuN0jZ+JSfP0bTe9Xm3y66nyrMp9mIcQ5QZL2HMw/wO4sT
u9A2T+jQUxJLYkngOGg31dMmHG/MNobXYkeW9JJnliPEUV2a6fu4KygKlC43B7Oi
4j+mQ9Q+oRt20diDj+Hh6VcJoaswFQLIQcC9pgWJ0WKuMDk3enPOVIFUdXhdLqIn
pwIXRFJmoSZhNkLXTncF6751iadYde0rg5I0cL6j1h5YE9oEm44QDy9zjPyQBCfV
3/1YqwNHs7AcIBBLTi9uEZXFFA8xX7T6p5IWow2wYKtDvgTgpPdFhDG6mxOME4bR
ORl8t4Oe4+NKqdL6nS2B9QP2YDs/2t0kml5siRjH15iYWsQUPFV3OFqQ2zvVI7o3
30j5F6XKZ/hBBgjRD1rcBkPfybHMpEpJLZbMlGZx+tB4R2RO7NwP6rt2ToWg3aeV
Zqw3kU5hfYXFQfqvqmFE5+B4mewtapObHc7ST6h4LcSWe2Y8Wwb3biqMkAVenELj
VujGVuSIJ3du16AVj7/EQFMm9ngOlvtsHvbywK61a/adRjAYZ6uiUQ0m7mHZf9ZU
wDe6Uj7e9jlxAxA3OWIWLg//LzpgV4jrisxVcEO42+uMb+WY4XSxD6zt8gsHWzOi
el9j/DmuZLG9oe9txSRfuG5jELhxv2LEwgiBSfsxi21PI1wv3+CnyBPEWOd06WDp
8XZKX5UGPtQ5LEcKOzJU52TLhlLRoUVjMcHO/C8owTzb23Bt0OIFhb0FCYC+nBXj
U08ya9JqnrcocYJ793AIuf3gV60hGIoikrG43QuWI9fBwu06K9/OzOKj3E7pgDyP
EdoIdyhT3cjfvH7MnCQPCDTSOih2tIlHwhok8re/qVZaoQL/rmNX7qsuPnMj2Hwn
/T6viywAaGhAXwOqgUtcZDu8xRNtLL6Y742RISBwheUBSGJvE2k+4yIXp5CC5Soo
f9b2FYnjayuiJKqmhivF1cAm+3iuG3zknUJ+Nleu4FTDYnHhUlReIhhte0gtgwv9
lKl2H12XzZA4/nB17U8YLwbpFLmgY4Qrs20pTYDyUJyrRQuvk7Av60iQhQCtpvvw
6Sp85jEsy06041hcsmJfIvBYDJEEkK8GTJz6V9KfPHRMWywd3RKPgbScF6HnX2sC
1djdWPLLET8nT1QRVbWHF9OWl1D6vySimpuRYHnCHoh67EdBI/oLl+cAJjQfBXkT
YA/bixBDZd58wQOduTquFkxo3PZxqI0Pu74m9ArNbG7Zar2N1ru4B+y2b7qmhZnK
m0HWPf3dYsoHeW51CfynK3AHWRdvQKgJ1mekAVFNNIawuBk5e4ivBXgQGuO001iw
MDk5tmtPjZRiL+Sl+y239rNOxVlK4m7BDZfn5nLFiJXMUvsXBEkbT8jiInCXZKFh
qSdpHl50rr/HNPKviSbP0wy3YzQJBSd2S6RGAmMgZnq5H/GV5jISdSQVHmaaP886
3egeaXrjBsMbyqt5N9YMsBO0qqah2Ty+iJg8mLhUU2Lw4rDQhZiY+wBSpFexqSl4
3RbYdOlHeA0QAvnCJ6tvIsBwVTUPXp1sMNADVYI5GRaehsH93yJDMR/1ncL+bDF4
TxPUF0sUyaOQ5eKjUXlgTfD803FP99znz3aFU+SDxq1+OWxqs5IiECd3f+ZiO4Rg
FJzi3dMv8b4b1SW/vo1YbVHSDqBGxvpc+Kh4ytV/Z9y5Qcqwc/C9boNn+pibuQwH
e419nzJVvEbhJmL0AMI6JeUbLamfIGvN3e46q4OoYEfiZdZ9nAnrp284iLOnTma8
/MswF09bQpRb0P+NQFE/9V2a2pxnFkJ9y4TIVE57JasNwznPwsvUPOhdA84+5C1B
YpOxBJPio/CQUbu2MLe+metdtEjPcn9FoA8CqUhC6j8W6asFhrd53v1L6X5yg2KR
S2iI8PnpizDdppfUTi/hRX51TjP9roVP2rUoI2abGE8b9gJdhfCz6Oc44TuRLS0s
MEu5aOtkDRpSS0CVoHhHinRf/7GExC0ZgWC0WD3Zt3+p1IhZzVP7PSyjF0Q2G/3P
XxWPDoSfFu71RR4RfO28DglZKqTsEMD9hX1PwU6l0alRw8lLicAd26oDiVPvWel4
b761beVhhYrzlUTWSyg9/pHSd3fzgrjlY7Zcuy9482Me0TTMiR1ZCSeRiNMsPnLx
j9T/TvarcL2RFB37reDfPCTImpDDYwJij6INgW/XwYVmG2SBWSSVn6DxdvcxNZAX
YMD9XToJhCCDqEm4u97sT1YVPIYSwgCTmybo9KHkeY9YjnP04W38dHBdZKE4SQmQ
Dw9K+QbbylYRjogRI2T8Ndoxmi8DU/By2ytLZOZC9nsvIX/s8VCBxazZxY92zecn
gJ9OS4gkxPMBsB0ZXwfxhDdD8CwuzlLGCkygF1+tfZI1SW6ypqmSXaFd721i2T7T
By7hWCDE/Kb6P0C3krOgxpahNid6J2r0Rp04D7Cj5dOq5IblIGu4LI6ju1BNMLDk
6rgr6L4FZWfQh5EgrB+qOJ9JeLGHley2dupyJjsw916kPqBheokJ3MOm2gUEZdt6
nXnGBs5ewuui1b+jbOpn8NAaOg5UdtihvnX1QUi87/NSW2pL3UYBRSERTM4c14Ur
FJwwbghhAx36W+xYHZA2glA8QgpQ3anbYxien8JglXN+zGbHFsh+PP/96Cs6gyy+
pJ7ZBzWN5WGaef7ekVpnzcQsr3YxIt+/pQJvJ2hAF19xGCflhlMMhpAHyEaEN5PM
XURp/HDm59tXAY1KVZj+SbtxJnGfOOxxLnrB/NUnlbjbpWVTIt1Ww9wHskw3bsRM
xeeFVd0OLBvtWOVcsdVFC1Eaq+J78viCnf1HbbTOrkaR0vEj9hwxDSAB6QUTMimo
W8i2o9Jpr3zL5ooJEVtqhdqyZmRs2kdDXxXkLSkSx6u42mx+RVBGdnDk41jp7W5t
jNqpRyfq2+nRW7eY74ioKaz4XABC0jjazjthLVIjTCySsTG2FeU4h8go2CsB9A1J
skirNIrjcPdgL1+pNu8eFtb8y5FJp8c86CsDqXBrSefBNpH1JolLh2lkkzts969w
WU5qnh4obqtolHbY3sg9lymoHD3jE17VvwkAGpR8fMUqBo2C8rVfNjyVSgFegZUx
SDOE1dqpWZ6sMYzNd6eFxvUnNt0Gs+qBEUUYOor6Ki2S4rqhfxF6CU8NJvfeKfLg
3JzXe/yNPHXaJiu3qvi0lHMNkOXliHCowYctZ8eYMZoSNJOS/0dXYhiEcYYP+14x
vnBhXObopHmhjPBqOX5CN+ugRhy2J24GsGp3C7SshugORROj17AdIqCYPVoP4HbM
tn+YK8sh3mGbc6ppXv053absM76JqK6qVXDK9VjKoxL9O1algoW/WZrn6ihLdzuE
aIPbhRiRAGyBjhjQU5U7G4vtx6YMaVGHvSz8WzPI3GxoN/6eegb9emH0yZqxmoLT
jKf4JXwXirFEseSozaFKACZWAPpnxK9c4wKWjZoR4lCkCpG0FELiGaX+Hzk1wfwk
CKgQ7dBDPyUFm7L+Idu881HyODWq+1Re9QYZATu5Qv7ZNGMfYgT0lKF53OP2a7/q
7zh6CmUC1QzWphPv31lryg5h+L6fcvOgm5IyNr1ksFylR7UlxDSAOpXy9aVMDg0P
mZ9N1CjDY2MqFpeNUll3+2Dj6d3KCFQvrHoMzi8oAq4VFomJZB9CIQZnBiLRj53W
lX201M4yNAy0hIQ+GOLbIh2M0gkLz4vsySinwT7eavytPdYzoITIRSR1OOMql4UD
Q3tEho4KR8SfiCzI47Dqw/EH6xKSkps2XrPenkJivqsW18vnRUywcuOrmkStCQRQ
CvScpRKlXIDF8VQ3VMJHEElOBQL8gOXOm8OoMWCOgS1nLtAwz1V1ZSd4cueYgkx8
AML6SPzr7c+APY2X7RfZ1DheTMvLMQI334ejLhQvt26pLXqYo8eTDtQPWDR4I+89
V1KRB+GPkXvjRNlq2YzMswAJSEH1D/viCRJeiObnZPoyzanv3djW4PtFr2p4Cdtm
tCDgJr06mS8xZdXIYcBoowSKeUqi5hOHUyhd7gM7Rdiy2wh6DeQRcGtos1ofWsB6
Zes2HctLA/JTdzmjFe+WuJHX94gH5T6bODLSm4+P9/LkWG6SlYPcMoOizixcaIzF
QEtDgShhmwZcdFykwBMEZW/55Jd8JsJM7u0EuHrUour/ZTWpztfz1eDsND//SfQ9
7Fuyv+gzHMKJeVGCRL+PqJFxUtUFKVzCN8OlGPBJ40nzQj5FxTxdtAcO5EhX/Kmt
YnKhRiyyJGTiLiahun4JPPUHa5oJ4nz8yvthuvlG+pa0iYFgFLJx4GFV6Mvetloz
P1hG4BwaX13nfM4vwtadHxBGDmsWz1N8YjowxOjH0VJgmUcwQlThioQKIKbmxLBl
hCILuZhqws3A2466yVmPg9iPa8eJQYRCzwFSAM9Kb72uLaDPhp6DlcL2m/Yiwnud
jsbImuA7sVb8Y2I2Asl3wwxppJQ2jxTxSbrkSFU92ileSciNqm7mB+X5W+9HTLEk
RT0wmpeDoX7W4eAOW/vnzYX17Ov/oA2yTDpkpSwkDogOEXT2hl15ogu1OW9E/UAo
sK6QYp7q8LEciWtB/f0cW4UpGtMOQRQRy0MoMHl81j0cPERfkhnn5cj9gJeLHL3r
ixcYww/qmIPhEyQU0EVe5Kk9+N4374NdygAFWTYGrjyJMv0P0lPqCKHqIGnoTf7+
vxQjb1vb9comJ5gdJOH2WGLHt8FaMVxFBDdmKRXxjenIsImkcatbZ1yrAj9A1ExR
818olqhZJ7GTX4fsPGetFW4KO4rRa9Dgq0D5z2kt4d4vZ754G0EuApieb+FbZ0Uy
lSENwXBTJ/av8RAnK/eexQSIROE4XNPVeAS/jGdyVf79mymRQSHFAo0EYr1ZIiQa
+kb6m1fQIj1jqwMR4LTEjOMUyliLfX7z5AHlNXoDtGBVyZiuac51ARcM1DT6tG+H
017zI7S6m2gzKyGMsovl5VCl6q2qOI52SP4Pv5lSbSWUlNr5kOiBIqB1gpY08XqL
BrFU2SStQy9GUEV/N1ZKRa8vwLUFN+ad7mE299o4ZuQUzsKWficqi1Nnp3T68Mh8
vUq9acIQYx8W0omjXF887wHFUbyAuj18K+kbR6ZLG4jrOueNiGv70AUfiXXvEepJ
E7C9YyBjpVZ+Alt//5Y5nmEN3xGi7CNqsjCV5qh0R0xG6bKsHjG9Y06j5WSMe1Ci
P1y6Darl82OIDlpjkEVqnHfOwz/+qOo+N/LebUPMDfEtYrqBiynzjDcjkFXc/cKr
PxLV2WePU0QrTuapmdrx/XPjH4vUz+6QeVWE1aFVPn6MBt9qhOTVeEBCoOBoy17m
eQLrXBMgcxovxXK6xaDt14UCFgLGvAD6ccd1D7an3b8/4FdS7AdhYvC1KB8NWN2O
kO8exQ6cCozmTDxeSdDQJGuDBoKWvSCNpNzUcXnme9FxLMRvD4daVPcF1b+9D1Am
BfviBnHD3Vg/BTerbPtR/yi83AvAQxqPr6KQ9Hma5QEcSX6r4riuk196SzGMDPy+
949pY/4gNzbaB0mllLFxOmoPpy78VbbVnxzbeKl/YctkUoHejjr9ei9bS7Kts72C
NIdOEIcIk0PbwM3FxN5bWUMx+TDTpHPzXzLl0DqrJIlR3V03GAw6zYm2qzEJYvVu
LYoJhA5w++A49TzPJRjvLTnroy2wIkWNg/o9BstrLCUPMbPnwAr5cqZYQaGZmEJN
SY61XvOdt7lw7VgoWqnXyvtXPKNuQEPrwlTlbpu+rWoQWgoriJjQWdX+Jx5NiGjm
x9CfHO/vfbMKZhvz+ukWgGHvjQyuF4IX0FMR5mO6uvmXd/llfmg1+z+SDtYeeob/
hd/Ed1nVrm2b803iTIOMUM1Vnhr8Fcc5j/ZQagRO3nFm2nghfsRbXx6dCt9FeuBP
GDifRYinU4aLlZ1Ed0jJasYpLAffeeRzGvxdiHraCprV07W110Jm9nWxAeJssFfP
PcghCindJJBNg429fnsz+qpKb1SzwFhEVBJyI81TinY+VZMmules1y5WRyRwtAzp
duqW/5B9xl/BNF+dvktUMawLh/Kdf9KkcLVMCYZ+EZe0U1jE9ayN+kYkoI0gq9Gr
98BnT4cVzcwVWY7JH3aIYeDdCc9yaNGZ8D4SY5Vr7LOpEDc+HY4sXNKDLE4f0V+O
07goHPedJTrPO0nl+1qZrql8gf7ffIrENNVqolYujMCNk8MPEPNtAhJ/9NXB/XcM
o1JwnAV5WJjTP9MQPZn6Pf4MWIUXyPe7xDuR5ykVYtWKEwWkKb965F4jWd2JqUP3
FoCM5PM+ZABMqX9hVJbrbt0xzzcvuDX1v5uCcGOpR9ex0zkqkVz5d06EB+SmeO1F
qmdcVbdvGZ/IWxBEHzIIje2qkG1nPkTsVFwljMOCuur+4OlLvhGb44FnymRzW8OH
e2yWoGIAoh7CsocUm/kpGUEwXpLSmq9pJkrkSFB/mRNA6/9Ed6nTG4kxHWlBIxI2
AE+hrZCheunTkhZMwpqDL6fx3P62pWECyyhSsK5Ssq+IQRXpLMutMEuCizn2IhXe
UMAo9vHa9osABAxuJ8PNTjtSoZgJpE0RLCONJ1AXXOTOz+qCmD3cboXsnFx76r/v
9wZ/wmKnIty/HSrNDdgsEi6dOJ5bioDIjsghVD8wgizBeOLwUMIWrrdVM+pRVX36
jrsuqhER73SpqEeJRcJHX73zVLC5JUi8u9B8xHDu+ACA11oyPhWJYHqKNVWBIsl3
QDx2WHiOmZD/b2UFCG52rFHDK180qLB0mLOwhowuYKYPEHX4WjsCDkmYUDYuS8J2
e6e/5BAl4qhBBmfjr4A1SOMe9zc2hiddpsFUgPdJ0p0bhGTWqhwNahEsF9cch7b1
TKfOMXMGKouAtMnj09UkqiY/jDZV/sUR3w6WSvB2fnjL6f4cNB8HzvvtqAZyF4r8
GWUBDMce/WKW9L7N+MnDH2Yo+rPGxlG3mLvWlIt6DsRM2Mmw3Bt/2k9wNKxzdrhy
Qnvba0QcNV89u7nWTf5zzyI6HwXgRz+brZE0IV+H5R946b7i7FKtwxh6uR+xxrT3
zu+Twsry5iIHvMtQBQDKnih3W5tX1LQkOHz8tkLKPHJyaKJJWc3HMHxxFHS2aohn
0gMUCEA4GP1Aq4NeC94RRRiBvYgfs0kXmGpaEyDMtmQg2PMc2GYbVaPeh58l6NrI
V9sYYEtWnS5jAzXKXjos0nUqgsoF9iulw8UBft9OPa6/G063kcXvlnTg+8uTEgo1
VbWGtpv+RqkuFfZgSTgr8WprZs5w38LCtuN4kcz1hD6RydumOaZTE7whRYvBHOPT
QWJXI+D5OTb4Nys7TQU5ePqowVEqVR24rekjdygUrpepisWxmF638M/g/1WqU1UP
Eh5rtIwN/x3WIVXFFRV4vFp9ZbAPheulkagHVSoVxPoLWIGiGl2KLR57S7CwSZMh
0DgC9uDnakA9eKuuWnsiVtRjzQicNbFLIUBaRrigxHrTZCjTU78nCgIjuB+b5UsI
/cB0GJMc6rFWy55TMNBMRf7B6yztJKKoQ7NneWtYBCWfnapJ5Dgzw+Mt+H8zJsRl
s3pDrP2YypNMFX6qVrq9tZPOkVORMGXQlTDNPQQ+//TPbisRmWu/6G+unWcdUjVF
eJHeAasyDBsQ9ZbwCUPRspdTp1uxx25A8zdFOMY0DgkKtDHdpEzvN1B2V4q86uyK
WSZZ8lE8rEpi5YNmvY+F5zL+z+x7n9DymSFn7aI6JgfsoLXqV5gOEQTEtZ/3AWRe
eaFjcrC9QAgyx6X9K9m7KvrWgob6X6KuBtGvflHkns9orGpiWayBg8EbkI0gX9OL
/bHHdYMIsVtMJ1d1j0aiL/eL5bG9VT00HdqLTDjj6JgF4nEugN7YfKt9IOTmPNWU
pFRmd1QBV9H6PJxyJROWtOkUJGdgCgFWg74kar8rAQqhHAx55SFiQsDsNvbtORfh
uI6ZDEtRP67BAI4gOmKpoq+jkHBMlL4aHTZGHSY0rIhzWP5JSe0YnEKHQtufqFO6
auiqhiyUC+OWLklVbqgfkG/5cPVgnZrHehBsKYE5dGI0nbm8oFUekqNIs2/9l9v6
7l6ZfRmOo0QQkBkDzMAIAVMuwMl6DNWNY/SbIpDohCkOU4rTDqSdUwytzgFkvQg2
ppaJ4bZ9PFthxPQV/AgJRXku5urp5Amoq0s97oLH7O64tCCnZDAzaQjaX+Qkcmhm
sGziPVGc/8aI59h2GnEodNRjNbjhayXJGyeZw6aXWEmGENyT2NX/joDS/9iBojEo
xtlogNRs8Fkf2GN6OcSaDRuk33/ZFnaX6Kva8XX4N8g8uwdAswFb+W+fkV8ohkLy
G54EneB+KPhUK3plvjcrIbSvpKXWeZbKQXD6QVMkle28+oV55flLxCw8oJeBPf8L
o7Qy446pL6SACTDt5g5rlDdZR3DyAt1SZzltdkl5YPAgM9wQh0nveBU5nz69DTM3
BOQr+mQ/aHv1ho2M9i5L+sqIWLMfL10KZbJcuplk5QUx+/hrwSjaYkww1n4V3rho
b6lAvssy+t9Po03ZSXRWv3LfUzBkR8QSbrusYseSiw1v1due5uzjj8QPty8q/rCc
LLnWbMfTaTofcA0Kkf0ijP2pSZbYW0Msr417hFxSfAx63Ts2TbuAeL/rc7qJmFWu
RbsbR6+BQPoRVWa396vB7WB1zPYI5J99cGzTwCrn4CjXQRXhwmkYtj0wsmJY7JoJ
m/xRj6nQL+hDIX8lPSgPxboNqumBCwqMR3B0H5qHakmQPRfBv9ZUt0Qqs0wCyQdN
sbHgC0LZvcjx2gOfFYrZl5jDo+zVFz8uIAhszskSVMmKA5yiBWRi5sTEbmqTu+Wv
KL08QIScabjsAsccQUfb9LuKHVIarC2OXQ7J24vfaYo54XnL52YvLlA84raKjpmS
m3bNWPLEUG07bCbIumSrWyJDtGv7Kl5n7jXHwJJVVyouvo7R18zPiJaTjorAujPC
4QdLsbZ5up/g86gy0UXAaZEoaOUnt1iCKwX2DQ3cRxOV5OkXi7U2gKf48gk5wrUZ
q98P6/05gjmSSSsikDVDiRkCENwxB3Tfihn6BSf0Ymk7tOwgK0mwog36oaUHB2zX
dfSmD/UV0Cdyfc+mc3lNMKXFauzv1tHDoEMyquO7k7aVlbkL0U5IvwpqQUX5X4l8
ZFXPn8y94ZLTvzU7RxgGXb9/zSDEXDSQENEA7lyCs9+YJpb0G1acwThpcGYuuG/6
h/wa3pQpbrLLinKI1qkflFpeb627LxSPyQALiqXs8PcY10E7B8USZ8h5UPlgIIO6
gjeT6moG41C9SfWfvua2IiOJLf6cx+ujfIjmjJhdrFOXyjCpLJXq6TgxCwRTEJ6o
DPhDthkD9OANiIV83SPCC6oKmdwcZF01paw3EIDdOHG/+1WoG9Irb0toImLvDJUv
EjaCS2ZdynwngR5fhY+g6o/vGMBpEzZ+GtVldWyqFlh/wciJHZWS8KR9Y387G6oD
+ukRAqx65KmdPBCkmiVvy98A2rxGAIXoXZlZYFmPCBwWccBKvlLe5kTdjzL6AUBU
KB2cbTaWVP+phiv2N9st1Y2DvdBqYHMj5LSdz1cM82gX/JN9XNCcEMNbxWCONEjw
eO1/dWx4OA0ggcb5/GjrzE38V44yrSKduDkKTErtOABr6ANQFqpmLnyqugjuOMV7
j4hX0fDi7RJHVlxMG6wwaDVcLXGWeUiOKw3CApyTWu7gf9+o1HwaCyQ7jwFKpxsZ
eK0YfLAs9hLjViRYfv/w02Cu9DdKx8KLDi2id+vkJyI8getu7y0eqnkaQ116/uuX
lQZtOiH7KqZu5l5aP/ip2sCHKR+esxpN7jNe1i69FT8skwtgBKKvz4TvPTlUq/Ia
qJZpC0syOV1kgStmzB5h9XJg0uuqFijVB/r8nWOOtT+eBONcKkmPEDkgI5Dt8Gip
LWBcBFZeU+Jj/4ptD5rMVT1TwVOc28MBtH0Ks/ZY1YYUyVGU/+EfDBlBlcw19VDk
N+xYVvH9ocL4kXvAL9U1DZafCoZpdiOG++pk2p8DCvUkY1XotcQnMsutnY5xpBN4
nuut+wprCr5nFn1gpAvn0SlRn+nw1fUwNxsTI5x+BpByiJyXXtOtvspGoz4rncFy
mRcW8nq5YqM3VRZzHp9YbxBVjcxPZjvUHrDqd5Kgli8lwhyiyNoTxPtKSmmGf11f
1WhajAgr6D4wclwibKqpv+2dRLs8tRVi/zfrDBUnDOrmNyDOHZDd6yCv0O9np+ZG
+8JPbSxqBg+E8Gdye1nflcZBtNQ9Gg7Xp2GIxwUxK7XeX6R8S/rLu74ugXeIYtxT
/33SH+ylw0u4Z91bUbQy+X4Y+vjOvSmy3FFWQMsJKJDHxL0vbq8chQKtVKxyImL5
lWVEF2VYNRlrkqd9MkWSUQ0NoR5A9znxW+Rpevq+69rb4nnpmv+N2473Pr+YveH3
oS62ez27cMBRPKfHrxOgVx5eenZhVtoViSX3SHysvyCZUV21Zr1ORu3QMTgSj4j4
ivj3C4Aw/6UL+FmIIHSEqQ2V3OQl1Tg1C/lr1iKOtYwFbEIbLTtD8qCusA+dk0y3
biXz+bib+ksf8OJWolahimLqFBQicEt45V1mRBnZgoEwj4fqLi7nVGGEoupjqBNi
etJhXpmt7+AO7f20p+BVMbjkwAD0vumL2v5mZV2yeF1VI+8y1aqLCq8w06Th9Rvf
pbPON0Xe9U1FjCELpgYfsbiuYlxkc7CLJ/MVZR2BjD1FSTd2serwfMlZZ9TSExgV
sfnmVS27XUTnTKGU7SFyLoAOA+GjAdmXARGf9HMWXbh3Bjty76sggDtg5DvMZg//
CpDxkxD21lW0z12uYjakhSNHmrUaHsUUlM889EVNpCr7nmZCLjIE8QYTnDQ5kq21
m4nI4znKo8pAiHp/YYX9ZDj8lYkrpoN1ZDo/Lho5dwwlkV7LrFkrGl+B/IURPRMZ
FWnHUbBdeLy7u9Jii3rna6gyXGWMo+YzHDhMHAAXO1p6TLCj0iex0wlUYs+ZPnbw
626+1O6kekv+5MwWwDxrLeNqLulCrd6szipfwAk6veVb59hWcdEGpeA6qEW5rVlS
W9vKWG4rJbx488mqRzxsMuTemHcvvzIn84MHayx4ZUl6RXMvi6CTVitGJJzZeBfE
v5kUfWROIeLt2t1yl628GSmM3UKYwQhBqZX09gfwJsb+6UqkNqwDCy34pRMTNWG6
Fhe+fMh4j5WPdyIrSndpIk1+oJWg8YA38Xa+PIF4LzZWJxZbp/4b9QBiCbGCaar8
auWH8mns4CMO6CLThKE7rmkqaToKub1EIxXpG0Bj1ExID22jfia37XhSrKYV1mRF
Dth1B2b0qt00A1IzHIoGZGdZxGohJUouI5mO2ZQdF1erwIcvmaD13AEL3UQ+AwPn
mzi0qNBGINU6/5SICfhCZSMwBay/NIaZs+NjUl3uJ/BSir+SPqO619lVlklBTry5
oJKFsHO3AcpRNy/ECu+8cVPUqheO55flPQUQ1l8GIoYwAEgvRIeZe37mMm2qUwjV
/goc516lfFVBt1WDY3MsJ3lPakMtYeDe4D2sA/sTfaLkHX0SBXyO+mYATQVmO8pp
uwF+I3W/AOuHMjyhdJa3bQH/y6lSwCry8GiZkNH/4Mn+Xjgu53GkvvZ/vg18y94S
FoT1cWlkgJOB+/JeXGdakZBpsPp36WzcsREPlfd6Agztl+qXya1kNv7BynaSI4zP
h6NRC8ETHhehog2KH3PzoIMsfbNHlLGtI2gzp6pZk3amQY1ADFtnFC4SpgqpDl/l
04LiJQ1jSaHPJn2DtWWcqRyoB/N/QkSQRBpmOZipCZx3JUiNFC6GvnPvpn2ywBmB
MpBzipPB7pqJsSGHmtL4WURpVbYykGWbkd0xxmL4pryFbdDDijxiExEGmzJCHPlo
93uwtomj8BrUof2pfH4c7HHI/Drk5MP8t22JmtSQcxFFX3ZokLTvsVVEqQplZdZz
rOfHcQZwirAqGqQTYwLWsLZm6sclzG6YI0Pz/CSqWuX5cybXJrpfIhdLbB59Gvvt
c2U8KmxxwfsumI9cjNew6rssq83bW2cIDGsEV6WF/f/EJeXda45m+7YhH+uy5DxK
VMzWZgWByspdiZfjkh4FCCM4awtY5gsXiFN+nfIxC/uvV5vMJFQ082ohmGZ5EKVr
dBlS31oAbANtO/rAB35bohaN23UXDo2Koc51uaGeh4tNbaJFFS7t1oGzzZ87lRLX
rqEqcsM9Aj8uFQpuovuda+8qafJYKcdBASQZWztRVKPVAFkVN8U5pqi8K4B0Qid1
VpPoj+Fm3PPEp2aKOPmtqYBT/Z7aqpLPUOKWhmDXNu8llcr5GJxjBX2xyrGuMglp
18Uc26/jLGzXjA3K0lyNzZhyRYADeCC2uruPFIbfC2olhpVhajI5OTrRUXKK/6xY
+9HMzsEhadoB31zwhX+lXtAUmeiiDxgyTo3bwKBuE9PVIgEbIJJsM7NezsvAGFw8
1ZqHaIrGU7ljSQxS20ypOR/vuyeqIesegEF9cFOP9aNUvXiDUe/KpbEaWDQfvIW4
72u0GWqb8962b95EyGBtsJMWeyEclIpP6wS8i+dyxcCjq+9DKA5OrhpysrvPJhDP
B0tyMPn4+YeC5LUsJnp41TdGJQN1QxAisPkaJ1eoImDJcP76D08UNAUbxNN+95P6
xouVXADfIywqPHPFlI0cnI5XoFCRt9SbiMK+tP7sh6NOB9QeTtN29JFdafKeyqfL
wOq7Bf95mj2SD99I4E0YCiw0ZqhxOBF3TGel2RX5LHiNheWRWXZUQvsHrw5F2REY
QKL6N/UmSiPye3XD3TBg7SLKx2BUqnaDKbVrvbicfmzcJGp1vGU+gHfrF6JnOih6
wvjQqQrNhT8V+f32TipiZXaO5zAaAxCG/oxtbyndYIyETrcPoR+L5K18CEcxzsWw
4VMuRmpw26o5K8A96xdnIF8ZJzBUfTAq+rgmC6jHUABvzkBH2gsyr12lYpt6XPCj
V/vJESa8mrCx6u+j4NmP3aYKuRgl0w8kcRnIT3M604K6A2z4D1pcJPPzkh/9haMH
g889jWC3Q57KeDewKF+3mqE8nkPQwUKER8TFx19HFcGNUzfc1xCfzrWoxdK2LUWf
6UYfYcDMCnnklX29MLeXSz3xaKHZylcqxSY4MTMtCFR5KNLjZILjU3LA6slY6G+z
Uw4BELX5j973c9Wpmu3y9OWRCw+ZNyuxS+sPlRA5/VxR4uHDuPbs3yPEmOUafrJI
TkqT/+xfG4/xj9AuPbadsN+bENORjsthH5Xez4XEv8X/cYCXCObkAoYQ5PClQnmE
fjhXc590x8CmFXAZdWMao+YbKQ2zuM8LzwrO9BPR3v4ZI3bcu777jvF0id97eQvc
bwj0JIDJ6jaraEQuAhXkXJCsIBoF6RcApsv6n6Ntn7122fA37d6m0BVoGuPPoH+n
xeAE7PWqboF5vvkRwM7Lydm7iAtxTAMEyxaOzH8zbfaMzOtqZ/oTfn38mQu5mqOX
IMON6Cl6avJBxE9lEtVtDxey7Qc/Mmc1hwc25IUxkS8/zEPPP0vBwBFhrtdMCW+f
NwpUR4317FkGYtE55I5ep9Hp0Q6t00Nee+qMZG+GvmIy3n371dp7BbRTmuTKNgqU
yEyvBWrfAc7/ALkMz83LKy08AeET0RDFH6ewJb9pGcRMcOXPZzw7RHYb93pOjuuz
oRv/LR5kKA/tiBC08iBPK0N/k+Y38aTZLrG63TdoMZjeQKa6Fh6DUFNfb3OwX0m3
1bIEp3xYvCoDtdWroyAvX6XGZeK+cSqe+ddkOnECSKXoFe+7HRQpqPsdDAsgyE9p
JppyADdHzfHQ2OGBFWeKIKKOXBbgp69YoWLZP3LxHRTESBSDhZgMs8URB+cLW8CL
ZLXAoaXuUKYI6TGBGHMsbmTS1mWVtEy3j/uHPLzwpUXF4XX5D7X7YbAIOwPZ51wE
oM2xU2GNSCeznvfeyaNgrDoz70FsXcVEoLR5wsOozBXs/RukpFBbR/Uo784YIJSr
Ei9v3qtbHx/FbOgcZbJLgzWi7bvpIue9drTjDFKOQ41xrqtyooh7YMMaBCO4LiiP
Fxy8yj3X+Qb4dvH9d4pH6UxlHGtYak6Q6DlzkA4S93YbwB7n8MK7ZX+xxIO2ovCq
6vylsAx7KSiApSs4ZqlgHq2580SBYTA78KZuDzikVA9Vn4B2syo1iZ55DaFX7w+L
7ECFFB1YVk5HBPTEXjEnFohOfj9U32PZf8+qIK1A9+XT65DIaaj3uUI/nko3DXK8
6VxGZl17ML+/ATB8sgs+T8dwG9Z5Br3h8MF9ulpVcTwPfCwCPPn+e56pQ/0Axo6o
ohl+p3Ot2toIRz5+8kW+3km9pBJlRJMJnHgo0Dw6Awp5iZ8FefB/2PLoRav0llGr
6scCJEP6C413q6sexRL0GcOIMeAt6NNJjEIfQcqiVT7vMrhv9cFQs7xgxVJCormu
i/7mzJUMMFH6Q+iJv1teduTBqyTr+L1qoQc6qlPxPpW6F9xkYGko+TMoNOeNGS9n
ktG1ABWWes4c3QexsWacZMXgznwNZvNVx0K7pXmlMSd9Acl7FZoYLcmSPBsNDgcP
Z/4YqtcCja+nEaFa6wGnehlKsEEZPoNK/Q0UJmrvhpfeZKUiB0+geR42TcizFRoO
2d63CRysuSfK9iABVWcOfMfzWOl7uwyrWRm/9+TjyCX7wE0gvCrZFJbSCBmoGFC0
9Rgioh1psmatF5zxD5+2Vq9er2zHdxH9HfItPx1KuOg9XCynZRzrquTR+0XTMGdo
KzqGJBn8zwptfkpnzOfJlnKx+s1S3qoUJGucVMY9Ri6MEfUVxeApWKaN5PAQa7aS
xWJCho5iVJBOO5F2zWvIM3lfdxfV+ANPzjh2dV2aycYVotcq4DLbxYLw4EDWjLeZ
U2Cs7saEOrULKvpphl8dewsnI5yXPwYzAGdQ8AS/XO8X3dWgXBfAEU6fObwFCl/u
kO0ajaokJOMPJv4rkxQppxqEDUfEEuAGTY11i0+vGf0Bnuy6zb+bDc/5WS+/BTt0
Xfsf6+9vUKUKUArXeHTuAbpMmIbbwiBhRMWqliiSWeZ9uRDt8qRBvfsewFsgFDlO
dW7EphFf8/jyblOccZjuYCZg8bP9UQCIp6Wocr02bOA28xwHeCcfSzFJ4R1rdmwN
QBED7Qhhzz6kFBI0GbYDDWmXD5qk2Lu2qn2HYnQqzehSZf6sAp7NBOykQCsJZUoy
xs6w34UliNI0f/hfQPQjc6CdFujIvWaJWWmfg49ObnT4euXprk2Fsnb1ajKlKb2q
9QsZk2VMQruJVE6PWVqFeitHhE6WNLCJVaVp8SCiPDX4Fz9lC3+8n5TOuBty9yeq
dwDZbRDElXenpGrI6ERMx204dzsXVHf10aRZjgARlVHEWrR8h5JDTIw30mEvl1I9
ydJpa3Bfs2aitQmQJmG2QYgfVIGeMxKzTVlR0Zns5s7qlGa5vfUUlpftSY54eZ2G
e9dmlv5+/ITSk53qVF2dDNztcuy7u8i4J3EP0WQTokZgKpf0iBXXkEnYLAx89xd3
dG/VrcDKJrKN1UnS9OmkLNY21E/bpUhk9gcxk/0qhB+yhXe7dGSg/XdqfdU4qC9k
WERc9PCqyzkzFucLJ4iA9FK+euH5KccBskWAXKvhqJ3Kf1nM+j+ncg0zjUSDLB4A
LaFc+Bfjm3isSKaFR6X7r2J6g9U3QtHmhN4QvaMYtn/YBFQuJx4wjA8BQRb5cdoa
dYoDACMiutjysZixP/QoKo3Yud3ApzzHXML+kXbAFF3sgrPVEMl1pkOnssq1ZTRq
8q+7PP0wcMnYuKmDZ6A1T7p8xgGoIazxEDTvo3d89fZIa0zxefelX74IW7XxFTbY
BLY+2k2rupMSKFfABQFcBklTO5UVO37JFZkmP1x/chh+v4ux1MflsTIObeN6EIxD
v68SUNCBDHrle1BTIzpHUCP5aysimND+/zfQf13pudgJVahNi+ojPxr5W7+FL7iM
xvmBVCV1s8S2ohJTVd3BCZfsS5A1VCNJCntMFIYofXi//C4/d1DQMyWQpI4aMIyy
16wWZiL9zvQu/OrinT7y3nGJUefNQAkQQkydD83vWU5xSrWghzZ/ljxCy0q71cuz
oPuP6zrOx6IlTQhfdMGpFwKqS1F8Ey/EIz1R7zFpVEw+x9320BhsmPPeM8amhJwc
NlVW7pL2SDhHm/LqoqIiP919yIGgqr5JBh1Z+RI7xSgEnqCTQqHo75etHtfSIfXq
dKBqbHr3kzvGsK991mmjhZm0vVMrUbBdGzExLfNvEpEaj5uDrie5z9rliHU7W6LX
iY24vCT+GPrmrYuqs/eeUvkfE46hnOJcKk0CRpbNFaCQyjEYKj24CsxVpUGL+5zq
Mu4EPLvKSUqM+GEiDTlSSJqd7+DOL2S4D4/Hh8GVsSr1YtE/HBGHU9dcckPmhRyF
qcZYWmzYDD6lUmb/fFW5JA+ixziOREZZ56aGc8+HSNwGjNnTjoGKOMzFs5YSyoBR
qBfH8OCPip6SULkr3d3XER2U99fOZrgSn/SZ0z+GuhsxuaFUQBUhmAmwqwahM6Rw
kmPQSPps7brtCuOGamOo82gHHEHntHJ5YwTHhR17q37aQ6R8b77lkvHgIF0MfKt4
AlTJxWIXhYHFh5yEaaHf4fDhR34glaRq4JxPtNm0fCUqRBNIcJgDGAfVhYDNzdNA
3bVp0o0BU84Kf7UyEOe67VCdYUl4aY2tHKSotmVHyAsIKtX+byKDDgwGnQ/DpJqe
BlIBXby1utDGgA+upxKlClkqmCPrvHZvyuhfIdkiGTYrs33sk98q3GsCWz9TdAch
bN3oltTPSIiqBsDSw8JwK5LHO92PSFsyuOChOg2f7pNLayDsEW4l4umSLRld9FQE
V24yFaFkFa0G6t65bqYMFpUPHcK8ETc2m8KIs8Rh/nSZtuvVaxAP5pkSpBi8c1/P
GIcXLKynLXTvwMa/OXlp4sP8p7+oPDBagthuZFobNvH+u0L9ZXGjGOPhhNMOzJ7I
yIi1ka62osR4xQbtYWfqWWZLTKdHiQOlJbQUc63NaPwwZ9Y/lBA8I3WxrE8K8DEa
mwucgBQ+NCsO4R/lkyV0Nt1rYXZ4L6d15RYW+r68STaSkb7lPPT0ihTI8hydoLks
eno57gu5v9T1FFd0OGt3T3ugpn5NoxwXeX0MUK/WJrjDftNF9t54kd3uF6QuADn4
XHGABPAmhtvhurW3PPpRJ/QxjI52tx/Et9QJ8FpQ/PvQT4zhYO0AF+5P/rFJf6vu
KjlZ/WJ1g8fQJC8+plYBJ8byfhSmTDOLQGuB9sYx9qdbzAQlx4IevfH/DEjhHdsP
YoAUc5e+HHan18n5YkZlITsNEFYRyEy/pM9lp0G9LQ3BuE9YHyuu/0gYeSTx4m5C
L0MS5+UUSl7S1bkzeowbG2qO1xWCdPBSTrHRNKo5+LW/dpuDTI92M4YspKL+a5fH
UKzPR284r2Nqwki3RJ4NV/kUSoVXR7GOwDjygMinOD3S6KwR+hUkhe46zZMmn1Y3
oQL6N5MV36IYOSELczbOKGecRG4HYp1Y2PsFr9pxyh4Y7Xg9M9KFpcj3JdCSjAZX
rKKkHeHnnzBIGPaeFrTTwj3poBoU8GN8joI3wWmy3PniPIuK4Lr0ZTJl+x5FSj34
F4ilkXvVglMqr+8LukSuVz/N8rvJnCMyqlJjkl1iAm52y+XZQ/dmdwCvNuJO31kZ
m1U99wGdsZ8ce4NKTjWeARn8E00eo5es+Vidd5fnJbpPM4Mrfi/UGpY8RAQPGCOz
k7mt4Lfd5A2RvbB9cAYP/qIUzU5c88X3xOAmgve0G9JXZc42ZFeTRRSTQOzN2eVw
yMbrxXd5Lu1FywB5ucLOuF/Qt+mXTZa5ypGZiWKLi/elpRQ5i2YjB7G/oU4Ql/j6
XiidAp3dj8TqAfvEaJXF2ipkzjrav6fXT4CIh+1fuU0Hd0/L8R1C8Ud7Tra4/dkJ
2QtRWTptaHYcsqfHtR+KU1n6CwW5AiN51Z+0+/VNBGCsbR4ywBq0gnCdyGXk6+JJ
SvJ0cjpaBKSpTQbl3D0bVpKysPa24tYwSIyszX6JEBL1eI3J6EBJm28EzIp3mrnZ
D9ACXWTuOY3YxR4SVB0HJ+fiftmpaVHZnkMYxGKjeYRo7i+TK/l3OQCfa18HFfUk
10tei9A3wMPD26JZMhc3Bo8MHLg6Zxbuo1jdm6avNf+IL+EPi9L9pyH8WgskzOjl
/QYkaXE8hH9Rf0jSxwD4xLTp7BelWF8LFIXyq18JbgZga2rUaQFriOWr29jAMtSf
z+4nCwCt5nT06sEoHURXenFvwDeJt3BN0uSLG2Q48yk45gZ9lA4FIlKPoLzZ45U3
gDfMODVBGMY2ehF0oaxkR91a5zAMiagBSLmSmqb+eQD/YLSHyThe98MA1SXLJjkd
0e+jJkm0rha/ICLGN7iRDyZwqrecl1A6NMwfag7ulEC2XTSvw7R4veUs4MCIuM2f
raFBGkwGZ+j6dbhNyYk0YilblGxL1EGSSUoh92UkERPCd7czsuljke7K2kEsfSJF
IyIA/H+7wOmAK5PVrKybDqZPpvjia6a/evNfPW7y0sUDyEcT1ejSQ8/gJumeXe28
kiV88VktivsAxRnBJXDYGbQ67fJVt1T4may9rY060I/T6wzrBnkdxCKGbvQH8pRn
9e/l6b1yZsLD09KlCLGxoJdkqkVGH1PIsFzULOF3xMqOmpolknwAMNPV3uHnTool
ZrSqNSu8uMcpg8TigRf8Mqu/d9uibttxpFOJ927/j2HHX3731peQ1wlvgp0Mo4VN
e0cpPpdDSQNQMVWiBBkeahcs9ldYHaEWgYx7sKXyheLjycvHvn7P+zbN1eaPaTkT
Z75rf3aBXwe2FnlSyA1g+IE9kVKBdRTiqCYcfaLREWpMZ8jdEMVn1JWkyC3KUlKc
6N8GQC0UbiKuG3DWsMo7s4Th9cOf7Ilur8QYkHVGxQRs1Fyxa0HhmSD9Gi0mMqy7
tzAzAZtmkqlIuLs8lxw2m9OX6FhQotsFbz+avX1OjTL9U9X7Icsx6Q+fJI3AoHPA
ggHKiBlf3ZVMm9cB9jk5y01ADBDZXkBDaFhVT9mIb7bdItr1HDobGFr7nLU9Cylo
gorWT3IiYz6OVT00R6qxgVzeymBy+ikhrsZ9QE7lMVX1TdTirT6UQ+dOGvWQJUIv
/uSvkRxkq5qf6VZrKa505HPR1Y2r7dE3UPbaFsl68OWGred8USC6yJYPo12L5EFr
w0GM4Qx0B7XnrRCeCkPA9K5DV/fBW/osqi/uoomj6oo94HEpwXOyM5SjdovvVDof
EktiP/pT37umIAM6h6DpAel7K4VtU0+KPjP5qQbZ6X6EFWH/c04QbTLux/qwjNAJ
XQ6JHYkHygF6mOS4okZ/giES/17ArMXOqkks2zijeBXlQ5hY/twPPkMTHEgHUER8
LPqcB2qyxcYBmLfv5eZGRSzGlCieNwa3ySr+6OgUz5bnLbSytA0uXdleT4UppeD9
uNPMPkl80jOHOveABD5S+KAkti2MtV6blVDW/LCkZS3YwvFIq3THUkxPtkpSwvmq
hZFgdJ69W3rM1wj5xQqATxWBG8/mmg7uBsoztdEpm9zZpn0fKOsvDMRIrx41zntE
UShod3gXiEgurZayvsGHSWitHVwujGo5pmmEWkJCUJr0cGvuQEil9EkNz7v2jgPX
Hi/oYfk8zIRyAWVWg3sDitzaA8wAXbnv+nmnvDh7kJgbWm6dE9UdINJjJ9BZoYpr
QUhR0TcoUdfCi3Cta+a8f9PLTh1eTi3mE4e9Uk6obdc7BHpstAurvdwldl+k4poA
XnYQEwcziWba864dTFNUlKdtdfAR6mEo1GeDnk91FYOsNMHKD5TVrswUiVh8IuWf
APtIOc9uTy6qG3r7YGtz+JbhjeDxXzE2Ai2U95FyMXeGYxo+xNXZn1Fxns+7/wYR
U4FmKGGV43Q0YLURxXUtBpi5SiZj6qSZr3Q+m436NrSd7o6/sKbcGS7UpzbOQ+qH
Y57t9opfsgBhYQ7S2HRIJCXNMLkitwo3yxr9sHKkrDcWQY1xqXtuF/o3vgPSQL3c
DsK+jcmdHDy4KdDE/twWseG4/QDMjaERutNefcRErFB9rJaaXmdJB8relop3ILwg
LKHPs6fEjDcnIwHcNptk3PmzAffNmzFam94rIc7zZcQ7yex9/BSkcob2S4vP0+8o
CwlinuSuv3XfL7sK/6c19QmiRiO6SRu10j/az389yWDo9JtBRlyihh81qrFtwu/v
E1zpmrTaNkpYI0hisfqImZR5cARhGMrQU6yNx6Nf30VFCUk/ntBJtHvtfFKXNq0B
Ihg5M9wSpAeG+NCkaNn50Oaz3JNYGv5mQFG9fa7VDUUBLnHV+txtfKykn/Uw8KRo
gcYH19l05aeGyXFenxCq9Orkm4VYSXTLIJiQWv5OZ4isQPsrJMIkqE7fqlxm8/ef
3B4QRg2LFxe59B4ORPpStJOLKeSdOxl8qJNqvSngNIOWWeq88phed9AZy5qhe+Yw
xlHDxgQ2BtSKaWCbkxzgMyzuRJMFI4tti/oTdz/sDNNkXGFuc0EGrf8VPnmnwqXq
X4EBJQb6XNRmzDRBn7lA4BtkaGkyRs/u4+Ct/wO08SHIgounULy7liZy4rD8V8IE
KpDNhCdbGKwpIwm9VKiBq7+IeQRyCJXC2OnnouEqPzkI74IzVB3XEu8USZVUmm9V
fjlwvjl+G3VowXrw9w/5y4yG6l2lUyureL28OLoAbkSuFoq4CfD6JAdV6Rk062un
1XzIlMOdJD8OE8aV6HJPczrYemb1RYwwbWxEyPGlDTyvXc9BrD3QwWYsp65YGfow
hcbIS4YcDNDrgt69+aBI6vfMfhNjgmyA6UhTFkB1Ng1jLYY1rzJwDkB/1jyAI4Aa
KIltvgLRpGTYUty+ylpTDULjRqIAzbE6KXERBRh9IBsQIYMQ3L5dybqt0VRU5Rgu
RsCqGMX354VUyxBeuUoV1I4T2iZaPRzNEI4Ag/B6ZAvzHI7HHtUMxbiY7GNYl4fc
SLoyaaMzLpxF3z8hhuNJWdHwvEdHHmVh4Kz318b+q4sJOw2iH/vBNWWIsYeE8Ibb
tfqQ0dHJzIf9xuNVQUK+KBIUgGpe/0PQ6oY3QV7eWVBIz4EYvPxAqc86wYJFWs5r
14dowocexGpXPZkqrBKb7BKAEYkx1C2F57j4DlRB55zMURNMO+blxGW8raOli+mV
gdph6PoONi8gse1swLguA/yfNP5B49oZJbg1rNjeH68+hjkvDYnfDnjq/+E09hB0
xufNwoq86Hd0tRuVzLMRixl2L7D7zp7k4zXEDOLMk3qsBN1fNe6txSJQ9lZB1UKQ
ih/+voqi02+nBlOCfn/YQ6jhJnJCMepAuP2673JQznDPUGHOCYcS7JgJPIWikwa8
GgISHtlzfEJeEC+0Q2jQGS4bHB+5qU5UEf9BhnpvlvGPV8UT0sHJ6ZIgcTvrFrW8
3iKk88OZKvAOlXxvGt9hcKj4uduzjymvrngG50U1CWTeevppDeuOfyRl4sYpotOr
lBk3fjy0GOkfIK2FoXBN7aVNt30ua+6EnYCO3zxrd16kbkZBvb3yJsRyhOZK1b/z
Bt5/SPwJ1ocuHhWJClOuG4Ih7l553CVtQj2Xfe+js5GL5Uam268N5cDgzxDHaPwz
E76IhDsscU+zOaRt380WGtp5rxXa0tNrpDVFZA8EWco5Tdxi2ltgWcMzB7j/ILsP
jCgA1KRzGg0p7BnY7SkmSV6ozDpCYF3MPmDnd8iv20gX/URogkfv6JwcsALxi0w7
c43E66MglzxvXJBmJnOhxR9J2QvdYZnext/zIngaGpoEtL6P68ZNfeC2QShFSRJ2
+IKzsmXeXTGlxsT7SKpxt7TbI4EH+Fmkra92XG6jnjtHvXQLQG/IDlQjfB1f24OR
LzpXd2M4DvVzQDYyTu82kxntIHbb4plpoggNYv6kraIyGvXxHSA0/Xe8PQJ96dof
VCOsKciSIcYPzXECljDw3bLVlAwjz1vR3HO2W2Ao8iXl+8JEiIdgPGkpw8t7PcAG
DK6zyini3yyNzQ3TSabgCngFtZNP2rTAvveMuA3kiJTv44qOtaYJMlBgflGKp69B
o6HONxgCmTaPtD89itgFd9t+sez5SLIiF87jDvz3UDpxjs9jT+5n/qdTqz59iirB
YhWIkp7ECKC5EoHLBdmKFExMaGr1Lm1ndbPunbneeqEQHepzDS/mPWxB0Dky8x7S
1eATQ5JiQAAUF3mXvLRiOt2LAtAvpU+rJc23chtjHUk9HqlINi/VhMpftov3vFEl
Oi++a47sZA7FFJY7vtdTdQgsPFI+Mgdcu82hzIidA9Mjhq5mB2SA8s/aGlzZmMTV
wi1OXeHwLARhQxcrGymOJXUkT4ebpN/GKzvKii9XJ1a5RPFFW8aiYyHsVSExo82b
iLEMK6W/6t0OB4Blp82EINFX8kBM+iOV2HLomMODvEuNB4Gj0QpFiELf+jkUZiSf
3Egcxsf5Yn7OG6Z9pUa5cLrFgyBIAfCNP/cr1DKJJrQsQmvdwcxcIQokkm9mcQvI
6pglHwKTKZJOsZt8aGMGaUb0onPxndF7hMmwwKjn+NXQE9wtlIqqrnZvPIREwkVd
HxDkCoLUhE/Mnw2Crmfdy7as13ZvhP93TCeXAczc9OyqtvwrRaD9Pyn8Qh22RF/H
SgpLniUhk7dPKNnPTRajaqj/nVDsvGrCEom+53Lww12I7MW4B2MKRS/1UqwnYkOT
B/DogVGJ+RKPdgRLZoWr5lWI2O3176PT8dlATmv090PG8djAxOMq2yOUPLsRis2r
19/STkzFGBHBc0W/FE/bKr7e4r9bTpv5bnJHWFbaifY7tYw7Cx4QYw5/OVxIRJ/K
w81laoLa/RsaREgFhTo0BxSZN22X/xs/WEtXGtx3PSKuimzcJdjFH0GG2+AVc+2d
YFPgVF+PvJk/TSIr5vTr1hoegajI25uNr6kjAAWIr3K+Bnq8RAHJQqNEYseIXri0
kDQsahlyGuNb606PAcMs2oW8e61ql93OXBeP4N4MnE0SGrpE4BUNYU2+s0e7lzJu
fBBImFZKdZTNh5f3oroHhPXg/+c7dyTMSrSeHGOcO/Yq0cYO9VWxY8xoYSzW4n1f
xMEA0LT/Y7LzJwnIWVFNpb0KYvUurFgELNDX6JEUaTz53gCTgZkkZ9B4QlidOT0/
C7szoWOpEJZGjzEPNAYkEk/z8Oo9bXMYu2iPaY9xoA95Onas7vUES1LlEmYs/ztJ
Mcd9DXJFSBsjmA7r1XaMNUDThn8iFcm/iV/wYoPc309/nhPlDtSow+DY/xLtDUJD
JkLOngiehe+jkxS/Kq/J2qlwfwIzxuI5aWToZ1HZeg1MfkKc1YCCqi+VKwFsgBRU
UdPfB9hJdIyV5q9cFJkgSqhTj7XPax5zrd2O6VjKEpsa/M8txrbhWm5OhAg7Xozn
wHlsCoVuKinQHeRzvFGIg+ccVYpcGu0rEPUMgc284QYMcC3rM09q20/4x30vaQov
4lD7IyZX2a0rs0iJEf4p66kD8f1eIQL0HL7K6U1RtOoV1iXIH9eweudtcMwIOizB
cZGFGICULhEBHFmurVJhpOrtPksPCPWFRA4XFU09J+vD+Zwg5Hz3P50Sy2MVfMdz
MOmCux0sq02gkZVvH9LScaB+m6Ksak4U9So57jMAqLXN20sdIGgk/D1TScJ8vOvg
XMtKOQ00QfiFoStJ4A4qUyBW3iAASbpQQgQNU/eTTo2/cMYGnjCz4OxEkKSdJDCb
0Y3z59gNx4ipvcHH8Qg0O21eIl7zwQ8mpDBBlseb2t4pTlBPuG5aJA/xLLu3NFxd
+BBG6k5iR1L28Ig8n6KwWVD2MsRkccRfk9AydaNpfHgu7yXj1TBihmSAvBur3EJ9
PShd8+ZiPaBCN/HF0sQw97s76dAFwPfEnF+verWbmawu031raMoBIFS+76BlCOlg
QemYUIvoOZr1uEui40DbrC0XCEXNWWjIF45Mk866vIxApYynrH2jXsy8jlMhvD35
gIT/twlzE2dHMcq+r5e9tHK6La+/ijKuWshOjZfzEOGPH2Okk0WSTWcEcYjlGAyG
HUhuSnjhv1p5xx980dOOt3vV9ZzYLrJtVbuwB8PP/9DVeDfBEhKV3ajUdzVKFQzg
kmADJKPconbfLv+ERfYjaQ9lm2k7sGX2U5oV8tSQpDJi9Iy3w1+PITinWYBZ76wa
YhvVGvUV/Dm/J5jWXxiG3as5ldgPB+h5LZDvqVyMBdcB0TR+EMkSWaROY5j8gtKP
xagwY3gy9l3/xwD/r+bxXEPIUCtkk9D3y+yh859VyidBJsyyc9GOvRGIyIwBEsTx
uD7TYH8nDm1KTtgQWMiA7ALpPTTiLzH4Llo3bNVVaRJWKXk0mJZUK0kD7+J5PomW
G+jqJtsEB31NkPSh46ABp1ygKQ7p4WFqxYWauijbhHGZHIfIFWcmt3cEmYXduGBP
ZfaHli6OPGdUWO7M3UZTkFvBj7H9+cb5Pu//cCEcO6/duej/feYsjxeyh3iF3AJ+
W7hbby5TJRdyQLLmiDvOmtAr7EW6/OxhoHxnrZFr5hhiWCyDaXDzkd4D9b3we73o
mTtkaDw8pFijIM18/+pxf3LAEWZt3HEN+8vmOadeOEKlzI2TCBL3dkIw8MVChnTf
w5d7QyqVNdh6U6SUeZ8ckAUyeSf6gNtksOvv2jz4kASTKL0mxdgPhaqFpRvynHKS
H0OaS19XLsQjh9PGIKsrwf3epZwzXaJwLQ14CLI3LwtWlujFMwQK23dX1+cuZnJr
iqjXCu1KZpiIIDPHhkDn5dDApJVZ+pSD3T9YNhfteKPlRiKIDpWVBYF4RHdG39wf
HqW2/kcRmbtGbGkgtTOEpZ99kXm/iKHn8idYHP8CPaWnLrEW8TZJFByyvwsx1Vph
9zOg9A0bug5kx2djU8jqJcN/jEvvdJhfPo9EjBqyh9rg+pg2m/gAbAqep8idtSfu
CSq12lgfdwIruAhJcOynclXSN/vIMszSr+XG+KPUbwQ/iKtKfdS9df7LKsVI4eH7
ELIe631c5TwbHqsSFD6t67RmbPCD2FDvDpVFq9U+uTyZaUW781dstpy8NZGwyjDL
MCN802ph0EesDrXrNcsdUrMWzUZAS5NotmJ7odMV08nzcG4Nx3wNgl8ML5rL1lIw
+Y9pL5/AhBn+Fc/6X3kiSE/Q6T+DlvtfR1qSi84tUStDLhGjy8z+LLhQyhUYMmUg
q9hL2CwUReh7ge/xYX7csoWceZwxJWW+i9DIzjGBb0zd6M273wQZNenvnUugnr3F
01t1GkXJIj12kmRq62yoEzjTOFyvYMWQO4F5n4UaBHvOVy94r3tj8hy1VbgudswK
NJzUmvrySgYBHx+gkEKGiVTWxG99PXvA+h8nWEB4MxWjyvMNaNS5mQFPuwspamVa
kxRUL7xSA/VoY8jI0M2Tt6VPR2mvvq0FEFsG+Uuoo3r921Ul84qxEsBgg2gvBH7D
96cmUGsb1oeJgdu2tk1EfWoT8OKW6t2fmlmclKGogZHTOnd6xtHG6GPwnrqABtiv
4VX7opZw6NzF4LBei2G3yA51Fj1Gtbnjl5I38KFBxbSJ1FvdinOx2GD9hitSI0mF
er+IU3Me1Sjp+L8KVVtDO+Bja8oqeFlce5VZ8TR+MUcXDPctDAcIghJsiA46o9AI
NiFwILpPeswqMPc7ZLxssyd4QA4RFUBaGgdXpNbk38Dv+NfT6sKshFCiedKSerN1
B0RpiV97PJpCXfUaWJx8xDp27tepApVYvB9xmTvdlEac5swz1yi76mdezxlSg4I6
X2DufQUz/Vt6BLVtIfdHPOoMUFEECvkQbuZqFbOHHHgFyrNwe7YVBEksBzIVtpOb
DRE1K8QGV++JqVwzeatIKxw2vDBIcukoL1THa7bSMKwlpZDbBs+5gTVeD04H3xCa
2eP8OoJdm5PFVCx37Krtv0kqrdjBPqakOIMXPxRHh9mmv3ps6t+qXw57zB7OzjmW
RALBvNr2XRhb4OQm2Kb0Z+gmHncB4wPDSxC8anhEJlh76WH4lb2Y1waUAyEh5p1/
SFL8iiQiNW1LxtgnfarRvPmy4iKxd/PwA+3Rhn7GYSmqNLdsD2wKl7Xps52oJe4m
hYA/eartlXGiDJH0gmrRMQbdWTN0aImBcXk/1r0L2bJ5d+8OKaGf880G/IyiVtXE
jweUCx3ejv7w+++5gPPenVAYFu08dTNGE4hmxOUfo48kz92tcFseQbUqx2GuSzB3
Rv3s68fkMrOOkepTCfZJ5C2cd4Q5U9imvLR88aB+Y4MW7q54/OUg1/Z1qJHj9qaw
95+PQ9PFk6AtaS3lJOkpTZKBQYIQWuMTgdSzBmVVFMDasdj2HJmbfyfXpa2iy08d
JsyPGAJiDDrmULWyEpxHEZp+XMlvzKBTWbN9ZSKADi1FRfyATnDAdpNDBHD0MiqI
BqVHqHb4gagdsel+cbVXrDfy/1gfSQkYQo8byCZkxMxjRaJLxXxnk110MDA2YvYQ
UA9Y3lQ96lBJh9jCyWlOUdtge1kWTPuW/cAAk3ifo/dHBU953WTmGCOTGjcE22Ea
THeq6zHWCOEzjVfGLrySTZq9e3/CnPF1QoCfOzYAJcnVYX+J9hbtyhdt8b9a3nT5
KFSi7Dfp5A4ODESsg1Kp/nx/a2Ml5Iai9Pp23uQ5DhDrD9vbqRsv9F1bKd//BZPS
Egs95g+/mpSI6xrIbNEcJmemBqmZR0kmjE0slHF/jxflo4IQBf9zcgbt58IGfoaJ
i2uN8xk/IB2NOMwfXyn0Tin8yV5w0JrbTuYfHMQXNC1Ho/2imv9j2X2ehvLK0xs0
83tX5WrRXs3Fvv64btYLGGsQZ4lizjY8pJvVIUHuVMTcRPoefmMCBJNfKunXXpin
q3KQR/WaN/lTL4F4+vkE4xx89MqoY/hP7Nsmhb5eog2C6GM7dWS7UjhbOSy6em3Z
/TJ6HLwzoMVV3ofXJJdKZLDTKaDMv9QQcrLrScBxQ+XDFCzaVwcJab2vOG4/U7HW
jikVdV93vb4WdyLK5yyhuIKcYitNz9+MVpQDP4fHQYh37+AjDMgdr8ZkVwxfp/CR
oqEwyn5fKzxm8KMbv2Pk8qgyLAVSwwC0It2/InGM7H18zWoXf7xcIUBi+mcEqf1c
6TTHnyoa2olG/7b09GcLj2ZwaumpyiqAzavf0497gr6XT9Pzl0u4eh72MUsnIdrW
+jjo4ZT3bUlKHyLGMSCVTo5PxgB55g9WQm6b2z/BdVahTFNng2fQNGMjBFCqHRoP
0KQpS2LSNpNUD96S8+n3i0+n3XvDXDRh3/PNI0osd0xr/quH56rwSsZ+Ol+4Yh6o
96XjOy5DSQso8RXwukr9mmQIdxsg68epCaCVg1xSdLhoefftTZbcfvgUeYvMkobx
esufHT6W0LioSmdfrdJfJA5jEFK/ZuXAAEbobYFHaPXw6RsUYgFLohLhuV71lVBb
0tnV5cIFnWWnxAtkZjq95Ap99Szu/cbuse5oSvfcGs5StYhO8q1T4h3kZR9mDrDo
leZe9gSMsp51qgyYXUKmX88vPc2l5KfcCls7sBTlFMyG9/60A6wl2Fbk9rQSr8TE
o8zUVvRS8KK7VrJ8BK4LO9xS9YamR2qA4lqmz/XBjop6+2pcw4thQdsX9FX7hzIl
M4fkGNRbf8qArOoxwdfVJ6WcVX7DCj+4UK7tjYogYr8vLf3ZhvTSbFdyyTdgxJS5
ltOsv59VwpuFvelqFp0GfdDJPDjIvgE9pPGOIJMJj8/i7onzZVAVCoRXvdGzjcAX
x5dORDKTtydXswC/p6Tr65CC7lG6uLRmg716oojHmAP0BbKH/3uw7OOFGvixIZAK
czoZ7mWjI6WoHJz4skhPePPQ0QAqgxJtYroae9kgb0EFUkBbaUptkjoa+pI4PL29
OHlK1A/V8MLbHhZ9izS923JCXkm8PAVhL27N92bvjMoUH3h0FOY/3hJvFQXK86pE
Q+wStr3YipCEcn/EtrxqIIoGpFxtkwxRWszWKgnkg5xYiw8l7J+zv/4QNDvGvmXF
RdRArla/c2lUaHW7yKx03Ifi5OpLMOu11ikt5zYTK+xXo4mAQA91zCzI0d7+H0nW
PgQNNLtMW5kVUn2K+tvoGxk/PqTsw2Zz1LJO7PugolEII4I9H0YJ2yGNQvIISKq9
sxhCkLGasVwfsZVDwT+IQJmS09bc/fljZ90A3Q07bZaJq5tIXuYpCxm8XAXD3N/4
qOrIklvh6ou6basl+OU8m8oqL/pEk/fO+lQt04AyDX3/Og3ILrnkr3m4qiooV+Jo
iNgx44wjox4yqjXpdk2U73NBg2lJWoXw7UaCBCKOuQkgPWhTZ/shdqkNaW6yRfXZ
rDVlCvf/CcZ28lQdrvGFNtbFMkCe6kOnnBGqBrWWKYvfGCQPSU+evQ4ZwO09KCa2
S7jBDru9e0p5+t2vqyhJGUskf7yDI0OlzER4H9D3GEuMWenyKqRHMxZB2RNRZrBu
4yYMhTNviJO4bmkIArwX5NIGjijRsCTi1OJYC/75KhFwZHXErManC9IRt4bV/aPX
ZlKsuyDXEp3aepMOfMMlHlPT0SN5kgDzr9sskDK65gv1WQObl0egKPyGS5CP3qxt
Xy6f3zgLO74XB9vN50mHBIE2YHXq0URE1uVkv/VvbCifXBOc4/gKwluLrcwp+FBJ
rF20+loETJIVijwUg6vT4/Nmgc67sWhaJCb9DdP8gCHfF+le3vQu9GV5zBedpZbn
M0Y47FnVAl1zbF7DPzi6/1tgDWwK6vpFUlgmYbjAqf4qmwGJtJogvhsa+Oj0oM0c
Sdy0GCDenLTWvepaenlvvp8qMABL5MurDmdBUyZRRRj+Iagogo5IK28z/H2IN7et
HoxpQ58i8/6aDV9aw3x3bRXq5R+HzADuIQvOUm4y3okbrjHRkNJmigiyJp3xDbud
P8AvEcJ6PnGDOVmJgrSGP+1MUAQfnBpdHP/9n1RNex2dTtNLexGeoZ4KS4m+Mg4D
dngyzK2cs7gV4oA0wydATzLh0A0P1vGK8BWKT/KN7iIUzbb1dMMhEHPlbzit9/r7
AdKVnGZ17Pj0BowH/0QnKPhen/20F2ycOLcigOD0xgC5fzbqWNXydBqFpFRI3Hy+
3qoYhi9OqCAf58YKoZQl11B9UBmv1/pjjY6gYhQ5XVT3Ds6bc8+udOknZMwPUAu+
+r2Ks0vivgHSM2XPy4Fbmqjx1KDcBxd2XSofBuj/+TE0Q2/4aViB/T1FyKVte6Yh
cusOMz062Nob6GdqISoGZXN/37kCS/L8WD5doXNyQViVpjYoWjpEJY1WNt9F0a5o
JUuCe8YNtavEPtde2gBdsGQ9kmO3vQ1AF6ZA1rjvolLwGUdOhmed9x5dHJaAMFjU
M7oiV4n9sYGNJBX4cDeTGP0/UQotFN+tBmx7jJrCP4sYgiOVyq2xzTaMOBJMg7hG
N5wkoGstfH5Ez8raY480HUg8P847WwBIFiW21/2L2sH6mtRNxV4SbKpYyvofUo/p
BtBGcUBfX/Y7dc9xd5/fUyvK70m2Hu9badiVQdIw83s1P79ZXPEMI/fo+BNWBnUR
lhRWLELgGSZgy3FmpenhWcMHFwk1J3LbbSRZxS+Z2VQ/NtmTpiJOFBgjNSZNEmRR
lZMGSDofc6cqxpGQNcZSYaYR82zJ1T6E7kxUl6Fi6oRDJezcoArI47bQeA/cV6dl
SqjGwXm9TO+Va5knCLlXNxcuVhxtMCEqpiL7jSzwGH+JRoGvT9Qg89LDf2z2BU+x
Crtb4Oyo2jgtrim6hVTelhrnsOlIcUtBhpXvkaYvvGJsLTjWHdwzPIj89IAn/mqW
NRDnunZEWDefmQgAooo1Po7MSXQakm7OFhnuLq0+EgVcoQOVw51T/kcelp6WR9t8
Pa2wPccZC3onXMlsTMwig7oQ7FakgO/viZzTGrVhzS9BPLY9cFCDFtf9kS1XbcHe
Eoysx0Yp8Hod7qSFD7z4kfaQvX8xZDld38LuteW5hp2MbjMr7WXawc7KmdD9XEHS
p1FzUqIfW+s0ta+WEc9ZCrRR/79/qp+J8fI0ZgW4ucd08oxOSQ+nnN4RzZmRh0Eq
/6izTanl8jitf0G94N7wkvALMn/puJ/SRvCqDqo/xnP1hlDjLOeVvJOrjI09dE3Q
syJnw9uK/lceBP1unCw9uB8D7wnHsUk0iN1mOVbaNmHgRYvzGtSl5dgqTe2/Yd1N
P7rxE34JBUogH0abBL278JWSMx2y1BgDmKEAlWuypCJYWOWQO/u9oalSSlBaQ/ix
jzXY2M4htUNwJZ9nf/6pkbFMc3Qh7U1XGD8IXClJuKSkRQMrnOZ5Hs/sGRfWAI6V
GgpwMJEhhxllp1NV52YoXv4hZBQl6aB05i54O24qI583VbX0mrTFa9zYtHSLp7bu
4Sh9PCJFW3QBgImJYiVyRBCU9gop2uwN1i79pyr2/CiUDIz04az5QG4C7Ho5hkYm
vnvVVRSqSok3iHr8JPBO7sZhGBO2Ns9luQCquLZzJvhas7bYRB+VLjRQdNyxys6w
Pwfrp8Q0zf04GCRXc0yuEoCvWIguZ97XF1QLcdI5KpxSOvHLokyipuTbndijfwzu
LLmFVPV0BGV2VaMjlI0lCF75xXhm50Uk6ycupnCR95fDS54cpFvwsXe6s2HpLaRS
KtKYapjHzs5bWKYJSYYnssDhr3kewvtjtQLZd9te2P0w7r3oXOR11T63A3pzUx7d
bDeXtnKHegWifAzlVxphaxEFkOLJqw1ObGjv/NeZrwEy8OWfhplvMUwC0rInm8TQ
Ar5JkDPKEzApvBt+LgEvV0nQ6E9WBU8dlsKjkj4p+ZcTNsp79t9qvRC+E7Ymngdb
1OYMs3pPbPkZPhrIkP2laXoEIBYfM5aisVOuXZ20akmb7YFEmUujHEN22qi5Geh4
oHu97uEOcikV5vq5f+DQZEa5dHAdzyJBLowddUPeZgtlNcElV7qLgN1SKGgYneGq
6BXerXfUdpZOqYteFkZKhkm3hQLcDlSHtgp6vS/aWrTdadXuiitLpp/Z4QqPbW3D
RVx1XRTim/LOwF6wppucnL6zsFT0LRjaBYEm4bxhJJIHcjU1NLGaOj/tlx6zJF3I
BjNb55UAMpebM2NRWKFRtp43zuHr8Gs3xmCm3llEWLVO/2lLk3n4ajx/Mb+6uM0n
qEQ6Sxeq5Ikzyyz+lglWi1Rx8jvLbkVyqpA6q6NoUJL2twCBphyazdcMvys6eD8U
oLhbm65ikZWxIqsncAk/BNsuosJK1NGqYcbyMqdkFz+l/P/+o/RO4gMKMNhQy0QI
gyC0feV364zOfcN1UyjAqawTyaYzcWdEcPY6H8BST6it33SvQJ6cWd/T0V5xGV5w
UL/ZgEogoCCwAnZU8ghMo8XceRjml7YpJO69V3XSzGliXkltFtY2+3v1nkljTKAX
ki1p5C6uGbJgHbV+aQvoeT3gB7ei+quzI1x6KX6qX0sfBZsWNz62xu0kiD/n8fBT
7eop/9urYmUJIAKH6wCLNY0Fy020eHFmES7HaYDrVj6Y/ZhwPe5zunxARUc5ndEZ
fP0ukDzA//aioEjKsfnMFTis1tfrG/ebtTr09s6R1ij3Bkc4/3FHb4EM4orraOtL
sABLm4Wj2ykBgO5Wkz8oK8eyLBpaIHZWygGo2L5zAwY5y2R4mz3Zd0wa4LGW87Wb
MImyFPLhKQjJiyB2MUr735qJDTESL7m+ALEmjTEKV1Y+4QZ456okjuu38M94qdAU
vuiZzNrpQcL1d9L1OK9H3oxWEyN60JE3gUQ2ZAeW1KqXbaZeEezGKkdQNOhecbtA
So7LbYiRitz3yjwA3YKbL1eRIqoSleauag+xYKaUjXirzZXUgjIJFPGQ4GS2x91f
pWe8e7NFrMn8ynAWrWYRNIm6fpzZkWu1kusIwIAlCiG0777ZB18cKJBvtfItKO+b
jXm0GCjjrHRxkK/+qmrFojrznHZCXWaDaa8o4W5Czof1UBtLeICnkDsPllZbejC6
1gu0WnmfexdAoSKv3eSMHcdUcqAtE/S882RxOf3KWLAjD9oTXF2SKCoAxrCZ0t+m
sJoccETYdOzA2z05/zfUJ/GgmOD7daT/rRalqHGHiUbSsVT/T0CEiCBrM5wi+3Kh
j2ZWub0S1ryCwqqreGUxtHuTT/KkkKLnOm90AMFX1EaO5cY7Url9TSjqJl+vMG+k
AsV8qnaYAzU5oJjnvuch1ZnfKEmsk+9Uzundz3jfBI71zOKgGuvE158c8TXOFp3o
45BZyQBZk82SAN0VC2znL074dhGBeg6hRUPkeshMM2TktAWROmPjDsA2BphIR4J6
15DyDYei2keDIsoZP1TzBrZp9o2gf+n3gLB8MahcyMqx5pHST01tWDAdme22u7+k
tj+LxjFgEdWLficfk0gbkHmnFfoeO1QQS1P2UiMrgOyP+w/ZekT04LGDDjyvyMI0
QFxammT6ft4Q0ye9C6JNBktaX0vlO0zeaZPLeHfaXi3V0hCoLYEJTp2ITCiYTXQk
oUjrZhTIKbyf1ONjq8JbqLB8JQB/8e5JvQSF3QfHee1oWk+IgDzz7yrkeZXJExTa
7HrOw9+fc81MyhCXyAd9EHDsWWiNQ9NjThwX9JVxFGw69wmLRmWXuGdRD6T0bomA
kTP2trm43eTjYYurYQzt2LqxdDSMD9SaDj+hcGEnRdPZD55dn+BKcC7cUL2Nvq0x
hrZaVJz5y6TxF0jmYqEofHk8DI+G7T/qWh0001OSbIA7nfjj0crCB+uvsSBw0pUJ
pst5qmbLGBcr0FV6UtuUtbsylL0A9Umy6zPBIp2ZObtnnNq13Mxw/GGMvduX4GOu
wq1pgQ5xwZsbiFEcGMjirbljuRZKMGvUp4DHf2GWbnqXwL1ZYD+w8WweRkPe+62k
N53bU/OUpXC51UCK9HIevf0XgjoHynZ1nXFoCWa6NmMfv5xeSXddlqW7m+TeQjB0
+GxBb3U7ISs+u9armbgUB/fd6hJIq5dMCB/BACGg2T8Yzvtoo+mnkoWF04SiYgFF
zWa5bcv/nZ29PFhGj4BTlmInGF/zrr3pN3jemPNaZ2iKxOFNjyLxgpfqHLVNAaYC
SJVSx7lvdfBkOhNDYKVIbI2Ho10dSKnu7v1/g04KF499OWjQZDRwVgvfZ9T2EfUN
ONdDNwjn80aDqphgYUCL1TI+FedGWgN1ngDopLQRavM9sCg/8w36kRCm66j3RlC3
rVMNIbJHOEOZEN9AE42XV+XAdxQbPpL1eX8MoM6QK3jo8sKR+y5Wh2MXt8l9yFGc
hexcLb0aPSrfTf3LSnFGmY2ces+Is4DfgF3gCgOCSih3w3+rKc56Aqt1HR+qGDEP
3ZKE5lWhOfE8nF4hEwC/dsLpg42wLgEEfwhy30jtflzY1yG1WCsV9Yw87WQD5qXS
pbZchQlZjpkdYQnLPdEf24HE9ddsxRnmCpo8jXFqJnLwayfE86o3Er+p7vY6zreq
p6tmFXL/AfSc4ZHkywez0NPGn27ZW9pwlc9SM3XPgcTMqqqTFPR7M6VCVm5to+uF
2gA+3J0JxJtb7JUhdpbXRuQ07vhZNRNy+UBbd00+ru0traD8pvwDeJG1CWwHM912
2pXjaTqbHLYBG4PTqZaRjDVg6qoVL/KBipLWW9Z89M05+K1wjNuUVo6nkhOkvm5+
INjMT9wGMvczqHYZm84CtXkI58hO0AFGsIs3TnQsu9iWDXa34zynlCb4XPzh07EM
ZoOpbcaA31xtIY2M64NEjlxBW6IdVTYptw/OhTMJQ5WwmdHtHSHv0zowq09TBO70
PlFervpLOlFPFauSqCvnnifG84axq4J8P28qEZ1S+izRyQcW0Ww2p/rA0otvd/1I
x+C+8BhN2y7tzQ+IHTMjjRDG5uy0d/q9bJ+3zE8ByKWXtuRlg6AshLBJfKar7tjr
mS8dYTL2qmyThhpMk9aD0E2Q8gl9LeMcTWvUavSwHAQskD7tskrVeKf6ZvieE3ML
+snwcLpg8RBVjNdjGPVfLWKKeWJStvym6QRd/D3kNuFEkBQc+1Gi9L0S4mUBD1q7
6I5b+6zoZgXiMaQyA2/D8O5xC6yEwHTzJezArxB6QPE0BoOF0kWfmJckqo/5DE5Y
4+dsSItH46JuDLdKGULJ5L3fcJLTW9PzFHim9QxX4RVxIiTbXbXHxw8UqGhDjCls
dfYib7sC9U1G2Ip5083gI2BaGZUpPDwE8fK+hEfUc/eXAs1Tk8LD/+jIppd7U1Et
huu+OB3qkIWIRIa9ugtSCdlmdvG3zDx9pG2ElvXECev7JipAmERKoXO4xULGDKNQ
FEtbRmNiGJERXfa4eYm9U8EdYGtq74Th3iTuLNMKeA9VfdhCgG9QY5ZjURNi89N7
ELuXEBKC5fR23g+knfFphteb8YbEmOnCIxXi4lLuf5b6g3bQdg77FufEgM3L7bJF
tHFqjMBuKdu7shFE2knCD0pM1iMlkv2RMGWjwtejonQ8juV6jITk6qRSxQE+SUj9
76g+r7w8aPWmTA3ZBYhnuCUUjkJrz2rAoY2QF0/iYmDbJYTSCzdKCRMop8Cb+pGM
RLMGQY8YuLGyHTALDTkcVthkSlrWfEmo5MceZAYH29Wj7EVX/ZLlp9Ah6vu+RnJh
MLIrm2UXtP4/NyVYr4FmVyFq7yB91TGlcnLfLrjFT0gjNvfwkubKU+1MIwGA5sLm
wkg+2LBYSfAgeSZ2rC0dss8HF76yWNDfMvtjmbmffau4AxplgChl0L9Sug8zDF2+
B0jffuAAeiMVWxsa7+722kSp3F/Foan9YwROuPhSfYUCbI5U3Tnhgkl9G4nqQl6/
Vie/GOCBpVJFlHIXYmIHAHuk6S8EGJzmEoUG/6iAvNMg9n5UN+yn5AXJNoec67Ps
Q8dPUrlgkaHFn6mAhgF9ZhjUSfBrSiPCaYMQd2cmo/pOQmiuM2RLaq67H+/IsVmO
VwXAKUGujiUybgKj4szUac1PnYEObgKyy+PYuE6P+NQQSxa3jQ+yCxJoQRm2POae
OLVxIFcn7YM1oi27LgGsnQ+yVS9+4TSFQZo4gRIcwIZC+mU4xSJbcSa9nmYaVDT5
3eMGGvX2rE+AHYJLZry1L9/cEPhHC+K2lZwUHvU1LQmIaYZZL6Hm8ZG053FS/ZaS
zaePeAmic6yWY+DI9JvbJoeFNTqY0Vfd5WhbJEvFbGGIPTxntBckaKjRCVc2lHEM
J/Tn5yIPUV6t0+7spy3fAYD6NnsyHVggxBCx4cRkW0PSp4w6tbFSKyocfssfn6pG
QhNLa9IBGOaTMwxF5Ia9+8ZmNOBAf4jCjgUntWzz39br1B35NK9Yth1vCUb8rt/o
0HS2/sPKHMumNsle4ZEj8rb+pOB+wUcPwADfoRVsqSPFzzP+qsCVzhV/Xy9nE5Jv
dLLaaeKZSqtzBZmexdmJ1tfKLlMkS79mqUV6t8hfRbhg4SS2XJupEl5pPjeQwGpn
ll4GBxwZ9x+1THWA2z36EjX5EeLXUGLRH1mu770WBO8nBvjcEgi5lNRcu5VWbUZh
XrRNS/0XT6nRs+a8OLs4/AYRHWMiS5KazjLv/SMMLs5mfaJFc7LDwt09Yd+0FjEU
ItewSvEcZ6zfQSjNZCPWFo6PtwytU/uI871STuHawrIrdfPoi9RTsMuudqgN6hZH
abmYSh3FvN1aBmWbsIYZp7Ycf6YJs5uyvg7v473vM238NB4DskNc1sFAc1lu/S7Y
X+QUkV0UiyBtQh5P3Ke1D4UWijxs1siPuHqocPE+tJ6pqOOdCS+Rt/+ykRxd+VH0
ZKZ/YI6yIs3ita2RSvbQCcnFvpDoMWgRp1yOuQY87vonIesH4F0yrmEsenvEAedg
vBjiS3PMSXbznyoTS6S/Z51Q/zB+sR4c4UAYM+uoIBliJUCNwPShg6CYDUYziVil
Z/AdaJGREBL0k4UW0/IC9I+bilaN/noTgSi0OBF9rQJjvON9oW2wsKsppYm0CeYa
Pcw1qX1WUaUZLjTyt8scYcHq7GuTKMwDUEnslq5Xbrqs7L+LUu6F1R2E6D4jZPnU
7BmZDZyflPwMA85/1QwtvKgRWpAoqghlNHAKyfzrVAu3kXTmBlCvtVCflqBzR8EQ
GBICMe+FPmH3UVDgLJMPSLY/WsYMyTgBnhFjaA4O6ZXUnBtKgPH1JDfmutY7LIPv
Q4hE1hZnMLX2MILXsY37GlfQz93pV1rjtUMfsFAdndy5kOrldXkiWkJ8on1jSoeF
oJYLcMbmJer8Ovx/CRdIFApt+vmRvGdrc93V8pudwH8BWFz6ceFI1JZGLtFeOJCE
q79sVfutVXT09wcvdRE7M2HkDliVptuH+h2LPTPxvyZ76GnOGze6H0RkoMSWO9IC
G0bzEWPuH9BweeYhhzXpBYaWtQz0bCgZB6Fb5HgP37tH3l1GHjS3FpbZzv70tkUL
ARVo4y2+bJOq3NlPdX+bux6TOMx2f4TK+WJ694Lj8D+R/ceB4RQHhsMQeI0SUbm3
C34Hx/w2tYuCYujgjumXWlcrrgwsfPO8KAxgCSpxNwdISy5dbY8NHTdb3yvzrhZg
Yv73vtI4b/Q6z9aSacXcDeu9Whscq11w4yjmi3YtMHakAXIQvVTaBncyr3AJI0ub
METiwbnlMsgMPYLLsNwbN153ImmAfMr2OAbLa9IWnfcE9BnSVmAmKofClMJD+JMf
MGlvzle2jbskyq7FQKZuGm/375DTlXX3aLTJGRFOowbqlWF40FpmVrsAbvtQ7DvQ
hHxpEKJwzeJCOghDwOxPri3J3lKlflzeJAACZwqeHJjUYkKHr+wTsfF4Cp1xl4st
J+n9f66J1sK1C4WFhX1Ljq+ZOfBnAS7t39sjikcQ5/i8NJYNUWcJOGB6KQYagP61
ZB7bYM7AblqwKyU6oWyNIMUdf7+BuSUP39dO5rYhGjz2qi1UhwA4WW5Cbk5Hs7bG
jKjvJMdxeu4zzqrMGCBdRIYfuZeVnCOb0V4k+xQ4D7tnVZh0rNM7V817ggqvnJyo
sP8+8kjgjIcmkKM7qx7fmQr+kOXdCDbx98Cq/aFHhbohfJwg9BR6JO7JwVYBvAG0
9iUle1+9KiH8pAeswyT3cc4D8BLGDXlADWyzIW4bO2hQlVoy3EXxvY6eVgloKQxV
UyEUKCTqrohvNa3gJ7wLD4dWmWeHzgXgE4vAfJ+VyVt8SC9xZVABI9XAG6YHkH4Y
VOUoOy26va02XemcrkCHh9OnG5YQWM7g+ECPM2x1cnmdpnK2/M9TGbMhGWhP0rDS
O+km9OJOKvt57IhtRRM2VuV57YSDMb6BF0/OgVjvKxgRue9SArIPdvcpaXAE9E6q
WuuQjaIJGuRKW9RAoobeDY7tgFzVmsgl4mN5Zz27736lTxsEzdRH/JezFy4gF1pm
joblh2IoUori3ashfgYcR2IzmophJz9QOrrPFUQgVmcIyPZdK5ZbElHgLUz7skim
r8NcnMjKbVB7ViwFyucLi3ZCaCDXh/9y6EeJOxrNdw26xDNJfig1wqZZ0qouXqIq
ykAjO8V1MG6yYJJ/+83aab5yFJzesiLaNRygRyGgJ7GUgGSkP1C+5GNMbHBHAKGO
Ui6gxSV3YHAT0MaBDfX8QHBBFQ6jCAOeHkzfAtN4F5V/LgnQj3faPj6FUkHC8g3d
+uFRW6glvFOJ5+QEyWrhMGcsFq5iZWuP2Ec4S9nNASroLLwhjVjlcEewDQgaolNI
SdsYPd3wAJ1csH7WBnEO1SdyjQB3B25dgC9G5qu9egl0fKb4eQvbB9pQ+a1iQQvB
TSI0h1LF1aewbSvoQuFoZqWfRXtRGSQtneXdLW6O16308ygl5fb4+assIQYI6XO4
wQlHG6oVcRl8FIuzNtCdHqV4nSgjqgyOlh2YNxp6XriklBBMtmEMnFo6PVp3zw4P
qkTtj7Ebf6GQ0uL8Esm+Cf8AsposHnqBe7i0L1MNtmMxtHF0zlZ67uiR4dkOpk31
ShOB5PVlolFmt/Uid68FVXcgydp3HZEw7T8N7cKRsoaIbByEYSrRKd0QYohyflQr
m+kICh9ZedMxJ41X4pQ0FCAMyQU3OQmIuZOEN8Ur3+ERdvPqIAM1WLZ+CMSP7CJJ
NKfRbrffFPbdP9rHLkRu40HNRECXMEBB5EaQRfNAWmuJLlQfTwEwc/0GL7k3r3EP
/5PtgZscEL94Xj+8mSmTcdW6RiVEteDZsi4npjFP7BUC+fCgAvQ6FOnW+fvtlquR
xJ6FDRp85YTXx6xSgLWZIiNWWJVNQlIzrqsLXKn3/7hdhqlDZ40am3cvhfq+kqD2
SLCX2C8hlSR9ERaTleAjSEa0mSOKK1uTcd6uQTeI0fij8JhrkMrM/PcbkKlQKstD
cR9F+3NzUj1wMEqesKZlK5kaBzYo6sMu6JVA0/1jD4bjc+X06QlyLGUnbUKuIFil
PSjfhhn604vy84KDoDy4oppC2GehE3l+j68M+gtDod5b78Uk3t2Gvt8uLTlaUc0P
iukXRmC45g8Lwg+8ujDJUZyaEEAkWVgYXuiLHUwawV5w/2yWBbnwactvYagEAyUQ
B38A4z5Q7S8OWrAilN4QaBsMSSBSVB4um5bLXasydSsOQ7DEQ3kHJa70WCKqExPi
w7OVn5SAX302YntM8Umpl6twyjHwXVmmP8ZQ8eEAdeXptn6QUz/oVfPNJimYTxGR
8Vfp5fnuisdpwZsK0Y2YwuIDL2NOqvSVVC40WL604FBNWrW6FNtnvNSKQxanhgSh
700IbgiggBok4/CMwIubqs0cvzPo02D9WlA6rWA00QpKnZ79k6pE7C5qXJC/fmxC
pQOaWZ+bx58leHn5E2So8RvVemBNAFad4fbjFmpNFANaMLYIu0QPiJed2OgnKA/M
TZwXIqKdKrpAsZmOQNpQ7WebOSKLtYa53UDqQK3wkDg08YQRXeQfBvcp+lE05Dxj
XmiwI3t0BtyzbTo2n8g3mO2JILvj3FLCO6tkG22hfdWAKEUeMUpNFjNh3saW1VQS
94HiuWNNdtfHkzP71NqAbielMYcIGmqEi5/MszbXBnbh2k3newM0g1Os8m2+qauB
AXIDk0YRuE2gFtsDkw5bNJdWIstk9ndZ9lNwZrsq/c34Z/dW8aGTbPjAYX/hIAQd
omxBAFeXY1m9t9xnVqdspxoy1zBNC8NZwrrrI+BjYpj7L9LKqgkC01gThjX/vEo8
wefKIzobq+WK0yTXu/B+0yo908bfcqAbxK/79WLnQtwNM+Typx6IcVYlRGZplHWw
l+Hzlul1bDz8ml3E9ib0eoP0eZVdQdK5W16QLotLfb1AhOJztQHsPoAJLnqu3ZVE
PJgI60VCDLsH7x9c4rJ2ayMWBzoqnTg9bunYIa1Lzm+f8NGjF+kg6GGh2Vmum8lu
8mbhhsG5GcmP3Kv3yFlj+O9ib3S4A4BMNYHOHRbrpL/ShWXNrAuWJ6NWsdtsZc0R
y5rYvNwwiVRhMWpXp6ATgxMHUrhVxi9L8WkUdy9uiDwA4KTGxfmOw1HDTNeGQBZl
SlbjHWFpGlP8MfQA1+yM6bLvHA1MHnEyX4wtYvA7mctZIrFObeFCNT6UBhKfooV5
/qfO/Bo1t7HPHVKwJ8uQWiWr6Gw/ixia0QLklZptNV1gRpHp2vpDeEK3azAY0CN9
ZvKTCNhzvxQZ7PfkfAvZOnRt2Kvwi0yi8QUSOQOT0SgfuHSNesY/DPyiPvNOHwHu
QsjqIIaaj1Wle0hAWi8SEa7iVPeh3ZTDug78oFSLMGuFKnUFGbyrgHJl2ZfOs/XJ
zjcj6OmXLRtJzslzO5hmy5UYRfeXfFUOGl96nIgIvzVQiAna/HeJo3T8jGNH3Rtz
FBHC+saFwxD0o5TLKOUHMczv8eTZbUzubwS3T8iKuMK8BE1Mz58H4UJWqQkS24+B
WEmp3xfKhxWjkOGW7WQZcEh54OjFC7gJCepcwJLEN5vukFVtnhHcjCbRbNvi+LDA
0qQjD8lLzcNp1unmv4Yhw37sI2WHDMSUafJdqiW8FIdjd2cHBRX4vDD6VM6jRv++
6VoDOm0camoPSfIPI7gmCzvijtyY2+hJdPYaSyrtyDUfBfSzvUAkru9HIYBGmESd
gBlr4FgkwOcw502dEm/7uD6BKe9lYqaFtF8XQBSsWKU7emKENsSn2B35tsL3LyN+
eTSriasptMG9Ul0XAq+WyDP2j0mGAAlT26dCnZjOSGdD5Tiss1qUn5y2U/fqO8D8
ObnGjqnq69F88wLTovutI5JC/V37laitlB5NZRmO2Dc0qGEVYWuvmhtCXTSqYoSS
tkHMB91/ZsKqLNqbHe+R3rj8k1ZtacbZuRNBvqy8R+AjP3IskwZR6oB9zXIUclnE
0hZc+Yvu8R2OtA/xPmuybP9oOQEC0hiBg6MMjgLQBPpEpzGJR/YrA5a15HkVONHw
2u4YcBZos4fPY5D/h7PPnatTtW5f9YnDFZdYkKPQY051Mo6mV2n49gsd44kchx63
hyPF7d4OiQO5k0/eOmDEp/T2fDdZ9PXN7CmcAGWMfZK5IfgRpkrJXH2TJR/ityF5
fJ3IVzojpLX5tAm2rrUTQQLYguAT/cfSevsKC4x0dczlxLLKGyRdWUINwh05UJ5J
oPoux7wxmrOo7tTMUfb1MSd9wOs25f6jw/CbIiNefB9+uIPdLNha70wkCQYiiEZU
DousU68m1sSN7jDBiDn1ujHATBaysPfn2farwjbF5UUlSViCUgofS/gUE9c8JnEs
CXB4EGHH+hNXCp5CrWVLAeLJgE7gVIudfQq8I7roNYzeHalv6HFtpi2cZeB6hR8v
+yz5VFrD0BnsgYHOkoQHkaPT4Z427xqIivsnU7OO6/PABgL1buxOkYpZtGpNKpdI
53zXSH3TL0CM7GTi3r5q9iOg1HeDOl9DwoPEB4GTYFI6hTCwPzgqC1CDieYRDUkE
Xvk1T+CH7eb8J9OxKpuPWtkrRmoOBZLktwU5IDobdlw/eUyzBF+PiUFddnR7HUCL
twFcEGUOIvz9iuULz8yRtZYKW4ggujHS3ESbIjDmxGLd3BULfkZEANG2c0sD29p7
kASnRvpgiQcA5NA2+GD7eqZ8X9Cm1LzdhU9uL/n3tM0BaFkcm4+mSh+dN0p7Veya
Xs76Qs+wlfCzDEjcGj9RlpKspVO+tX8lE2bYZeFjS3PcLBOsjhmctuaVN0VT+1Wp
MoMaUOP+6mxwT8Jcpsv9ij2/p9hfFLa9moh5iLERqZiisgQvnKNEU6PHoRopZ/Qq
JOC6AlBVgSph+aSAsIEZYjJotkZCLFWdqB+tTjhg5/5ZSewzDxNI5D05GBtyHT8a
/54Pok0BvptsOf3vq+ARBp9Q1Ny4U3a0/cfM70lXjvQcq6gOZZI29z0U/Dfcp6sV
rlnBjnEn5YiSAiAEP4py1H00w2x6SdIsmkM+nT1dAUN6IWwYij9PgKmNMK7PGueB
ygs/ZWndvBsiyIQ//gt3U5LPMZEjeSXSajmKeroJRPZqSQN2HyYQTCHZVpo17Ajd
qRDj9uQknh+GNoY31sSEJXuTh4L/0DR62joT4t3qVL6Dg3fth05sm06TiSnES4R3
zZHkB/odX7TtzksB+5nlVrEIjRRnLhMOKCpfmz/geZzAaRxEFv/Ag1JJzb6hn6OC
Yn9TfUcExfcdvbFS19dhtTC3zegz3xugoNtzYLWF253OOv7hRvqk3cUWiKGEVofu
11fgPEl5c0REV+iPNKM9aAzv/mH6GKw9PuY7ePZxgDlyUj5AGnEMl0goIGjTrDh4
MvIaEmFBx/w5oxrZ9XU2ESkJLhWUHLxIMDQCc7x3znD+G6r5RaE9WmEy6JA+w3iq
FZOQ+56zSLdPdeDBkySYNvaYM/vUBzlL2pckKzc570YnE7S1b21nq2hRZbDKX8OH
G0TANEJQFVoEFVWT6VsVU8kbwrI3iT1FUvQWpQBgaSwR9e+uEDrpUSMS1rAUNUNt
xdLj5ULmnvVsDldgDP71Mcgk88LAdhxwgJrGqrvZ3WnBtlCXyCkIO1G8DbPD+IbC
+IyFjXAvhX5YjjhyCcwbasRdBCiOW1teOZXlbtBAn4JiYpn5aQBSJdtYAUYQpV3N
glZX6shOyUG2a/eCTT15pAM5uoti0hA5cg62DkPzHjglOnrMQU3S7rWXQdr4DrY8
RrCGphU0QKgYOK8DX0pH//ZxSDBtb9A+BHLvGyW3OZMzsl+nl3KjYEt4vZ55vg7b
Vf9dD4B7gPa1ZRHmLywcUOP2DzyzWhG7gG2mS6Q4V57M8EVk2aqLT0r1HOsF59Jw
2uX8hvDxPtO2kDSgIHtDJSQ7oHffZfqoqc/rd5KFFDo0qiXLgVaYtnxZaM1Kof1f
51XTvxEy2FnVasZJRFCSXNXXgDi+0nXTh7LAkb/eG3dCjNzMzDr5kBlaKT7mrvf7
mgEpgPrU1n7r04dMwWK3tylVtQtGG8d2VKjMd8HkMfXmVuR83TMzoKl+56i6Rup9
SNX+j/NGDNBkBLoERXFncFsuctoCzNFGdQEDxc/d/U94nzRmxnkdnEXr31racPXl
N3XOnqZ6O4lE4XVq//L10TtFVlo5ns87T6wI915dgKd7tSaiT+myok5CIcoIWh+P
u/5nUY2Qy/mRYK9SxfBhhQdUCC/XeDrAvSEQloqn7T0cvbimX5LDMrB9vpcbIOoD
tcpdoQBheIqtj4To0gMJfb3tXKAmfK7CW1bIi+nnc+wAnOf9WEcBHfx5/HIsJyZk
ZgLzYdjvS8kRG2imACu8LZYX45TJkreWor2C73N4NX6QzHMp/qUmGqug0MViyFOT
372b0/np8lkFxiNRZUaPEh/wBtIX5mMqPKj0HZe1vGBVuFwVVfjaYfNgzNYsxRtR
Gdn43GNKKxeat/DHnUhnd20JLb8Zs2s2AYQKLytW9X1PhtGs3iIfAD7hFA2awkxi
i1FVIl1Qmer0W0uVuqaLwgQZgZySttllabWNWZJFAqslGMcB6aoaS4z5mV6g7Zwf
YJr+ZABpHmVCauwwVMkdfDl+S1j4wlFJHNQ9Eb518m/DGxQcvE/O59d55pwUtv8+
1eQdPs8p9j11mvo60yNzNlvRBbfyku//MF9SEbfcD4gFmJvicwLKFUsEorjydp9s
RAA6Gdrsj50wGanhInr3gjY+kD54rAmvtUGxFcNNSmImftzNMJrZ+yInnpRqS91v
CK7GGQOoGw1dTyqpJXtbMdBoWqet/qEOh2UAWiB/cbeUUkfROhxgWzYftq+wqd/E
jfIMyBbo8HRF81LVThgdeLQKhnE7uVf9X7a81obFFGArzE5DmvZoZSfYF7y4gstO
udwSjrJ99Z1r1XWLgXlIQeM0n+EEB7gY98hMZ/ZjRb7CTt6iLv85qJdvPa74T6EK
AA6zsH3TpHYvXLIZ0tjBgsmaZL/sSA7xrBAFdHssatfo4BQenf0jM60M/omVzukN
+xI8GdgRc0mmPqLi3Wtc7wYnfa1810KW0xkagLRM/cCTRwzy9MZQbVSZDxaIHvQE
cIrkNo4KOl9yI72jTdTj0sOgt4o8dHa+J5At+O7DMmo63vYkzDgSr+f5gZyjJrF0
8lnTDjYiQVybM2GlKzaG/wDjAtkCQMSyrmBZMigeIJ6Knjfhkn9JViyZnioVo4/f
BMVBOnWHwrRGUJ3d0QZC2x4cbY/g9QgD/F87J6M/CHRlHK1jBZpgZhkFAb4D0qaj
upEaw23wOfbeag9mXfWju0XVwnW7eft6TfRmRJkZljxXi+jk749YQjF46c/L5qhH
9qigTBvPwXDUfwX5/kSshCl4cokQoiWrkF1aJ1k9qrZYaru4IVx9FxXXuCHTE2OP
zPEDxA9O+cbiGGA/y0TdRf8Uxl7sDHz008dJ8DQmHmXhEfcsiAZZiJw5j/9h4QtJ
UMGecQdgg49skzo/Y8Lm3CFpw++PuvK+CfoN6HDr3u/fHQ7088cUtZp3lxIkaEN1
M5ivyWHMKTScMITxXMGy/9lWucfdnZvemKTIHRHuYnJ89if8h8j5HVCYxOez3V8o
0Lrj2rZ4AJmwZcAjznlMEvL5RfnXnBgwAfbdP448W1nQeGt5HJNFkkPwhSh+mAtV
A8GzCEY1E0EsUI2A5OTHN12zmFaN6GWgL5VJoY64c1HUOsN6negOHwBVwq8e6VrO
MaS5wmocVfIHQm4tK2FmKcZZtsb4KmfpvRcB1b9w1ASALsv4bnMx2tmDRXGHwPXy
9ErH9AynLIQD9JFcBP2PQKlpcJyRghp80S2edoHB1zhLQf7Ps3wcp3CyyNGbjARH
iCKMLQR1ZgFNTS75cue+IF9ACpsRS2tt15+WuKPGYYaE4aFpaBO39M3VwUQLb+ys
Pg44Itbh9uQV8wk8TY6FR3mBWF1nZkcmeIJTXdkgFXJXvtYpBLpn5AguBmYl+2eI
iTso+w+84p22MEbfjjv7OmXMN0T93omV+pnr09HxB5ciOk4DKzFkLY2skBnCzrLM
KfoI/LL4dA4NM/wZRO7kFomW1yZTRPncdH2Pmildfyj+oC+VmZWDVu8ujGViiSIB
So92TsSOYngd7rDX7uVeYSBZX5KmAKd2KiWkB904coUfrmnnlAzyXd8avbpO52ek
FjbOlRWAUg+WjpEEoOxWfzjlqyPS3TwEZXauj7FbBqZ9nyagtDGOovFzzYNmSpGv
lAoWcGJ7IEsmsNGcwKjlvvKm53ZpEqaS7MhhbTyfF19gLV3KaHE3hA1oIp+nA61x
W1fec5nJ+WyoFPnnQm+uJDexh1XGWsKL+CiPqA/vD4XGGNNNRRMlT722MO7bnS8K
l31TiMHymi8iT1n3Ml6rmVxovAcrsJ3QzA+Q4KNxtUJvRktf2QTRm5ety+A5uPgf
saFx08MNxspbNAYgUlwfio44GtM0q23ct+R+EkWyCiUoNG0ge5eFuC01OtlmOaCe
buo72U8ij4D9eS+aPrpxVBcq1qY09ixIVDH/QhRrBcjUsZNkhZpIn/xRyUCpYv2t
pR1EIFUBGoVtee7vM+yZKH+ydDuQoibKedhUvW7VaQ9sDB/6c/gIKyXdF5iyUS1A
7gC4wRFf8VdxHHYgzHlNUrPI9ixBsgDLnIzH/3WluFxiPMTiEEw+kZQsPA6VhFjp
siM//YmGXCe0lPSEJVM6+wTtZ59SgnGMpFLVYeu0UpzyE1GBxWkj4dXuYGHhYa/Z
xO9t17YdRsXXueztJaKY2Ja0fCLBjibqCyxrpMpAUa6DX/tlzmy/jIxI7Z9tavgz
4KnFHfHxpgjLnyPTUBJgEUiuXybTQEBohjh1Li8IpygselYTtD7JeJiST/6LEIP3
6Ktowy+9AJeGxFJZqZOI0ZNyh8uliPyVXoEzsckgC1l4/68+BdsO4PsjS8Q6Ydrq
VP8Q4nzeu2aONQSJJkGPdU8NdJZgFzDk3WZq5jeM/v3l8Ip4rXJsnb9VUJA806iC
51kM28nQZNR9lLuP7YQkNjjId4bqqGnBgjLpexcnQAXV9s5e5LGJyWdqJT8nID2d
Y1qvz1fy0jBTEEvc9sOPB6n95yZm7goAIkdifExRSDBUPfHSMFiqh/MsNBgf7ShL
devpSjwZ2Lh4gpz8fWYfbi3r3xvJgLRGnlHW3oc5BWyojVVDB3mSVn7vtDS5e0Bq
RZoiUVYhe7IM+ER6uU2xUrjFscu3ci5kps8XqexNEBLLU0oQbEy2tDP5zJAY/qAG
A4W0t/s5bFyyy60CIVB/0CNWUdcXlQlLEXYxdPVMTANp8Pyk+mUXi9zhwjF9h5RB
oVhAu5RJ3Mp8cGfcSMcWbKS4q/UrPf7qUZsR7WacuotaN8OdWfcah3JHvA+5u6b1
m+3IUg6VOMXGxJGiV3YNRNE1EwmUNa8hfh+r929DMs/sSuyyyOmfKJpOKyxMb/bL
y6D5GMhoDgA/Sx1PhsFTEuPS/n0908vcQDbHUzy8ZuC+BSQOKyxH+2pRynIqeqzs
XP7yaMahWHdyKReh0FIVSa/7dJxeT7ZMAd7rDmwnudfRBkSAuTQ/Gch4R5usLHA1
sYIIS1spjqpg+aYQPaicJ472Tv72UoQikmZhQJPFqljqsKumgTzVuaD5yP3O/527
w/GbdnZIl//QmPMyZLWf/qhModP2i1bk9Xsd+JIm8Gj9LPt3MkjoHlG1TNuNHS7d
JgAP4PcGvdSh+bnDzV/INBg7FaAcMjr6tDptL+w7p+cNz8f9pXy13WC39pJXx4va
9pLt+iOabnqas5tXgOoLB/hEwd7SNrjxsgHrPpfgC3fVOhfbZUn5gug9wb5LEgMK
IWBw4Qa9zVvjf3KR+aFpJUGFyh2YaIuCxX9FQNVcwCL0RVIc6vjRG8yUx0Li6exy
fhNQ24so6mehICHV44bht4iEX5pTRJYEPobJ0t2RTvcgBTI0852nOlV7x8hMIqkO
csq0p+sYSoNKodYNHkxV/CQIjsIum8ZphnIcLK9ztaKM5HXYHKCnyqcxtxORdoFD
fg+x7PH1p8UGrKc0GFpHHGMJLVqjLXuPIRtptw3mDiijSfLCxVFGiXZVUjKxN6UN
1XjueCEV9NVXLEgVaXpSuygROvyTL74U3hRNYu3nKQDghOW2RcV6FV1aGzZCwkkG
+afyyTYwjKv12+QatW5CiaIIuFLc87bJjGjTVaK/JRYW3qaXIRlL2dq3pLb+SsnH
gQw3YsnDoOU5SmB0dP59PTXqUy9Dach0HGHBUIbKlj1hcu4RmEU8UeJF4PSvexyG
OfsDVZABlf3d5YIJojXHuJSUuO10Q7rMkA2ju2ulDDTWuGriEkpnxdNld9m/s3mC
ORZcsZ/4x0mtryRYVcOXuXxLSDn1IIJv5vNTaF+17XyWChwLbB7bv43wlUQ6C9h2
rMeo8UJJyPKBd01FDfCP3ZATTvJ9Qy5f46tICRykVGd5dDUOiWFB5WD7jSR91hs+
Z4u3zOGsxX8vDzb0jRnh7c7h1wY9Pf8TFNfZxR/qMm5cRNrXRsZ5G2zAEBf99XLF
ll0T/wZt+GZzm4zMS1y/darpXSl/XVkMHfqOWRNuBzKLGN0Bzfzg16gGyrFInnMm
4IPomWbwj5DhmSpqeeI0Gko0cYS93W7NW0NhN4Pj4OBDitPfd30Bp0lLcUnUrBMb
1HfP7jvxFF5QsRZxmsDxT+ghAX2Ys0oZPSMIAaLk5ZzbwBWxiMzvZkG4ndrFn+Yg
AniYt44CWktkG8egaJOyxK2/dJYjGCHx3hBWV0KwIzrYqlPtfQ8lQHzL6pU0YbYU
RpslKT+SqaAjQlTgaEf/zGSN2me7ybZ8QTs2HJy1BpvEOqTVh9imD5KYN5jjI4/o
/K+82bAkeEvfr4caJrmFOKT9I3LcjYbrbwunAOrZoRFqxpBFx8VfUg/eBZSt/8Ur
zqhWMYf68eSiDUiAhs4/zSOdPGhMajaX6DS9BHgwcti31mvu+RUmyEfvAv7Mg1iV
IKwnAurhMwbnmr5lrIUd9MTcMBPksgo18OjcuJpl3YLMLo4GrJcrOg+DwLZX0RPV
qO2zT8KgRJTNy7Yplr70dJMalCIv4gkH2SKfnrd/FhjM6RkznXfXJaYvPmI4KG3r
MtYDhFKrZ+nNzQp7vt/TvhqgNZArmGSuobaiRVRanrYmVH9jhA+++2pcdD57PzIQ
fNltUD9MIFbzggHxQtkvCRk6u/oziXtd98zSqoFR8TDrPsT4apDDK77hK3GBsQ7l
JMCy5Pjj9iDHxpIH2uF1pJNPUD5tMGSV6tMC27iI8CkeISKnN5+3eINxEDdwTmr7
qfZQ5Th59s9aV+sTTvgAcCgp7cX+Kw0AHeErpZVopzoh/DfgXyXhYKSE8yS3AfLM
6gRZNAx/dyqFLBlL4/lpq1eXkSlAE8KkdptAMUUpvctElGX2hjpakBdWDHkojEUS
OOU9CAy77Yqy4pmE4ECGZnQ2OULXk4f0VYlnkUy9SaRHl5wF25yxnjJCR+3C4urN
rrDZhK4YWtNot0t6gP9cOu5WchxBh8P0b9UoWPSHv9dpEBBD2WTNzEIC9ud7Y0rw
LFcL+aM8TsAZqhuPYv/B2tjG7m5DUYuiReyS1BP+BLQmkm743qB/WhLDub5NnHaB
TTaxVZgqGQFgDO1827NedbztVcGdJ6n9Yz9N71em8nFInokSfIq5KJFdbCFP40vc
hOkR+vPSIlV+oj58dfaM5K2tcjaw3u1l6y0kdeLBN4XEhbCE7css1AFJ52zjNGTe
x3H3/ETgnvvrXL+JXsSf7LIFx8+S8Gf0yXi4yv8AotNq4C9ast7AERxLhBuj/aB8
yH/5FFUuiDBYlDk1MCOAjlwxy5N9piisCWkSkZeLDTwa+coDpcJKtyzDspo/odRl
vjz+kWyMSk5KAvTziSh544S5PLXY8ZqU86Gw1KZ70XCkNNLlzFiQd0k29FN6Vzid
DPk/yp+A3d0350gWz27m42wPiR4Nk0Qr32KNHA4CW2fIu+b9Ww9Br/3ad7Ds6VyW
UnYauqxZtAD5ZfCmmmJUk9kOege/CTnFFkCI2dpbIpuWW0Spnx6KSu204nUesBa3
gEV0F4feQxftguhuwR7D4OYc2ZvQUuNqM4Uhs/cMi4b/48AF67Lc42C8/XGTHHcD
n7VVHhShRJF7vJ0dOF3ZySs8eYCBrZxy+qPZKdH6gppnclGB+P9K9JAWY2Id8qSZ
zJ94BWdppaPgUXY2lS8JKNx8J205hVHBtxlOESifwuMgQfgkfRYesM4yAW3ptDf2
vu9uIP1CFveXwlHDumxDhTD/qDW/IvUAnIaxlckUt/+kMvcckZDZgq26i+/MWY7c
FClspnRg/D4iAFziubAGRPrUiS/mvZZQLf9JNspoZT13du9W/eYPt3Fz1pQGqEe4
jFWFdfPzULRFp9ik4piMxhNv7yWW7rKYFII8stdOHbde87YPtLYq0dXJ6vfCVkpt
BYrm/w28DjK9bUUZILjwNx+Net8ivwaibV5pyLPx4GePQtyg3ut8anEGqafZAohW
rLk1cnRIVDec8PA/7raf5qFg9bUwaJkyrRyViJtcrUqzG3y7Snhz8FYM14GvnXgC
IpLBwhXHuGNVHoJK/MTEGjE1zC78yqiXEYgMPrlnbPy6KW7fw77tXUUSuXCeQA3A
JU7W/av+BYyrIE7gmr8tVG5SSrb/fjtiTJQL3jbhg1sbRmW0c3KGYfoj4C0NYVMF
SHv+I0wMzUWld2by3tCNdWiyOaT/GmyUuPZJxnKf4zAYzgbZg4V/SQl/bK9aOMCz
w4BbnsuU1Lms9yytLWvx4Byt8hG8XE3R72u/24beTz1Zaywritc9NUX7NGRWeDJg
z7FKy1F4/NCXburryodOdj+RhUKWfFHf/rZ1sVdFvat99cFJK1VYj0ezRJfC2maI
1rg0nNdZTJCn2nBlnhWXdNf/EKnCl2keaaC7jzAF7EnD38/CV7MYzgHZNEFHxrwd
vizbsjv4k64+Hajl7kRw/JzPMA8dLyKXeP3YCGZMnkZG0AWtV8lDdDsApthz6WCY
ARDedtJ6qWzjFpBBmUEWGIVTqvSAhK2wd3rVYTbmdDzz6bVX4aPRxHsX1/CzTa+L
n0tQFDbQf6aqE8sTYGMCBFWZnryrqlPH2D2C+jCUvo5FYp0MPFCNDXLVaDPC3Io8
HfhBGjVhUlyaLxI5fjY3ew3yXVNlmaIs+BtZMTVJw/thSZ93pUdu7b/mAC3NTp6j
sQB0v+xyKcSlziFry2KJZYS2cffV2sVA5qWTofS8b6oQnbE2IJkU9YKLn0z+Khsn
+36vSGnQhrTb/osr14Lyc5F7bzwV5ox+teYTpQddneLBLz6+OWPbqJ8UjkjuIdt3
snzsX2XaAobHLDKvvUI6/PzH1+LOuGsTMJApyl84tpz3/8Nv+CidN1ZO1F8X+qCu
kBVUDpOuHqf3uzbcCT8xOXRkBx/5d4c3fF64ahGyKAFI3YuajoYplJ6OBzIKgyOj
fnpyhfK5mSbFas7qO9nDnbcYq/a/bk5V5bd1WoSpxds3M4RPFg67CWNcj3PZBqbc
f+ytWNueUigsVuBpeduPW8ZB3dpn6gpMQ32z9gHx2Yn6NoRKz1kFe9vnZVGtYd0q
J70hzNbZM5EjITSn6dqyOpqVmFx6K78TgIL0RW0hT3OkCEGx4FPnDmCu5U0i2KDm
tNZUCDRt7ju/DxaFBJJK7bAxXvz54MU4A1fE+lHJ5foO4kymzb2szoXupVuI3p2q
TKi8AIY42XS3lBQBqqRmzwtn9X1a5328q6odgzCh+OxpEJEJ+oXux2BJVaeqHAkv
+VuCPcZT6GfXwTDXCK1es3/Z6OomATjLnby48+64ZGNcPVqeL1ly1PfKTJSO/9Y5
rtNH3YjQSuPQrCP2o389mi3Ce9FFV/RCPnzQdlFkCQ2jmei0r2jhsjukqaOEY1To
uxXFrsWmR5TQczNZxpm82OeDBMWGhoUKxDODOZG2HYuMSs1tp5ABb8SdJQ9/7TmV
5BSJez/iBY02uhFK1odAX/JlHlh4zrzlKdJF1a6C8MNs1cS2z2L/SVtZ7m0BcE6D
d8fV3rFBRwobVVjtnAJaHpuDO/SBnoLfE5n1GweuPSrnL53P69zhwB2CObUXMDRi
0lLUr0zhCDlloKyG8LWNmVAj4vjeCLyZ/f9Df1cEIs7+aEeKywG/9cIKCYRVIZEZ
yZjQRji0yTrsT/akAq9Zx9vBBqm7OxtBa427yAxUETwpBAbnnu0DiF4HY+eIS7pv
Z4Yb1WvUK2v5/7MQxuguDJ/Fs8xtt3lHC815jTgLZW1IJ2n2oYIY/R8hmwvM0nOP
ww06MV9fdOwrh8ClWXeR2jSzDaI7ru3LXjRD5QMzgvsu0hbMFOns6MFPY0n7J2Jr
9/TtHKGFnfGu2Fh41ya5PggLzvJt86Mo0Zaqt4aql5nx5fzIBx+JPT02gkYswVKL
5z9BabY1JucUAZisz+E+TWElMULvm6wfCkuCLC5uaNFrTHhNZt9iMCOhaBZ2ZcHO
FZa7Qq69CmzbE6sG0ffZ5kvogT0ndKp86Y9Yv9/i+3PEyFsRHhY/XJhSwAhTBnMI
AnbZrPhnJCPJcYFqylAt1VtuDliZr8CKGqtfi38mo3aFwmoV4fTK68DI6ZYiie4T
fo2ZJS1q0bSXgjlaMndWj8OZZKFhNRB+rHdm1SYT3uSXjB3JT9GrQ/S2Nw2aVheN
fpe5v52Z4RsgxcYjGzF8+7R3HtL8NK2eJy8BedQFWFMwlQ9NIPKtmDdMUaW1L8xP
uZRAGTZakjfQnV/8mp6boFc+eFJnOCBwX9AXMCHmUApMV2CGxblpM4f5fv8nB8cO
jKQ7or268fhs+I5eta9ijxr1O43KJBKBB0Kf8ECkpx0CLIQ9n2rQWvnMX7bEpBAM
dzN2qgg1HekaI/PPZ01wcxah7OapJ2wlCaxkpgvcJRcEjaUPh4OrO4eWqMXwjiGG
uGLHmBoTu0gcJpuEFrhNHf1AhSZs1HdaDf3etiJI1TJPzsNLDFiLiYoWNZng5qRg
L8Or5mkml3SnxhvRsSpxlw9FY8lzMoQzmh1U2sWu1P6OhV1OnEMdjkcry+51lvxk
PX93q1CX6L5Bp5xyFKwE1B19KAcXFAFdTVDO4HZG7Qg/nYuSXe7x6XvZOAJmHy1p
OPbhSPRYGIxLmCEBxpMawEd5FJJUT0OjJlGIdqEMDHX1GjobO+wGjL6AjEhycmd3
DbKlUyN9ijCOEs/ZQDr2y/Th5vMBR/gs1iNaXtFykGrtkyO0lvB+A3uN6JCEsK4C
EW2ciqVrS3JYv80D/z9XoiWbm67Ec0lGjNeLpYRf+eRvmW3nCvPyRQIbrAYpak3A
t1AjjYpMj0zCnzYoeJuarSuAc8RQj90ltMEWwD6jaySjp+0HoeeeFf0F54qaRMIc
popaVqnkCgaj6Oin6CRNI5e+Z9Yg8yk1+7MBFIL4X5somnJIwuWrvQrhDXnEslQ6
svzQVhNxEAW3w1b/o4myhNOB9xsUYswxmj5D7bFlhinOZhYnMXeTGv/g/LcI/99A
zxlXXU0nGmsGL99Rg2p8W2XYYPfb86R5SkXuwgGQV+LIOcDnqL2wAp9vv9wOCsXk
LVO6pcXcJ4sVKXrVgqJq/ievODaUjpWrp9uTC3/80r1R3oG63H1MHOAgb6IWduJV
NrKPP/U5kFijbBp0ng8q+DhnDaYnnT+xb8aCtuXs83FjJ/4CiOICq+8eABcbGfFQ
qnIjatC5dv/yKWZD3JvEBQIAttlYKKYlOgf7105NwRnNIZG3qN1chDhAHAJymP3P
NyPYO65n28VDgZln7VdeJPekj4rl2Xp25ISi02JkPnBwZe9W0SCxWDs3ongrudin
g5wTr6a8SEEw8xdfOZz6rK6OtHJTinc96OFqYRVgdbZb/rjwyepXAcj2F18yBcxd
KLXyn3pvzB8QlFa13A5XPWsYwYJrlQJEAgsCua2BtJEnrzqetD2GXAUO6Kw83Jza
mQckjljReodkD4jioEiiM0az7ez6+7E7BvDpqzA6q1TFXZwu/SikKQ9DJH17KORJ
ye9viVrm2aZnJC9WASVS3xrS+GGF1w/DCJsw8b35IMQDxY8hnaqyJMRExafQO1I3
uV1WzIbrDxpzlh2im1eDC36ShPc6vEcjQmzbCwl76Y5R6mJaBy97v4eTfafK/ELP
i/vVtsZbbx2aotvmwHh6gNSS5jJKnBU82IRQvhNSGvaXz4USvx8pXQDo2oGahJo7
D2x2wVFbnvT2zyxPx9inDUPmYThUxXeARz47nu7I4Ip5db5S2q6hVURgBSV2QEii
tbF77MhfRLz+6NRze2XNamzgQLmQ+FoSgVWlaVlMRENAS5H1t0Lt3Jj6ulXgxjkZ
WsbAIbVOBclyl4yDhQ8FtWJaqZROWdFM4/Gt8/xWvpE4CveQHh8OuBsU3hasHYZg
AHjEen121p8qPmgYAFHVC5xCaFLDpWDKeGBEpTmVkK5kKhTJwgmkpAZIj8OK5H5m
Isk9jeK6OzekZqquPIQ5X2Ou7pTSImQZXEXGJoSi0ql2qF66h7Et0tqL8wFyWwlm
qgdB/ubv7PFGPoDbLshUgNDvUD94ilyCN8cgPT6+p67z3n22CHyXp9RwwxSo8815
fXO2u5yPwygwIgzMnJzijIGVwCXAVNzb0w0BeBwYdi7JZFd+qy5oQxF8rJsj0Vtz
QolbpfNfMj3+wXtL/wAjZPZxU1KciNPkvC1zqvVWJxuk1eUTfs2aZUOwBhuA+N2a
7YrtFB1vlOYOEAFg571JE6uqQmnuPu5T28uJAe4XBWCdTFoHUgYgkqeRJCtBjmcO
ygS70O+o7IC+u5oF2ho/M+7ns91gWCboW81wTWAZw0w34+uwVsE0hOXwl35tObKX
ytoPxb0KXzlaieJKyErJoJGseyj6g8bQIhVY/nii9Goz94cNkWUqKwnJfSqOLZ/L
4aQSmjeXGjcYlT5de/SpVRL5gS9o8CteORA42Se+LiHw+fhLgMZ1cxM1xtQ3DzAN
xEWZuWNwbpi3FiBTK3rvCxZzeo5cidqoAHm5UJmLy1Pba9+aYtKQD0i6OL4H2i2Z
y4qOquOHhGwRA4w/KaWNXqfEV3Y9IPye1GJnTwHj887KI/3sQ2hYLaa58NOJQEah
FshAuvyvx1/QA+dW6cRpWdZO5jMf2E4vmTetVFj/2EFUQzFRo7GmIeLS5LP/fpPA
kjgEksgJWAW2EPlLx+KHStWZSjmgE5DmopbAe8ZCl0vwGqBKiyMYmSVK1B3KyYr+
OTjr2C0HUG8orrOLiqtYig5SJmTbb4Ir3s1cyS82dYQZzXvk9AhoqCJ69mA4MJjX
MsorisvZr8ukiP7ej4x74lpSsG0qhC/OcJrfOmFx3hffUx4FooDH3SZJRSY6OJmJ
R0Mq4CCPQLEpm5n6Dc4oSZ50R5EoLkv/yJGtJtAqD2NIoyGFU8aibxSiAlQdkBs4
+PmjZhwgqTUI6ruNuvMPUn05wvWtAJRufZjjQYby1+9L6fd8odr6OtxBFILOuESu
EOaw8MYDOnXQEbiMS0vuBIzDJBr/QMx2obbC6tr1EYZwEenbGBu7YQJCYvQxUvRE
AfyzYkbUdS4eGM01cj67xSBf1oZmj9yf53CFys3XMx5XqVDHht5Tb1J9vOEemqQ/
/Q0Gf7ni12Cxpi/I2y8+1jUHityXilAsgY7URQmVF+O/oKm7s+Iox2B6XtQeGvSA
sLmIzq5k0FGowTDZoQMPS/MX+PyuxkL8JKZmczLm3waeNBi06q2/5dQqAuDy27RL
DowwWkzbVhXz08XWIdZbS6W41eYCxZk6/YJ7XRHhorQroQdWoKO7yF/YmL1TdiYR
+/NMrqwnLzSuoSguVSDd1e1xdcsFvlQp58f0TRRrnDDp3/2gQ0d3nIus+lMVTPrP
BKOljCybb8Jg7ISBlMG50qAXvshZ1GZ5UrK/9Nk71My/v1Wz5d6ss2jrqCOYU0HQ
253CG7U6v3hyzGw3tgWIL4ojrXc0StVpypSAplU223FMIZqXhz8AcpZkZoo5exMS
l4vUKofEOOQe1wPaMfafyEWrc2GdoxGHBKiaialXSvbzofLLnjHC2qTCLmNR5VAv
/SUFYLEl/pHdowsiYAr6iEudBHUFzLvgmoupZcWoLOybrjiWNHHDdQaOULNBTIWm
dU4sUcsS7XAXS/JQlEW8O1LwCL18pZ361JycXpD0l5us/wG1eN5gSR59PBGVzLDW
7UwEusTpR8S7GSPAW8iK8ZtSICxsqYwUsu1qfWn3FNy16izm89FsASLfM/cStB/J
I64g6s3h1voie+p08uUTcaIH43IG/hi6UGaQ1m6IBmSznFTNyHz0v7tfK2OcNjSb
E82gM4dLg5dhnrXFh1pEuot9j+mLVOs02SQO8OV+fjo8DEffH4TAdbuhRnO6qGP5
qRt5BNqIP8V3+XKLI4AM1f6fiA8MdXDewXH3smjUU9NhhSo3zhDmyUkpHS81UzT+
g4p7QmwNm8xPdBF15Z+tfVJXYpyEfqXYpUchQBHeQSInjHByOn7EMrL4DJRXrjsm
/HWqcPwZmSer/Ms0fXG1OJIYYXf7YSpMQFEJ1hYGkEF9+fB4ZM8lAur1AJPIHXtv
arvsqLLG9NZiRRRV7SrWD2fi/RV3ciZjskQ4P+xQLzo+ZwZvNZZ3apN+urMB43bS
ZUr0NfZfhrItP3P+2nmtr1Ihm/DhuKWELiMo2W8wuBYxML5pU/cIIg0Pgo1MqGDN
gyInQRGzamkrtD+ID4gmC+xsxJ//RtdTJ5aWZUJl9UIK242WkDJmKxcIA5iJlAPy
RpDNToiO4vUWu1eVZEipHHX6ruyxLePhSXMk4BEUe0+iw/a9AmKIGQQsUq4AqS7t
ZJZVF7ViUSvQ0Ey9bA34s6EdmimLWPZpqqkpJW7jn8WynwLxqKwnR8OysK12d+eD
kejrmCrlfL2/J23nB6iBdcSgRjJlSL0SPor1SvpExX08KTdgDZddioxeu2g+0tcl
XN3uDDlqDQeOh8QR7lYf4Ulg97jqbpdDT4EOly/93SfSOyHj4HqJUpRliWkZg7+L
QmPHPH7vhlA7gLH9Ek+n4x2Ihs9q4L+DWK3Pk2CnOjPKVyY5vlS2p7gU7Bb3sfzj
aihK7VgQA9rQ9m8RYICY/jxLC253U0/qkM+bbAWMQftC4w1HJ7Fnnz+wev8IGZk7
qJRoMyVYZ0XDKVU6eRCSkO0GcKLKVrkzD/t7iq6/A0TY32frV9Jsr/4yD/v7iEMG
bz3edZdkUtvyp7re+9EruSDdeEA+8r64UcgGznAsr2IjUQaQ5HGMJ7Ug31/1j1+G
ChecoAYv+0y8SBmyRRzYN/7P25bFEBIUMRcuFc0uGmK3KilFHMbnFkQtKU6MYQqR
dCIvubUmF0D01Qq9xEPA/FiaiylNJUsBSUqoO8iFBCWlWiN43pMKSO9x+rw5+449
MdQGfISb0tiJaxdHL2ccwDboHUVMkfZaKZOg3STWbFLgfUB8LX/8nCsztpIZ0G/i
NZUuLsAHAzy7PC+b07RAwlBmSV1UtghWJU7e+a1IV1QPJS2k9/ytc/JgghfRrBtb
JeNdcP4g1hvfa7YTc3Bbcb9wqP+I6BKg7N8YqRlbrLQUazwOLA2LZKASzlusC30A
QaqruPeUmsbjesbrq458QjZCuqvEiqYZreFNJ67IC2xVxncj+jAzXR3iVBa/MV1F
j5QcHFMLz6avNES+ztomUDgIwZkpdOyMb2wdyp/D4lJcxmnrpLTNvkDWseBfDzaV
lmbvwyGcFnigu17Heq/Mue3IkyVSDDm+s5l47JeLSI5B3u8mbsy0Z16oVzpayjKb
HzXKh79qcu9HIMs5gs7LsIYyl/6WqyeOCOAb9nL5UYPGvCE03S8+WYr9+hB01VGe
xinIz+ftoFwrxIzpIjgJMff6cf625GilRH9wS/ENlRj2CRr+OkwM7w/1Hh1nObPp
DUyTicyhU8rSh1M0xFbLh5XlY27PtF5NRze/BCWSvzi/3fpi2+LQtE2hnBNjOZx1
8woJOvvAsqDbGlKmUv5CUVHRzksKMgcNp0vttt7ZApsBrrLa/P8YGRu9d+WIeFX0
s/dHyTblREc7qkwXkYv7u5PDP2g3O+ammj3av9jyd9UOJhMNDVmK/lNTb7xxI1hd
g+N+FlW/+KlvBApC+5AxLU7+vppLWAfcdK5vqeY0lXjP+kPCAiSGkRdCMBPUkENh
xhEolQzq5eygzVZ8SNYfg+YF1inU766YEqyhBQsTFvRUViI33Yfw+IiXmTjwjV6S
KmCJGaFmfINFEzmduDHvgFRMAhF6UiXfyI0XtksnX9TLB7sm+N0VNnMA2IsA6k3k
ILfL2BAlFRpJU96KA5nsI7dEb+3YZyHKfq+QyO9ZFFIWHVVj1IGdUkp/y+qj0YtJ
9rCpZn6twOIg2lRyjfa4c82OWFH5JpbIJTxCj75l/4+Cn6c9AjckhxxquEyjOVXW
PK/0tAv67c2igKARBsD/lVnYh6lvDGv/27RbJqExBbhOR51afizZ1IVpX3ExZdPz
4F8IUt9UX8GycSTJhzvSjsMt3LDMXSZ/z9lvI5HSkFnFnCHTwapK2IWulRhQ74IE
I6C7RlyQDhMwcevGTQJQPf9fGEpyuZV+fAYD0jgW/iWc69htn9xJCbeBQVxOiomd
7FtZAAP/XQnW9wkpZdAmmIrh0LJMobNh5er9v2Mkkqll6RxtoRfDBTIzjKNPV7/+
M8ReGTh2ZbU7qF3M73VvNyxf1Ho0/wP/9sAmRXUq6GJ4Wv7c4ruqDnrsvwlX3kEQ
zzzsR99zsSdxmVDIdpn7P3bKo/k8tUivAlWQVBD5Vdbn3HOx1/RaCOW9KgaWbJKc
Vm/7spj1cVH100otlMJOohyX7q1ccRKp0CniVfGAfRzXmvFsk1WmeNCewHdwnxAg
lY2g8+IYJS8O9kRVZQPtO41hXFn7TaMRT1msBL0bb8vR/2xPcjwGHtEe2821VXcb
IspWX/l4EafGxfssx0wxrClTAEU3jTCRPaybxoGiZspfTeBMiTSF0tcxIUdXfwVi
rvgizpRw3VVGZ1MLDoBu9llPeq4MZ1ENxV2v5CiNl+r7Q/SyOYBe3bMgNBub+blr
8x1UaBvbOIK56WxNKbLbsa3X+0yE5W6oq76NtFV09uVHpHgePAuyB9dJDQdgaMjo
7ZCuLIWWZ34g6Ram7M5vNcHwVrxV99Z76pRWTVvFfY9Jw7lQNXI7cM/+tGs6fPU3
GFimky+xd8p9HCUdZKhDTKyz+8C598DYcvqU9YQXMxYUwREbsVSpjmCzE5yAeRdi
ZqRTn0gx0gqlaMVKqtLTp/qzkaG0KxiQTvgvYwItZU+OVRGYYB1gfw/Vk3UFfmJj
xSjjJYOetKHmjptGrAWVq+Fb2QxEKgmCNxEPUX26jUZz74IwSY9If50aVyFDXnsO
fd3OeiER7qjtiWXd8AmAnLvC3wWTfqQlGWlpTW600odeh+3v8Xp9zK35vjVrRsGJ
ulTd7s9zRuLWXqo/drbm4HLv19QJsdqboNy4ZHavLDB9Wqn5BWuXwLi8F3Gedz8c
aOenLtkupmbIP2/UTjeQnw7+AgWOfhG5VnaXb7/XbL5go4d8LONOkJWHnC7MguC4
x3KWKl0JnfNoksDdyD8isOF2ycGfPeMTGoRjGZv/Lt8ap8MY8x35t421tUz2vFMq
3ovun05/j3sdlDsNh6pzV3oRFH1QNVGr2xf2wF4PkTfO8e/kNjayzyMtcYl/y7kt
ePRwl/iLWmtwaYflHGJYDrqy1AZwzdl8GnNS6+6ZU29GB+1AvNG1M0VmTooY66TE
cDrQu+Mjhqtfvz/S5NBV5WNtZk3+tdeP+uGZ1/r95U8sS6xO0ON3eUyoA4MuTt55
hLSN6kdn/MmVVuXqnOFeHtsnC235X4b5MbAZGqmhPE/tQxsnTh5Q/YiNHqHqHtHi
s+deniTZkG13tzVZ3fH+tHl+44LP2LJnjnk4LEgLl0oO7MM9Q4IFVPqoVj2hPQLl
aHS6UiDwu/E9cOz9ijtlIzdWQl0s3ZfpT63FN5MuVzJXr4v4E57FldoJA2yfAzYk
a9vgrwYi8oNN1rRWpK2QXlCC8rfgLGcomUSlgPnwUiA6IkfJnfH7404lRkFEPYf3
JwbzuV+PjudrAkKvymltmWMyPicAZi16J9hLxiDMkN24cLnkOTGO4JBOL+vk5z8U
hDDf1Cqp+yS87bAs4BaZobg+7EitW+v3o1PuyHc7xjJJ5D+OC/o7+oUKqoyyMuHB
IMrnTRjxbb6elnQ+5X8UT5BN1/UHr4YxQ3YiusJkhrC35mII6M1WZvimeqMdj5bA
eCI+5AVAMsCmsh44YGpXLOsvygszd3K3tobj2GAXwBw7It/OPFMYkGS5YShDEqrA
bvlSmjgeTqVFeBaAFEt9koeZv+VrO8rKFZIoRxKbepeZ8Bdl9W1gPdZ4CMfKIwpw
qVd3L2uXEE7lOuSEzroAoZPdNoKkh/6XPyBLiXx2QxJu3BK4JJild0giTZPpXfKW
XABBmDt2JFH8bxEpgYOtCIuIFlz1y3HBT+K8OxHAAgoaRMTAQAHr9Ax3ycVSIaTU
VkTEcpJQh6DYy78j1GX1Z9lsZFiGijOS3EBwu7KkwMxGzDqkMdRuw/xI5a87QA6r
yhjq4zDD0weZ70gdC5U3WXUfF4xn10cGsaV6I9o9x0FAGVQTf9PJ2twgQQUt5HuY
RANq9p2EG8v6d7wkbhmDkWkjJ5SgNZYKe6u5UBYpJWdo9fdy46evLlRF1rnGP2yy
wc7ZBsqNzUjl7jSlnqVpi+X0CJOBCWySvHZnTNFCybFYx+SW1noLkTRXLovvmx1P
YIo2SQ3YZ/SQJtaaRcn5Wi0wuioNRPbc4mGlTrOod4oBal94mS8fB8xu+5WWm/CB
jF4N9KtFwXWjKN4FbK1dsyk2z+VH2DXDczdhBWgRkZ4kd8t26Y5xgKE2G9cnep5x
GF+d6ij5GM5MNQGbaBi9KH3g9iXn05fIFxftANG2UstoBMCJY9o5t6XekibwwMPp
NtKtxR/kTMK1d/j2xD10PxbFbVtauShPP2cdxtbLxGD1NchCsbk+zRofqQY864Ga
God+JHcr2hovFjDUoFDNh+yAJElti5Bl1E8iFvQUH5c/ilzFeDHLfGKUvB6Xh5BG
IBf/qvABltuKcfC0pJ49/jJRUdxJDrFCkzMqAIgUsn/ijyI4zybG/1d83+eJMk0W
KTo63BKT9az3auabSA/8il/mIYElSQLijETkmQ9e6wMSFREaAHvexIA2PCH58rW/
TnwvvsopIPCEvytQV0NEuXTFYBGknnMf6JoGouosx6aWtcYovw5s51FVL5cByW5z
ZwqVPkhxSMUrQ/TZAkOP7Lf48GnMme5ZL/XBGaMDwCgVD1511VdhHvPsN03UQb2i
6/eAOpdPircHntoxZZfm0fGlv4gOKEDrrN27B1fA3KDYn2OGC4E0GOMWX0PsmMM6
5IP+qA4xqJx0/E59pam+QQFQCpnZMfw1fuv7S0Hykiw21HRLepRfvC0F9hOHRMWs
2OwdCoJ8T1L42aaL/ZUUpWXR/nJozGPrQcovQwJH1AoEF0MXPJ+wFoRlDl92a6MS
PRlH08MboTSojdy+iLGyKizzqljq5iwd0po356/pHm7PDaOFcvC6oF2x3GT1Q0mN
/DwAQQatoTE9A2IigWX7WUGrk83YmFevK3dC0yBSL+xKQSyGbNw1asN/UPoUE85i
psmLuOPsJkSbXB4qxe/4OADMWY/a1A5li514Qb0eV0R0w4O0m6lyiaKPfrvSksMI
XrAGOD1mUEHtUxhKeHQ1lR8L9ZYPI4uzTNGsNGDjxGLgBUVnfcr+DPYP55Fco9CU
a0FY2MK7YAu+R2iVLAEvnM0xMccLzJR+3uCjwyDwmuJB3rFP93jNro3hekTWpWPe
ZsHSvYPacTR8maqQ+hEF2jpVNop59M95g6xWUrYnVavDPHQTgcivEXy56xaEAxHd
TU40Xcmk6FRQgukX8ODPKmPRwtFnUiBpWnZ8dN9WV2fY4MJzlb1RScDR48t/o7cD
qSBKvOrD2FaqdykYC4fh2VWSymisJJhnw5NjCClHNkdY9BZWsSgT/6oRLJjn8Ppe
kVIC/khhxxcBMkz0sMLuqIK+Oze6Kg3TGQU1Zm2ifn7bEXVaJ4f2nGiAjgHWG3Ef
o6bJRb4S/kVEllZVO1fRc+Bu8AMSlKwaAXXXfQOYBP6lHZqtznYij2DGdUqgiPQk
QVot8qW+B5i7wqF4yVetpGliN0vw0mOh/fWX9mdoDmaulATQzQc9/TzoWPQt26sK
/mG5fYytcv8OtM3zjtemTJo+cTHa2jT9oxqQQpxMZXpvEWVxK2FQeo2aPJdB9mmX
HMDaO64tISEvYRdkwUD4jDaNXjswMaPM2Li2rLu7XZKSs7CZpD6N7moh9RsC1uH3
ST7Up5IWHBY/9UqdomU8ghEJJn1blPqcSW8BVxAT/gVk7s34kLgrfpXC4uk3Jpw0
aqsNOPxqigvi4Es33bTmScKCTtpxPQM1pTyyoWlz4jIZaX9LMSHh9cRD7jJ7oUX1
ilwB7rWY4BdRP/iDTpBmgxtbHV/z6nDvouf8ZiL57sapAjMeLg09C2GlI9U65xGO
lZ3FSgxbQ74pb342NMzuKJcycjrvkDkpYZ+8vc205WF3SfJE4Bg6+pg56ZdkiUAo
wujMZVzfHXWXkkpka8CKgtJNzmW5dahr+IagqybGrn7bVbD1NagtxLSG5cdneOnu
sNyQlp+ZDC0j/APAzri60RSVQ5cWFvEHpRWWJxbF3xd9eGywBdr7fCj7hQuFAXWp
JCYg5uURPS9fL1RhQG+dFX58jHcNzcKRdyocN81Ky0bsD7tmVq9We1zFeWQTtrmR
OnXH3wippn6hLAga001B/xN9/B7SROYQrK8NlyQXCIQpwLskXvVGyy14/7w6Hw9a
t9iKr1l4u5dNhvGkQXglyrvW0uKSav92eoKDkfvkpBNQSg7FH7P0RlZdaRuZK6ni
it6vMfWXHRpvVQ0DNIluAOZPfzbcOY3tGDAoZveE8nn7okP4L1h1MrG9YcduvL61
xbfc5PoPmiqsg3dB75A8K/5vk8vDlvr9sexis7imfZZkOq77kafmpQ3UaWbjFi3a
8Twi5x2icyhgGHW81EyZj919LE9w68fi0t8S/q0KshUoa5JIpLXwJ8Eq5UFb9I7+
D1MaA8nG0VbAFqG0uvEFvyYw35oyKuYxH9guxSm6MaCQxrRehkbVAuLGk/ZyCNYg
3rfl6wyMpNTbiANe6ooUoFNCGCizyFIITQTVue28v19L5+V58Mc0wkGwPAFKXJ43
/SP3zw1o8utGpakiQRoEjoEaaZ/WneOvvvhTYAN2KUj+qBYH8u8QFpp/5ub8lpXI
0wOShf5zSM2f7S19W4NGzz8DQ8AssXbTz9db2pWOcICgM2OwIjHqrVAYIIQo9vUy
5N0w0wnsxqJzs5KhANrcyOyzaQPYO/9b3WQAtGKbgOQF8SrIl5A45yd8LLHi6KWa
fnAetAfn8TdRNjLXazIRTbB/peWMOajdLttKOvdsFDE5ciLVd5+i/GMjSrBJR0K7
eiyypzf47VqN4ab8h0jW9/j7OsAkjDx9vSHNHHO2/NJr+JEZyir6ZCciClkGiA4Q
Lm9Em5HkkWJhdkfEfX2Nl+jn8S91DX1bOXI/ahCBywUjEdzzgKhZOQuW/4H9rPuI
ht9WJyHYyiMJSLLi3tlEpXGw+3tuAW2M4Bn2YGDek+8yZY/9Cw4PX2YYKaySRPvr
/YhDAeQSR62le4xEF7RI8ibaE6Tzmh+WPH8fRE8ZkyCD0UkzS7kpnTFveqhKSuTU
VQHFYEPd+SG073FoQFWDfcp/AovPfI7YTi/oUUt9jQz3oj0lNmcioafLyRDMC3UO
Vbx1XJXlzcpxOmfNQIv8AmMgdDzQF2mIkwRTwT5hlCTYjVHd3xrh1jUqq8xwgL6/
aF6n7lDDqPw0+csw5/9B2h9WRrCCcjkUA3yJZ+JxrSQTn7Rq9MznbSg9Sm2PpfAB
vYDUAXaeHjj1b2uoXNObImRffj82TAJSLzxI7vjqZKiSVki6j/Wm1FC+vJ9GNZgw
7ZBD8za4TyBA+AD/nWbpiGzDE9lKpa0bYIlq9lpxhqwCtMDcuEb0QP9bTtUKouV1
Gv7rfPncv6VpPhMf7ecmq9P4/Vw0dhwpzpKPwwu8III6JsFBeRbEF+9eNYn/1go3
ce7hIZed+bWliQKkFKUXRA0mMS9IveCK2tuVMMt4+F2duOW3C5HdmBdCpSK03EDL
GvIY63px/A3X13y9yAhc0jYBGXRObPMKDKqu3WlmAgqQphYNnDDipLmDuIPJwVp6
DNMTOpGu7ygg+QN5fOEWV2d0aUC0nfNnSPL0O1d1k1Nm6SM2GISSXtglonmlkrwL
lRH118Hb2JFZHkUNdbgJoVgPPYvSXrP5G8k3NYGUzq5B6zbN7Cu5NLQuq3nu+Ro+
XcosOA93CJGRTja1aNLdQj1/x4/7/gqZPC/KqV+NiL39gNM2bqcRyG6xgp9+vB/n
ep+cKVj3eshcCAUOQ0gGTM3MGCPs0s+E9eMHXNbWG7cVdcxtFux4rwCA4ItHxQkF
KeZGosFwztQM7Gr1ejjtsTVgCFfWt9MOCmFZe+zFa6jDFGK/O9r+qaDoVd5WT2nV
aBCT9BTHqnY6LcNYZJ6B6NjVaFaT7AWWyg67HpF/RiOEeG2WG/SH/C2MP9DL0jSS
uT+i5cbTQ8eb526+T8zeCXx4BnU3I0CYiUUfpRlT8b68czvaYmqov6ayaPnC+ifa
h+vaqz41xs/rW9uJfuxjgx7BXgP7vOMCRjSYXLaZi41DngGMgxFJ00FMMuzRXXEw
ZDnEVXeC2CG/IOUz4DWfWGowmabFmZabs7yvNCVsYvbIV5rYBHb5dTlXlzo1mJgd
jeuDkrA8usVopWUp/AUdqlllWYNgztbmG5czSrvUq35vPL4aX7+WuS2+aXTM8FWs
oaRSdOcQ567g57PPfyMq2EdjgP+UaV29jgaDQRySgjiSK5iYuo2ZLm4JeLNiA+2J
lIi0AyTJHmxMM5hx00uuZgz68oD4sk+uYAfhH8tNd1D61Tz4EL49ONtjMZlQba9G
XWkYP9M9vw2u4OXOUkhJSTeNgxmBSgHVac4jVQTh+vWnmZauzdTIytBtsRiVQWCb
fVSDXL5c93P/Wk/+0JJNfXlGE0A7uGo4X7Nr7b8YOnLdwtZOhUNBGBSgaZ8Gqfr+
dP7RXCFAXi0oUhRk4utLPp+JQp+r0G7PB8k0Ii1xsZYisHaMYRKMqLYs+cdn0cpk
Y6BlyEXIuSraI3bTo5Q94KzL+3ccvBwYESFkasSHcYaez4R5Az4URd5iMtJ+aZfm
vYVAuutC+dvu16EIBnbc0uI/L3R5qHJ7c8tXfYeBf77xBcqWiNUEy8hT/ROYZw3+
9LxsuXK+15YVVqVvyKsL6O7haCN7UaZXw+8sjuWAtv7l8wyh9BPbEvqrux1LH3kp
lHXSOg/Jxo2gL+UYxPEqrLJTMJdrNrU2UY9oofZQOr/4QBv2k8y4OgzmIVnOZBGV
y4s//O5/ekXYMO4fzYPyFBfi/SNBGIzdwcOJEl7GfFYs+HnaVZtegtq9l/Cw+3xS
6a2XjWP0Fu9aZFxH3GbY9fno6fRGZA9h73q+EiqNiUssmVxCOTMbZ5+HzQkvYqwv
NpQcklH0YLL4s4O7xFMME1z5CY+7E8ScSyMCd+6EdY58iOiBIjn9Affoo6RcHDb4
Y2NeIiBaLoI0SRoToPpgpHGTPCsWb8KiB+5TmoruNKM72BNk3v1Evw9ZVjtECGEZ
Nk1xowqSY2j0jz7cttJQCWow18R5//FTBTb5sEkncEo2vAwdZ5kCAJ+T2NY1f3VA
5v1klvJGUt74GcJHTr4TXv2/o9RIjtUhbJjNrGz2Nbckdn49lo4c+VP/2Sl2qj0B
AFs+swPcFXuJEXQWLc3cgmMCKu0n0x6pazfr18LYmbSdZlFapPqmZCSrsNZIykZv
USioSB9WsOG9gWIP7AvxpG3Xqo3V9MBN+d0asREislsztUz+ze2WrQi5CyL1Atp5
RdJHuO3fbRynzcAY2MJWy2gQYU4yKkrVZQHklkNgdYLh2bHG2ijtldH7vIIM7E/9
Xa4QMvMrYogimDTgrmsYYBIhwLBLW2W4ZXD+KMK5ry9EnRtZ5V8WJSEqskhgLOHv
6IQgrMBOlCP7aBkq00GRm6cor6WCTfZkFWsAsDe8r1hEl6J5Dq/x/ifEEi2bBuJq
FUcW/AMmvZew4TkBQ4Pcs9iU/dv1obZ2puJpJzPwpaiHqdVP5hCz70On67pRxb0l
FD8yosE2gMZt6AJnpQLz8N9iBHOQMrADlGyghZPsBv5LYc5jS8DHAIzcJMcTTCRI
YlWOvE9aLpWdcgOwrG5Oq83miwyH9BPOJL1O1gVlQ02wL1hSkXRMjWvRHzhYjScs
xuoYAxO5AnAi0xLrg+zRq517AeKMx+8DS1nduN+j8xnXobr4uYMNDGpFYY65eb1v
5f6prg/owXX6oGlw5bBM3wfJDN+8RFumFofKXRbAhbqJ4eWKdiiqbThE8JjHMq4d
qUx5ur6JUPF4Xv92yVbXYX2xxYdMhAUDj9Z2NaIaudxsZheMVWtNAt2WICPApzf+
BFiYCKaS8LZ3XAtYQ/JAHR6cSW+0fRCe7Ku9x1VgP4XDQJHwF/zhrAXRUJ6MIQ+c
SRKbIROqCMgAAvFKDAl2fBo/gZB0kmJ26JUSx5PI1lWSnyzzF9aDol65SRrQgKmY
FDWaQf6vtDhKWXaO9Bt5jWTX66eu/YMcUxREScLE9nvUhfKfTo73SOOF/JQ+VWZV
f37pxQVkHRo5IIEOBFBIB2VRRIcT4ziYwEnWnnMZrfODDteEoTomqUdZ9FK+5T7Z
NRzZxCY/IsXFH4RtuM9wcjM0kBtXU8n/lhKG8ZTJUhnBNbnuvBGcoZ7nAAW/zWFQ
RbV0t4D6kq7MvDvH7dOCqovFGBdgNm72GvirIuhBjq0NWXwsqr3aNGhGr3DZ7Ivt
oPVffpZflqoaBlgbXQdrDEJUdsMnk3ggIFVTpZTAn8JhcdBW2l/iYaKZpav/tPAW
dPHgbBo9QzJnZYYV+LQCrI5kQsWKSjW+/lEAPbi1UdZBAVum/W/5LCumXLYShxHs
x72RtTvc8TgXIlUR3nN5YXnfLXg25ff6i87PwierhKmvgR+7mvrS/24lQ9atrf+d
8y1xzs4y2fc40x6NvootIH42oWzHuNdUvmkqSBzS6HqvRjVkjGHmS6YeStmm1y0A
lgEM8nr3WmtbVWvcVkrLIUT94/QMWxnLBXSPfhw1OH/ElIaXdcT/EkLNM99EToGB
GUvXLnl45lApSvW8OkBv0/y6CHWlvatunseSlAcFleK5ylAWJwioNFEgRAA8dmCu
4zmsY4RN0pIEPZJaS1odKG/1AHCWzhfGWjc0d6fd7WYzZHnF87L/h98Fcp7uPWZO
y+xai6nXSvjKfnt4ACneR0dO4Z3dxrSw27VGr6Z8WuXVmf8QPUb6510U3jvK9jBl
ODKh5cx/icLDibVUx0kceB2IoajcI86z6Pflnd03F7heOXgVTH3aZH/rAo57Db/U
EDgR9BdNgsE/bq2xT9YXiNrEEvVdbecND5I0kJhAdcy60hYP12HiCSVXW/QBjlEC
e/BF1PVTp8Z4J/gAb8Xj+HU2VZN2FUBzKIa2UQl81MXEx3mT929bEdAyuF8/qUbD
fpLyt8n3WdMVseMMr9XA//WjVhqEz0Gt9MSZF9XhpuMelwD9ANwp2WvxcLyHJPmk
J0umoE+mtuhxse3DklyRCNot01M8mYoE/ed5lwj0OCKfH2YYwiwBSKWnTZQJysn0
23eKlaoJk1Ny5X8ruHYjn7N+O4LdW5ObbxZ1+H2Ab3nvvqZRmggXPTiySYbw1z41
D8UBLK+lWOltaRzri9DH6nU0PIUDV+I4lGwWCWEGIzKgma3OY3w80kug//kt6yp2
3auoM7fEuiq2Wsp6AO9R0IQNaC/bWep8X/KEPQsNpweZ94J8xi8mIRK+RmpTwEp2
Hfq/sx93erkX3U3rbY3fF6LfS6Efha1Bq7blFgvZ23DxsGLB1Iur9qjpevK7JH52
SMmfIAHsvAQlcjwz88F5S70w2iZsw4/gVmTaFo9MX4LhEUhPnQuS5sTMbXaRMLrT
h3LoZ5PyzB1kLrDvzxYpVKV4dbODCHORJqHXXTxIafKaCL2gIjOE9/kDZgcyF/wu
OHHEWIs7UFH8aMWSTC9UeKt2y0/x5oofJ8yyjbBjStmGBpDNKo9HudFOrstD7IvC
43nIyUBW8oFu3zJaTozrxyixume4k1Sfdw4qVtr0fD7N89aOM6cVP7i2duyJ+bky
OHt557dQMPr4J5IlLPiPoQuvItDk3K4c5AXQvhZzsagZQvTORTfaG0xbEdxRAgAl
LhPvn0WRkCqQZzajVKI8KgJnViZ2n6WZ1oil3KpTtxAssT0yT64UJzEtBT2QtM6k
yDHPlkxM849ifzTjsVkuPPdVfzvm0sQkaynediOdaNL/7ywKf8E4Ct6YnPqTdhVV
03yw+5AKmWmNf/Eseu3dImOc4JdplF4kF+iN4eM8IgNmm5PCmmDYgIJy/+hWG9Aq
UeUjTSaqBwVKiYomJTgVa4/WZADXGOx4ti42STVxhk6OSMm/h9AlajJBUT5X9q6t
7rTUbq5SFYKpukIsjiyyS3liU1fJVcOX0jX8uM8alHLC9y2p03jQSNqR9kzHnQvo
svFstyEslKsyk1hKh7qIjtlHfnlLgscYSsbx9qRO+tDOzm9KZ1ojQFQCB7z/qVnF
S8ghLpporOid8AE6F+5RCsJmqinjoBL6EVawphWRIO7jxPUk9O5RzthojWjdzVh0
JcVWycojTqodO0jhaX+QoLJZhpVEnPlHTrPSxOw1LmVNgAYUO6MPNKfjIsj9xUbx
dZdTp/pgp4vgi2TpDJMs0VwBH+RJMGZtPSrFXK3kgDTYlpruJhoCnDCmkJyedj7O
OMp6xZxt8S3jMCwAxXZxJ0IOD59VylzYsQ3PLkq6QUHj3ntzIFgowsGBk8TuiAzw
LQlnfp37eL70f9yA2goNQXsQVIvw0ZnT2sIYu7TFl7A0ny8ta3MWUXziT1RxK+oP
lA4Fq72vW//GT9frpGsTWaUMBhPuHLbNESLVnOPXfVjU5hqSsTjFdM2eYIzWsSfo
3imPGlFI9yia3LGYL/O5DUOkgkCH22E4exTbocHqv8Ev9eNAqAiPCENiYXKfBz8P
1zDH6x5uRtj5/52+oEE1jkflN4OarQigpiLgOmnCmcbuIT7npW1iPGLGz021/evy
zMidtVveeD5G9tJU1nrLNBhIIdVGrROrmO1IZAv3jaFbRCTyuimal0xta88pfUub
WYh0s9Cp8Esyh1Gu9rdc8zu57K4PUbTLirsfTpw1FUX9yrZx2DowjDZ3LMi7izf+
31OP4mnBtL21EMiChg5wrE+9L6sP2RVZkGTiy+yWxsSVyQi2KH6FlB8g3+Pu+Km2
Erg8uhtKPi7ZCSabyDpeEARGZFy9incWtvAK23k7O+Vi85Sj0tifKUuvysHzyk7k
kL711gsqa+MRCOAGv74kfyrUD73kDzV8dD/o/0/Bxdg4iLcdMCZ+ioBhKSr7SquV
3xr9/Ib/F1oKrsPSiHNzN47ebqWRNz6VhPLFYx2AzRoYEtLq04PYaEhOQ+k5y6pT
PpuA28u05dtdvDRz0oBqcxjFLtnrknv+Km5pfKgzV79fC5d9qlzpWqd3ngHKFtNG
WeKqC0XfWHviPRKcT2n7CrFCELYEfnNYcCTgTNXGfvtMaZ4OKm7vE6YMyRhaxKl/
X4JVvg9uvMViPgkjlOjpk14SbOJ77QeI2Nl7fu8scSYfAwClFNZ2RunK8qcN0Lfq
q6UuFIUj4l4idmhBlFEGbmId02jhCZ2T/+Qf6MiP9aZlhGywJpNQHnVL9NESoH9V
0GSKFBIyztvXko7AM3flLGORfnzqi6GLjXE/eVGOAbyklPhQoR992DBDNJ9zr8ry
07sLQvjD/tMM72lysef1iICrJ8rc3ZWY1GnMBl8VMuQ3Zi0Pp86mED+SA/Y9ZERj
W3jkZARWANOqqrFljLTwu9usNS22WGhRm8KhfBmKuyHsg8fBZayjeUXyDlb/9mEb
tVX7gUdbSwGvw5S9yY9S0N/FbD8lSy1gHEgirtpWcliza2pz272e5gDXj9iP8Boo
HRCZrJkgjPYdxb754g8j7i8ihHoQ07I0jWXNo5YEPQCdnmffx+i9PfkZ6JSsp9Cp
CXdUqxjvhptxL3RaivPbxtlu62YrCUf1NB1YNyAvA20yF4hOB6PgfPMNs+a3xh/y
mFRwh/c9d2LNpYTxqkmg4SSeSHZPukJ3QUawrSjWRm+sW83QtXvs/n5fbvIc1aFk
F7qCUmN8UhCDFNwQl0tNc3emQ4yRBO/gCq99MgslhRVksMoyVL8OpW9+NEJEH/SZ
0pa+YRYQws8h/qkE3xWTlf7psR2Sx/TLTj/mFETA0aJqVnUmqiq86JOD/M9+ebyh
glulf3B/tJJsnLUQ0F6zcWxgt2rkJboPvEW+Odfal8VaSOhbH0mByRwTx6FWUCxu
nOrwAJ37lRvG2XOp7PtlWLv5JmL2+wPon6UJ5Ex8mNaw+TLt5rwUQ1cKAMBfUdSg
B65/vFL2sw/6PYAvdTRBARLjSp9iinoAUnvpB4zMQa4ZiEIEOjsCRdHmXqS9YFpX
6AkD0SfV4WVt0Ha/Rzmadz/nk4w0gHOxSnQoeQWlR1wwboGC/MeGBIQr8/l+UBYd
hylZc7wlKyBVtSXcl7IwxEb+xH0oPwph41nzH98lDZ7uCHgZvH2kx05xADXN76bd
bWNmeZwXOY2/9LNA0c5o1VTA0QSEdm4tnQVP7+TUscV27Uv70JuIHLw5VVnI2Syc
G1EekRYgN7EAM4x7ozh8q1TwGfUbn+VW4B3A9jeycfhFmlEGuVIFYUsJmdKXJ1M4
7QweeXRCgb7LNe4ojNrrDbgt/hryIOyZXwkoY0Myn1hTCCkaDs+32wc7uaNXRtZ1
KXbtPXMLc4ZDrc2zt3LANHS3aZP4FiXzBHuahzr+qIDv434yc2RGAafeviAnlTmf
07lKQMCY0XnXTgE/663rvGRJ88bwhWnb3HSZLpVuu2zGf2l54YBNqLgV0iaG6at8
oHpWfRWhLjAeBMzd19gp9wehRRqAzNOMVbovSnImyEaJFsQRcA06//ebxTH71/9X
Dy/FVLrAJvbonc5VjdgqIuDJ5yo7/CJ7GVb4bByb/YAbOyMPNOR5SvU7dCSZ6OYF
CN1tG2+NgxZfbEKk9jMX3gkgm1ADstz6zR9CPJ4IC8M6X914xSU/QkGWnEbu5dU2
z3ZjIniwv31Le4J0zeECxDiC3sf1R0d3N1OffoedSonT6Dh3fCuZ132r85QK0oUb
oVFSDlF3EQx+ap9APXFMRoYqkOrJXhwRJEWL2qosAutZpllDrZ83VSwuwuEMkO8l
pk6iXiZ+rYJfEdU8mSfG82q9HaPHUoZoXOY1OhWaE/iTIa5DEyqFd8tzbaxg42W/
esTF4oBCxeM6tL8unJ0ErzM82BKJh+VtDwEa+e9LHvlwtQe8ndeh3h4Kbj+Oy/BP
JkwH9Azi29unBURiSLJU2h7U7g2YcVwNq2M3qQWJ0VO0QkUj6MuAFUT0mTdKpJWf
K0H91HhhQmLoQPBkkbfrwlu1tj/K2HJcIk7qXj+yJeZuIW8plq7EnzACC2cH6qZl
Hw87ZLVWHb4zWj8c3aNdySROZGV7riJlNme0e5ndH3rJqW7B8/H1mOmCbDjp9XXE
Uop8QcG2W5yeYDuGEjXsY8ghcFRk48kF+kt+MaHNtBDX2BnFQxJzF59ycd2digX9
bAJTcbrpYbxsO1fPdazmxb1zDuWnh7rBI8OHAqLqP3pq5bPEAC5ILTfiOEM38y/H
mnS2Jmkqh2ovAkdTc8EqT02NkDpt6M2UJzcDioLscDYNwQ+vykgh8I68Df09i8PA
JRcXZZ3PAdf6+ia/syvVinLe6lNYn5J1mesyVsnJQSduLvBdOFA4nQtIS1PUg+Mt
9dcSPKXQy2l1uowjjxkjTt/xZZnxcHiK85oke7NbTjAfu+BxDrtVxEp4G7l9BAcf
Dyuz2FOKHcj7OOE/2Mzk7F4LtxR9W3UNAVA6Qr+pT7caO/SzwKOkW/9eoujkLjH9
dr9nmi5bNnrDqsUfdIdNFKfvuT5XHDjj2yGw3pWMYzE=
`pragma protect end_protected
