`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lfd1mP48LYsN8InkMCZKbiXS+a9xrc/z4HO0zWe5ebOimRuG20aGeLNVcFfMuJrD
m2egt2d+BjS7vop2zs2bRBv+lfC7XRGf7ixd0ez24XQipv+zer3OoAtJi14eHnwb
hVi1aLsiNvEba68RlMZ4oStQ6E5lXuDHE3R48BQ23Zc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15584)
oiBc4tsnTkk8OnGHNW1lhZIjVmfPMxAsv0iPJnABrqmgeg1QPNvbamnoZEH0MJEM
L/PIFNAtQPTLjvIiFuw4cYixt4NkHnX3s5Gp16s/XBMpnyKDlmVG/gmXqzTEpDMf
NDKHyJJMick+9sZZLKCAirf/y5bda1qeWSXEkCk1JsZ7c4YqbnSZIB+loNfiGynP
e1wVhw9+s2VI1dLYBF4jF4xU7gAPsH5kqFom5Zmy+bpiTMPNZkCPJLOmqIPlKekZ
RUMZQn/pm63ZRZjxmSKiKtArFfwucQxfe5JcssFzcrff1kfMidoM95F4yOBYVR4N
heyT8H0oHXnMPGLhwbM8ls6EUva7wOQCWyHIX5X7UvIxiOXBD2Yjd0rAdEttQD+M
TB/ccl46gKJ49LzFkKSAcJsbX3fBE75e5bs12l1dbSJtobTRYvSZ3/XRCht+TL48
ak45CcKkmJcUKqcF2nKi0WiMnugY1wqy/Uv4X6vQQ2xXgzUJxpLmJIptRlsDJCaS
5ch29qiTcVaQzryGaKD9O7bxGu1E13wTw9LmxNjQLbF1wtRvjP/6KV2H9ksECXUL
ukpW1c8ZArRKu6qjJ4pBuV5ssG99DQTznRNmRlsHp28UrjVtrx082Gn8HUy5O2Wk
ystL3ZFm3qOaXXl92eMHKLfNJRvSNqut9MupjeWf5SqvF1ZigDJHzYl07DFg3ZtH
IN0l4juw3jplNbTNXr7HrbTnwmo7lSjgwlHR+m4TukRoom4UkBPbzaOZixhB26L6
hU/bHAkRwdGfxOUwTktG3iQvPVA3NknlnCzgK2Wk4JGMtrw5gTx0lpcmuMsI304h
E6CZ1FsbDGRAiKp4eVEwdoAKitEZV/Ct4YS+P5JBH5hUuRPq54WUkh6l5Bnt0a04
0wIiMdUBlXHAMCugv21DG3aK0dX6l9rEaG6zhFE77H80o5tTZozPoR04mVLecZfl
/jHlQZlgtiDCOOVO8GP4wzQ5S5VGfbnkNtc2xKswlBb4N/Hjx5iF+GEtryplYPzh
EdnTD9YR96GCaorMOdr51QC+iSUlSCVJ7/UylGUdhY2hrk0MINWatE8vr01WR7JC
JWeU/y0I9lVATLJDbQe1Lu6b4u6p5kcLRiiqzi8dJzr43GWM1YWUplrCtMRU3iDM
9zH90UtDK70+lEMEquuzVodP8ReFsrYbgKv+MO44ZFViUaqTx0qgIxlNak1Xu/Tj
96WyO6fmyWY9YBNFCxoYr8ZXQ9lOoo/2xsf/4LgmvOPeVsYoZH8GpKQcXm80Jplm
uDkT2WMgYyINhyOyE34MRNGhNKIt4tpOT8Kq4VAP3ZEMcyvfUUXncH8Jej6k3SwR
EXFAG5BM9roKA3wgegZBdW5oLs2X0g6hG1RJGBhFkKzVf3V5bGr95P0Xli3cVUod
RdQmdRWdSTh6c7LFsTD7ABT5qv2xS3l/bL+eYkjmksndHe7bpu+QXfoVBfXrXu4J
HFpFyQM9lU3wcCMRV0/6FU6WPqU6TzmGob/eU9lykfb7lkjG0tv9KSfLuxvmi3vO
gfiEBDHpqylx/zjvi0zTGojOcc87rSonEG3+KM3wAmtQxMQQ4HjT4fRogVt1QY5k
5+WKrgls9tfXU8gcZQ2Q2m/SVtRwWDKxlG9AyOB/d7WQ6wC+ax7C1v5UzaIvY/V7
GIZD+hkdOSm1O/lf7kEiU/lLwo+RdRFeAvWbd2NyjEXrREZfPB7DX+Y9cYHxiHda
WjGvQUWn/dcNfLX0ic7A0kyciUMpD1jCTE+GCP5r+aSJHxngda0exNkYTBOD6tLD
G5lorDL9uwZCBFp3XY4VL8JlqNVrcsorFbfQgU2kQGQnWFAkVFAQBq+bDtvnFJl3
82jyU4cox6XxYlYSy6OGtGnUl2UMe8EqkB4vM7iOm+MUKG3UP83RgJrU9pcZeh4x
R/lSzAhIXItNbj5LYguqOjkjrFA9lj8OixyegiE1OIiae9Uzmzn2KBN/BWtR3g+w
1e6WBexbnisJuzfcXakeR4GiNIkmSsSfhqMfbeFGJ8f242Gk0SDpgSfaN4UkT5aC
1ynS0IMZFPvTh4j9+puTL9sFq+OkU0Df/Vmd3LVFdo+VaolmyrXf0FckyyzNLtvw
NFllFJznGyRYCJwMYHe6X9aOjYE2QXcO28BBewqSPJP9ulqvNYxEy8s7N2ruzdcy
I2Jq4RrX/Vc3pJxabhwfuZXRp6OCbjuJNjY9f9xT1+Ud6karzSarlNv4NrUbVlGT
ibU7da9JL1udI6GWeJPuB89MCYEsHFO7lwg03xadEp0sfvN6rEpVZxuzU+jsfHnI
gXxseMT9Lkz2IPXXFefDP3beyh4tJpE93V7Vd4Zq/zq7R7p2IaGjI1ar2fCZ4s/G
w1BOVMoUAOuQwP6GtulUUTjlmKaSKwshJGDoF5BbAOFQgDIrSYumzFipYStWkO7R
+dDelTA7Lho4xFMe+OEqfjQQSrYlAYKeRufbDC84t31CGwnGPrRaMaANpD+d9U7z
J/hmGq+1Vbm+hQEwmobNDRaazdFJ9N6IlJDJiS47giCnjnuFYaDgU7EJIg4GLRZy
IzKy/NXlR4TqlTI6FltTFHcvOWYbkd1igv7VlR129aa9OXeJvWmCQv27N0tyRMKF
+2jNFz3ikXagw4uEyhsorHDp0x2ZoA4fqt+Bu56Bl2wzlKiAYj2jZnmNJ8FLR+23
1zgEvcKvGT8H6LFJmynscl40kGDTHcjcugd+0FzYpdnggGuGRi0slcYVTwgOqD9F
wPl2Dgmz2Q9k3ocx8QqB6HZQWlpdtMwl/BmP7pdaS4FKAsIrKKwC38MB47Tas/lI
Bpiid9LDuk16/oREgkxWSmI4wdlo8sTDbOPMfkAjpv9ZdFM4CncPp/qtLyaI1Ot5
XcgJ4ZmX5J61cr4BSNkNnN8f3mr/0qG6rvj+9Ork2u35rIbYMVVouzIfzgFzyjOT
bUfttFfvk9cF0WMYwQY9vUQhND72CiaH1aBAKrtFnz25NhM0fy1lpOOhgxten8YY
IdkcMbeA92fBP1rezD7Zq17T/zgvTtrZlU3IipJrP3wlzoJ1EyKt+UqYEeNDuqfo
8VrgvSIndIvKSHc/AuiB/S0QAFak/Khz1S5t8qDrnQ+rcUx7fR1oTocfkXVDUHk/
PibKRhQt4mhbkw4yiSuNTcEpUpjQYpeWKUEmmHVXKZRGSa5hj44tu+8+DmR9voPM
Zaho+nRR7XCVKTkAHK8YnPfa4QBJ8AZ15tnRZNHPgxfAa/GwBFzx4eOzB/qN5foN
yUIsivOyEqKDncTdZhyUoRgTES5tt6gKqTksqF/0fAgxshKrWx/OX28s6yrZ9hRf
VCuP1OwVGScccdUnECXneAkgJqnCmAgFWhrYAQ0qw69I8izxCW6CYvYfxuAvIuD8
BD2rNig9HS5RJfAMWhabLuTuC7AVvi39lz0jrn9TNRMiA96AryH2xwtdFB5Hs/d7
fHS32qWkIv+jvpCdsPWtn6n1Cyvf4tbh7FRiwSkMgKeuaIaQPHneItij5RVvRPBz
vYHr0F/kn1JJyJjSztBQONAWZqFdzSxyIw3/Yp688mFtS93vZN7l3pQpYC0hKWMH
AXBazs9ZqIUfCLIoqkf4L4BSgoffjPoRn9F5rGh3I4HH/LsCO//q2vg+TDrQEcgc
dFthzyiloGza0Lw5jx1Z9VK6LFDPQ2ENt3dv1QyENxPuKAucM7xfqmI02sYHnaAQ
W2wk2XtlCPsAeitsFsWVb9eY3mQsuzLi2YLizOlZzfyUzdcPfYnICekpIv2/dxYC
BWBR4kEJ4L4dBgu+8c62v03ecGbl4FKc0uPOVCTdKz0M5/wLCUo6Jad8Aa7wP+/m
2bgOtds+eRGq2tqVuVduXUMPC7264t9WqD0BI39+o5YXAG7CvwREs+fQ67j7/sa5
m/TuZ4kdJPFgT3MBW44IgfTV+7bjoyBAN17gU69jxqJsu9+7/QzFOFQREwoGmzFm
CgZZZlEN53MNn2gV1Nb9czgdCEZrzGreF7cQjpTW9hFoLACmvvmLEKJ95ls15x4q
SeIdnHICeGRDvzZ4DtYXQ/alW239+5w5jIE0D48zVBNAb1fFoF4aKxuaLN1MwPNu
707xY6pfxxA+ulU7xOSuyMGoNMqL9LSc/NJ2KqSRNm2kG2oang4t6aBmxLh2n3mS
zvp7w/FIbNS8rZPwIL2cipoY/OZbmIsuZ7HWuhrKVQhuy922sW2vgcB9cvdaYKLf
pgm373AOR7+kQIrfCz3BrZT3VfUZT9SKkJXOGljO8G2ue+tlSp5y2mpXhW81pBmz
r+7EZ7v2++QBZRcznQC0grDMKd+bldTFISRZkOQAAoVz9+gYugVJfX41rFn1fJv8
7wq/KSW8l3V6ry4ZcJed/eqXKROYqRfOZ1inswz8u0IcWZzvcFTR0S3Imp1loLwK
/iGMJ8o6oDlBFPTIqzH+TqeX45HZIAKUw+5jVtpJj4t9zqfx4o4dAh1nAufAmfxc
TyKbjdqeyQ9Fjm7udt5c0wBmE/TE8T1tX5qyw/zxqJoRtstvOeGCQhAVn6NakIVd
Y7o8gY8q3fd9Lwqckts/D1Cma+bobeVIE0XdS1RyDNq2xk8nKsHFJnU1yXOJ/KiL
c9Th2ObSE/liPfythxoHilPpQ9EaFyNbv69yDaLIHauT8rkQRr5vXCag88JN29rG
OdMXfh06WmDatVLhABbXrZ0dviaBMzVBq7c/JgSkQRvEfWfkQapkq48JqW0i3M7p
2/rgpPc/NsyIK04JnxAYWidbs7d94wnp0YTqti4purxkAIVCHidrwQV88xgFuRt1
CLdgo+RQ2cLqjqd7e/rp4m+AvRoxA2faZlxihS2IgXH+nA9brBCqoBbgs8cz7VOn
bMRtZsX2OaJp5R7O3Y5KKcBb7L2KFm2yaeXoifyKypku7z/8YIqZS3EOV2oMa3zY
H2KyZk5cVRjqIA1htJLHxChFQPV+oBt8g5cHxErV2jVi4AjQmLeKEluWDxgD5/ld
d4rlNr807Jh9ZVWahBFbXNDYPIOrwq67Z9qTKu1v5fdK6YIdSdoGttsHvkF5MABT
7gZ+cteBik/RP/z5qQS6Y+usUjHflRNC2FpVQEb0T2VJWJsKI0cFgmEyiIeNnX4x
hf8qXBZHxthEX6eDEmY138iCSbOC7vAr0OFDFUWf9TaGs0zyYZcs1SB4/i3HVD3w
XQTaVo15hiCPHNOQiayYstZTc2PKIg7655HZxsCmJNzbsLNaC1EO//TdcvczR/8v
NeYrnTCwOQoY6ZoXaClPOIBUwjkO/cKiAgv5wQlb8636c1x/OZudoTbJ4yE2NsO9
5533Ua2o/lv4P1ybj5BoB8GM/oa94CfrK4DFx7n+e8qHt6r8IMiTwzEyztEGLoQ1
BCaARrmuSsaILL1GBE0J8MF/2ou1kWhWDqhSuUFoUqbqZxMXsyhliOV2QjD2ASk+
g36YVEpco1/jOH0GblUEhqdEaOihkmO5WxogjaswocmecezVLYxgrF+M4i+KzD+R
4NQ5JMlHu8+KU1WYHb9mY+FPla/0v3MaABxO2ycNoWcKkwWHRelaiZiqVuOQeR1O
qt/vy2j1jKYOgK80sUYlhNsxKGftcMA1rKNYC8qTUUl1ftSbCgEwmGzw1cwSCqtA
RnjsVyo/sxRXJNk7iE3idYc/sHqvitKvd8ZRpmYTI10pj7643hvQC3Lfh1C4cIkC
Gyn3tJOuVI60+7c/Ri0AaBh+OKwxVYy/5FiQyT4JMz4ctdCKYBGsTgECTAV9dlU4
jkRE5e3rrOZFoK1WJa9oyyg16Penr2HG9RMqkL1bzx5RSGAo6Rxqstdw4KtZOc4E
BNelPPJMruEfvoTE0ArdrWdtCKocWYqOC+L2wUgQ45aLPj23qPG12gIPyqi+7iIQ
8qVRv3LgMLFHPFE+SAdqsgvd8mwaJEKSavOqarrMEzwbK75/ZVaVfdkE0ZJCz3Ia
OhWPDwRVd+mOOsc+IVBu/e9pLzJw5GhJF+A95LFdkDFa1O5dp8f1mOGYgbLsz9nn
fM0LdKOElRqLSRpSKqbPM+IdhgVPN3BIvO5kGqACaUnPrQsVKeO2YkOrK6JCX0Lq
Dua6ItBLy7hg7HPS4iDBeAwIURUpiMNASaQTN21rAvjYmdnUdhstDeULNy5LPSiH
jP8E+SV1VtojqRNdcVD6XzkaqAmnTgVenW9usyvOqm9Xa7UXXAm1yfkRajmNxBHy
GngUwA5m1eEgBzl9UOLrKhc6i9MQkJtA9O7in7zBqsQsDPHw7hrKkBOvFCYgMpiA
GApmRwIlnSXFKd2wEO91t9+PJw8E2nqlLHfg0C1fAIzVDevecfdZfjKsVXHYUIZO
HVX90Zxag08rEbarRjycD0PXC50u7Jfic56IlBI0DqLigGMos9YKUphKHUl6yuTS
Jz6Kd89Hk3Z4zzqZnvQMylm7TMuXZdZ/yVpXYjRFntyifvfdaWj+CvNvk4awqJBo
sckzrn84SwOhqNws5UGU8C62Rz7i1QWSZd2DIkNsZw0kI9LOeDcFG02tFqtmArGX
Y0yVnhtYoM+/jcCzjVy7KAxoOUbGNfX8NlvVtgp/cvBsV2RHm8avnv7JTPtThHiJ
tFiwlQV30uLjRrBUsizjKA+sLsH3spgyNDkGq5B1SZjGS133v2yqmQfxPKRtasnf
AZdp7MlIT37cT4CHbJaBI6kePpivGLSIXWJtKv+QgItHBkW7CGfPt8J7tpU7sSnT
WZJkHDG8vNyd7RmYwphrkYVlyLPaAn/qPIgASoix4cJ6h6YUoncClpDUSp7epsB6
bJOfOjdyP3QALYinStLaYqL8RAAyI6eA4pSZ1hks+SVRYJESwFxjllpsrp1UqWY6
vqyeOYAxIGBOxZyp2whLxFZwHQ7vqa8muMB/fN25VePt7+W4WTsejsXPPhMNEPg9
m9741HLj5LXjWHbLotPD6+4S1gnBhDGBv7Im99e6LLK+X0hmOxTqbs40oAnsQHJ5
GAbw4wSs86FkO/txzOE6WWeSDMuDSfYQCwYIivLoVR3VumUsxDBnUTo+abSa0PPh
aKS5xF/6iTNmX3kLrudtEOXcKSYQkdA+3UhD9BzNcfbC06vFyWTUEOqoA6EDYuhY
EZbF7cN3lL48xdbFiJ1LGwUUIgx8Fkk9HnjnAGWK99SPAI3eahpv2kiVGoiENlGr
TdD8hxKzKa68Q2KQqc1/4mbxFdb6zwcBbE4hCACkbbZ+50+98hcDsC5Evl2QwO7q
nCLD94NXwABhnFwybEFa//50IMUC/12AYToUOzRgdJ+KdFjxRN1Z3fXdNpZzVGw2
IzcxRs43X2XkGIrhXt7oZKQvkQvPxIX27ltube3mCXWRWykik/lEttAO3bwJhr54
TctkuqpYh07D4AsXWH8G2y5hQ4KQmb2qWHT4pMJvapo1Y+2bIrRFPwvvUYDRN/oG
kWOgjnUtBlGCJqXdYz+0osHEDY4b1+hw7CpeFMnHaga+4dmY20qnlnROh7FY7ytW
4UsuWWNwW99McRrwoonhIzgxwNIt9S8IZ1PNLKWeVGFVic+DamN4CB4XAG14des2
bzX3lrxBtqfNMvS7NL22eic28EozKzvDpEKqKfD0+ua/OQIBKFzsM37zdwY5dH1t
SgaI2OpcPNaqB3w6Z/gUF38sM6AiWDO4Dm/nhyVVRwcu+Or6s2cMgB0u9WKkQHV0
8kMix5Mb7JTye+kneeyC94vpGZCAJfpT/ypUgNuu+IZ7JxtQX9fy2Qto3xFvV7c2
Qxc4yLedwUobG1ZNuOLJPwae8mdhkA3IaTXVbQGdwiqKfbi6BjRtXLdVNeJsMi4i
aMVNNMZZyB9ESvD6C3c1gDhsJY9pUBv6AYcJtoyJy86A+eR5X27Wqoem5OHZ/bY/
24uJF3E6XSlk35wgMJHDaWr5CKrD/7/f9CNNcbApcIEX7UPska0eVPiI0H8lzt0f
KXXXZ29PwydegrnJc06vehrm6h0efflIcyhAEbWAu3KzpxnjW5n/owQ+8o0NX0kd
nSoL5DjGmqKwScckmgHq7wtWbkOmh90XsgfNc+37zDHmz1aLfexDDf8P2b9BEg/T
YmCfXzYLE7+AJ4dD0v1IEDag2pOLwVFhTgBKN61Nfnliqr2ntRAk42nKColbYsEn
Pcew7Qbk9/qq0sUVB/qf9syE2inDoTsYzExqrLr9V5G6Q2XkdtOJTlV7l3pAFpY6
Ut1mYXD/ZIgCn09pk78hFc8/ZyBspBzD5+SMOsD0tQWxEXOZs43fNPNgmja/OwF2
dUf/Jnr6Ii2iz0tPz2xiDlOW5SbcHZkmPBlYf9QpX4LlQ/k1oGvgyFxhDxjj8GfM
QSiT8rDYjWihiAen/6P4BEIJjhvl6uoM8txjgOJ8aj90lElf7KWq9JFRG9avRJlj
HuyFffDsDHekxPAPu0lrXu/GQ/X9ljgchos4j1CET6xO12HGf1euIImkAVOU15zr
V9armPa8YAUKXqP/nICni/ESsfu0Eph0vjASPPLKkirYNRW4ZVigOdOBPD96cyZi
r34nphF7n0CDwlbRQyzAaGjSixgp3RIe0f2G6pQfMLTKsOsf35VTsFLC84vIT8H3
S4T7iCiVORm3a0nUytdyXAC8w1m9cm3ShfFCymJEMhIk/c6aXzu2wGrJZyizA33T
y+M7GSfcHf4EVj2yWIjcwiOZqcF7cymdMDdWe4nxJUjra5wXhN66I0RDuLNf4hNJ
MfM5llshHHFq3K0+EvsnngNZltZ27HYZLezKwhGtobwZqeq07V1HL0fTqou/Sc//
UQRxyY3VXydnnxgnMw757X7Kug/+8GARE7kehVqgh7VJdBItLtddI1goyJ5ZM35a
AOUaMT9QVNpY6RPdfG8fudcdOcSrnRds6xSb/AWeAvjzd8FFt4NRCLXYVg5mIfRC
ggjREwtRk4OUEJVvvQawXopm3vCV9cD5wuLExxrM7RimrhXTJoDc6MmFiTSaqA01
CtAmrmoYKSiCNEr7ldUKNTvzjPFshMUaGOERF30VOL8tSNIS2Ft30uO5ZVVIieuW
VY0nvO+9sWnyg60mle9kTxeoxLUSgqqV/GJ7th9Sp0AdSEVrkElddc5IUKzDIr2J
bfvpcUUhZhCqT6g0+6CgX7UK58ci/Ceyv3UJjIJhk3NssW0dGLr9Vqtwfz9NjRsG
6EmiZ59KauBAheIBj0bA5GigTTWxzKIr+P6K7dc3WNMzuQfnBqsvlEJ0GRrryxxn
21cVZb9U0E8Xraaq3WbBYAfnPRTEHN6/pfvU2g9pZE5sqqEOiCn9EMfoPU8MYI1H
bMzqhdP2VDjflf1uOa10eoo2ryB3Q+P59dnZ6eL7uMtjqk3rCrAjVi8+xPML2AzV
5BNZWbxqIqzjwopVyS2i4fzGAm4aAMRzl6Te1vNjdz5IHu3CrBOq8FmktTg8Qn6j
MD4N0DaOApijb1NuiY5RT2TOo16i0X9MTYOOy1gwE9bcppQ12Q5UC5jqFy+EUAHC
qHfMxi6goQckcFZJ6RW2EyMOCugrs9he8Alm4ibWi21uOKVY50fXef9Q117omVwi
ggBe8TILZM1gm37x5Lo+6RGCs/bgxNcROtwv9QvMAU3X3OX/DArt8PWTfTbFfaaJ
b79qPdYg4Q9fg+LGtvJNMEAuFLBLGTcUA01GHAzt74Yyic+Ik1IjEAn31vPhbv8R
ufVFfDCy/zwSkIzbpE5w2pLw89bfci03WA1b5x0V0bp6NZEdyU4remC88h6nb2O+
iYGtl9yitCutWufcyUDxPH5nQri9GEOlftprMa4vk3g4+3rc2fN6JaU3xS6iG+bK
id4c4OJcd17SHoMOS7EZIlb9V3BuESUwS4yKLIcm7LHHLxI/5ogIj0MwAsXoykWv
raiZvO2FJe/QXxjn8pZ6OlSk1hX9mun1Ur+0IPjaSXNw/xqczrwJw0zFSLpKzyKi
nX/53MTaCc+KW11QqERMbtdENKKwxGJJPr5PCBWYFV8Yubca3HftbQjw7klXgrCq
Bk+1UMR+Rmd3FPLWQLSb5jeqWaJPiSL3amHZ4pqtlq8BvN1BSXfF6ruWGc+AigPO
/sd7Xal7C5icKcQ8LzyGWKrEDhkIs5KaP502J828QJ92YDZMISoG1k5Kj+GEpM4u
3imLK9XxK58icf7Y9BBXazZmeuK9dTvdzdtLQib/haylghPN338eKVRVsn/XQ0Av
/BSmTSFmjrxBLyYg1A9h45vcEVqBhkAX3KcnM2D7n/rmGyG1FrijOkckfgomNcK0
7NOVJomsPHDMeRP5aoncGyx2GSsqDFoFmsFEY8I9S38gax4ski8i4JYMw53supw+
0Mim5w8mre2CaJeXDS1qWy4jha23PdYSwbQO6NFBZzpUFFIHYX3LvhimwZigCd/w
PU+7ktsDudMhX1GshZa/BB94OgplkydZB1oLibQNC6+yHnLL63KlX9nIyxvFSO9U
xttL5yqf+sNOmktaoOGLohCAPTaoYD2iOh+dBQAEGiw85YTey0aMkTM4H1EZfQ65
djea8A5/jDN2HP9Ru5wcQDKdCU4e8gNVGe5OTrc6RFBgwcGQMY3yYYGAHoBTFtf2
aXIBmZ8FDLaWsOpfEDwvdKawbRYzw9HC0O8BUV6bnup2pyTjX+gE/w9OYFFepOSk
ee6AflWvaxuakju7VmKvFO2a80Zif6Fj6+NFaYN+87cshGJqhwhTiQpev6qX1QFP
wK+TM/wsHyTUt4pW/1xcvu/4cqrVM6uKdHl/CoC5YngQcj6gXAzGhcjc4A+3Q0hz
i9EYc6dekKvt0RNyun4ni2fuG7zWsiGjOs8/QYVdjZVZ3+cvlmftWL9sTtIWitMe
oz80BVua/WJ9GrKSoXJA4q5gTAKIl3BftcfJvpnFz8CoxHDCCajtAtDR4JHb307z
9kericF0/9imj+YuJDXUdKw/A0PzpVdYH5ejJn0IVI3f3iuLqeKMHmA7ANQSX0V5
4Lg5IIUXtEXMtLBMN9zmyTEXAPcg1b1n47Cpkp6+/EItLCx1JLHeRveBPwX68hrr
+sdiG9Gs3ARD1itfKUQkEP5KIBmK2G35dH83e6EPFuYl0VeuAHT8tqXWGx2vOGHk
yy/1eWXYrLyOELzoK5SUhm8LitWYpyUU9XKbsF+bJLg59/NvLkcmS1vjw7wF2PFM
D16D0vR86BkcfkYPulP8UOYeNAUwO//iWh0i6upJr/R2dBDULrlqu7AtsulENQ/w
Q2/r64A/1Pj09mgbarod83Ae1zxt9yYPkvtmCsTFzbeh8tBlg5m09zyfWsCE1qiJ
ygvl+3cT6HYW7rXi9K+HH8VSlp6cXCZiLUfU0NTMGHj1YKbiAX59P+HULq+Sajz3
FGniq8Q4uXaLPoGMftSWm02z51f/RpJoyEjobzsTFbN9AQhQAL3IEFYonhNU0ok/
D/m4GVGKXWzqZvShD/W8RcnjlFAYwhDlIfVbIre42ZgsvPLeiQKxDfcM3+HxbYIW
2JdhDxNbO7gcHiZgE8lenTn1ddFvON1i0F2/1dFvgQjWy7G1bWY6u3g1AJNYc/OJ
xZrlhdlFQLVONbvIR0fLPgwpGVZYfh3vuXA9ssna0LG36hpuOwOXeWgDFoYuf75L
OpAP8FysSTjrFG3SgH0G7CbaSHsQGoHzdad/ENM3gDcpkdlD4gSvdIXKvv7tfk4C
de/zDxfHODkGPMGGHPExhkiZCB3k7Izdgowvjy/wM8xQ1C6858BH1hhoFQNZB/Pr
N75AVskUhMyRojr4s/Od7dDd2kttIR0u3s+VZsv7YFyoJktHPXajsNDFLRp9EBZB
XLTExFZq5noscm/tvgIl+20Xx626pLpGLKg6AQgGkNGpuQfwJxM1f936FCIxZ3vZ
AUJmNfBSvfDCU44kik0lkfVWAu8Z5vn+kXV/CnSFs033cL7qr6JvmZ9OpFE3kmnB
MbSa1CAdYeVzOUAv5hmah7Ty6XcgR17UK600e8Fa7+oJOJTvF/9OONHcj4z+iFCR
InquwEHYy9C7lrqRQpfCg7f601DHARneSBjml1JR3HkChtx6LjNlAvBrotYj95wJ
mR7SM1VWEU+gkHZ92t2JWd6tWu8kWWHJiaLOZdkcmjUc1htU+w0Cl3xW2HlcrpfH
Nna1I/RXI5uT51dkzYtwpZlsHZ2qE7b/ji+CHiH5UO46njZEsLJWNaL/v5C9QDAd
B7sBzpE+JZlwPwGvjsrTNCKDuoL2mDB2tq4ypv3fKKtIm8aDKhf50m2uYu2ESPbi
Xodc4+4dVjBF2RHkBUhHST8QPsP+pSThTo0/E4h3ZuFH71CIv5G4uSj9XtVLJKC+
U+ufO+wPG14StF6qvODHU3YBNIjNv68WwgArTMr0IIf0KJeqckwwGnfA0vQ4Hzqg
NRQ7E/jUHM6/Avu65xFEYB1Ii87rAoOHbXULyx1ZKKN0FfPg5GGnx71dhUeZ3B+I
WPQ+irJOnI4vJ0Wv5stW8lJ3tbN+8BjPPgCHqnnQbmelYLcq8FNj6TFeKCBfzSFx
5Hi3tUSAtn5O/+gQquEdVeDIv096FKp1vLnEzBS+FJ6UOfKFj8jEjL6qaryLadW2
c00sNCSuuAdy2cyW+YOGOHzmcv2Uv66i9ds3ByDJklWruLuAJjgl07a8yNDXDMF+
wz7FuH/DLpPND+kfFMla3k22MEnc6ZtFH3/VdKKuYC6306ATnoGCa8C5OnOIFkHi
IPATgv4AS0O9jFsrLvxQ80V/uBIUGlXBvll/OTJduPTRTypVtvMCD8x/fzeeGsny
wJVCPxtLK1vJy41n4vnsH+kjpz6DyjeWaJpKCxkxEt8aDVvbCHEL1cC6GICtQn9Y
OKPzMyuusyXOb48mju3ikPuVy2NJVGjNMm5C0DNg+kuwNiCpK28FP4FAxz0y24SY
Gd/7sMwA93c8pRcpw7GpxzBmUbmyBpBy1EejHBX6qAEZEf0qUBYRfOx0bDehDD5P
yfM9MgBXWFcVtNmepZ7/WK37CHvnBd+kPkL8Fos8bfRtqjBXvQU/xZuEYfSJOYsw
g5hvoEaiNNsuke1GsvPYnlhlZ72ypvwuGAwZOxEFTDLJDVALkCg5MEqJTDncQGMd
ROYBBvNLfpDVz4d2cLqScXuLiAcOudSnaLwh6mZlpXFNl6kW1EShUdwTkV0abnpg
u4aJWEzyBF8cxBO+lpObAtaUp1ICZ1F3Oi/0jeLca2c06FoSDj+ixJRugJRgGFVg
+ZUlIEBjUAd0aHSDbqAsZ50vonk0KYSmYvTrO9LQlWoRQR0ikQuD4oLUg0Y6KWeP
AjMp7Oy8likxYmaC6GAzeCLg4x/HYutJSMlqS+Adlt/AvicfEfWaZTADhA7Ep7sG
xBbDU/CEBRo7mEydC5GLOkKRhE5d8oh39CoJ/cWgkLVcu9WXQVW2voPPSf7KSwjl
jUZ3NX7Vo9pQkYUIO+6askuw//dvBwN2S4XY4/vAYdXc1IYL7PGxJr3/KUTsEYML
dQBqScLrATqQfvUzP0bzhGf7Z6/TU6LEpo6pIGn5ualQO850MllR+KQkS5z9tDsB
8Un+MRcDA4SFiwxJ3OuekgyrQc+dOERnZeQ/M8OGyfbMPP/r2eFrDlH8yaF4EYcW
UhGVs33OeTkpZnUJohlsQidTvvcfhLgDALERprThbHnjk9ARTt+Nu2lkJoDxcO57
mLgt8KQ4f/L2JOEH6S6uPDlVqwS9taMdDgIIug8ULi1PpftmOGLsVqW8LRRI5MAM
xf3GlqP5d023G2D0PaCFHFnS/lNbp6JSE8T8vGDR0AHFeTojk8ani4M/I7FT7yQt
GllptVa9Uxep605Ubxw0EhhKIHO1IGyOB1iyYSv2qjbn/ooZ3WriBfepCRFosa3m
boUECpz26gG6UYxtVuVkuRY79k+3HCsFuOzyZOC5wlvJDrpY+cngcjrweo8N2haX
Ci3lnzNvWhQ0JPVEPoO7JNPdiGbyjJFkvT4BZ5RGsZmtREtNIwUww4IPrdZWj0ez
DGfxzNvDlwcinQNJ2Bm/bGSA/HjSLRkGYeVLlcbFuBoY6AqGLk8Hmq1/GTxfgFi4
6tZ5nGZq2l9A/bVyh0EWbsVN0LipVWoVXle/eVVEkzk0ny39gW5BFefnBSOIuuh4
TGHS2nel7mZDOOJ8DSpJ9AJty2xtGh62s4pH4TZ0R4XoEUXoakOyI1jVgrpY1rwc
wPsfKeTpgaCsrzoO9/nBIhCAEG+GovuvrBpcdo6/UXqfK0WDSh3Y5l8ZDbkDhWqr
PKuKWjgMLJ/PWeo5iBsOs6ER9SYzTvplF3IKE5SocwxlhVT8WEqySNdG4qoynZIi
mcKdwSxFaqG2jLPJZ9rJzD5Js9ZpoOi9ToXfCVR/OVHAkuCxsxq+QHiyEMvhVAMr
X8MC/Xjg8nO5TXgohpxRmbanXuIxt0KOu2dBFHM4I9hnVm8w79PWsza0CqAMUUH3
kC+7YEvfbVeSp5PAo7tB4X7RzVNMxLc3eZly6Dp36E1vl5aCy66+vnc+b0tQoSXm
n6HnXIohnS7mmbcE2jC+hxRnFplxvTTUTDJpr502SSUxytv6/9j3TexD0k73fN5y
ENV8OrsDwrkrgpXr8Dw7xMKmzaMqOdMCPPjd3DDoeJuqJIPkn6TR4lULCilFb6Wj
kCO708mOUmgA1oX6SbWAPz34W5n2B4xOnTgtGGiZRvkwPpCgS9gANyYWQYfxKrj5
gRy850GVDP4wg4m7YKb4xD5+Q8/ogFGf34shAnUqV76K+IZuDKvB2yhUIckJ9s7B
YUL/ON/MBYbtbnAHgFKzpfMWkSJ94eCzAioJRAkRL5QQ8C3ZrrK1tEWcB5J3UEg3
Bz/OoKthksfF0Ys9+2Vcoycz7fWLl2t1hDMZdKjCsIXBHlOvmJBMxas7rJpNoM/U
ry0ClHj/XuKTWd7g278DMg07THyEQJWoeKhqXo3TLPDAGk/ek83cT90SndIPcu/0
WxVA397LekxfJ6Z16DjW/Z9Qk3fqszQq1p+8sjF1pdjzOnY5GoTtpdUxb5e//3Kg
CmjcL7R9Uzpzx/w/gA1Q5+syMrd9Ukoh/wJ1k5qgf5MZJrTaP1P+OSt06psGG+3S
Ynj7RQU7wrbe/nUGoqktx2U1kJvqM8Ovfw4epb4isaNkdElsv2LZsTFgWTGsLoVw
hgjLc/XF7DtmVdKbxKwRnOk10+M12fXD9ejQEEUH1TWGZiS5xnGA88uwp+cQIQ89
YS3deqU2bos6IOoa0xEaWSMTozyn2Fu4iPwcDmeHsnTHFf6vHK89LwxNhp5c0gJ2
QMbqbBNgzOXAwLUnuk5k5ubmZsfcoSLk2vZXrALQQHAQGDT//iZHzwllGr9/gT+a
4DyBLqzFTB+qa5Jcoe2hjKEuZY6y9aEh5jxWCD3lBofDdwfJZgbN+1Ljy6Xj7ueD
YV678HwK8tNh5MmL8Ra/gg+PusMHN4kaMOnLKQLz60SYc/uDlJKqIKhYbHMZmes6
J1THLKlbsVoR2O2xJEuLhO24nPIccBqL9UPLFgpZtyutzHd+QTUGJMYlFa9mofjj
2G+F+3/gJBQuWAyMuc3hzlNMX/k/XnXOMcieTrUGrzxhlfJzUibO6UhyREAfzuzz
TeQaCEnEbIjOkNzXsECkEt5Jeo1FeuLfUWSuUGL+Y9B+a9u0M39KBt45mejQ41Lb
w6YRFvZUsow9RgbFQDdbvsEMUsSHGSFLoYPRmlrQ2n/WkGLumDGlSS1yva+ljHBX
WvloEOpFJywyKnscsl1Zh395ThV1Hiy24/8msQ7xK8Wfz1MPcGghHtWxfgWBTfk+
0Tr165xhzVK2f3WjTdSUhs6d2dw6RJ0LOKecrfL2LuINQcjMRAwYneEXluCEmRFx
Z5viUj0pSaPv9kxNZz7QKBFru7zh+4fKxOzfzWYcAsnhpb/ojfc2RCK5/SvldBKY
oZkWGDfwpid4uqlvI0ffr28qy27PZlq8BM1r5+kjMYIXrwmq1sN7Vv0RrPv1sXYP
TEMrhK/7OL2dmY19ssBUYdxldID2huSkaT1JvkyM9fZRMOoClcOKKFbKKAHHft/g
FjjXs68L2ghaUAoBk8YxjuyiYJmApSStngYv13Yp+kBXWMFIkfaFNLvgH/PiiKkT
xn/vNO8hCKoJZg8dxweY2ZIltd3cc3iX09bEWQUAVePfHeJ/RhIrpU90XJ2aSMJU
tC52O8vqW+yUsPIAXCEytTGjDXcVaJBx4YjgWN0HaMzG4dTkBkseZRMZqDQaERow
g4fKOmVTn3M9T9bUAGqBxPjviK28ygMpEVWnjLvVTcNuUu1EH8z8k+/Gik5nVc2X
DRVhK3eL9p+QMx5oi66JN0MQan5M0+9DtwAHng9dFrGx1cPaJKXcgKW0GkRfjV3M
57wmm7wv+AcyOoGLE1Eat4jX14WiH+rLW+f2dupTG0wxhg+Ld5EmVUZJgVS8Cwlf
Lkn8KgVOEAFI/DA+NeHj0qvI2vaAK6yCkwtuuKBKVp+0lRVvm5EhYNreFlW6cuD/
coC2kj0jdlKzNsIPtR/IhQrMDMEIB9DqIBg12JvbxZL8x0NBWvlwIVIM/kAlkBba
tDg4qdtr6lKIwzgXSyLw5ZD1eiWpZSXt/6lfZPTqyJJaVUY+dM/H9LKkeoGptTex
eN/n8t28oqmrTI1uSYvctiJWQN2KnUo/+lEIC5lAuSCtgPRa9k20BXOeHndeHSak
kKmaTtldZjguUXVoivnSp57ZxUkv6efzsUhNiYrwNt2uJXZNLvPgxXgMNOdArvMP
ih6kfISfHUh7VmlHnDh6su+3HpW2g45JtS921Gb2bxHBUthoIePnaHOPinr5wei6
FZUviDnnF7jusLE6lvuygNmHkix1T+Bl7zeoozR0R0WM6SfxUaLlUiD+PKOMD7X5
+REvYaszv58/MWmGsKOIjDCVdLMScXlPyNHD9G9XDAfhwXGDTwVVkUc8QSRkx5ai
/Q0sqZUKcGHc1U7ulR6DEpFTwhOqkYyyO/3WUFsIPht6PlQPef+QWlnzJ8LMmxC3
DFZkajemyincSr5OYKP8271Fpd4YChLr4vdGuJNESSq4IUO+ZgymsT+6K1s8CQeH
kwDRQamxYR+qzwDCL/+57DSDRNSym+GQjC5P1EFH69FQ9StVB4birYDWb7f2n3oQ
cnHeClWVoAw4yw6mbAjUkcfxzcp70sJCjBe/RC+Tlhe6L1KDsjI833cJzw103jwt
hTf725qnxJYQ+MECK9ONCjOSlIIiWfH43q6lKR1kc7c6W5zbSkLFTtWXmfVEg1vu
nXNoriTELw9do4j8Q74V+4utsROzXZo7sVJhnqEduEABwiFCDl1huS13aJPX3Sxb
eKyc3ZR6STwNzjGvRTtgQexbeZxBpRQ2i6Ahxa2zWHJ61JvoxWdHVn4MhalR9Akd
YfEnOL3C5jTc4uZXDUaRrB7AoCuyU5ox09EiNDdh/NQFDc4cKNvTMGJ7f08g1zCN
X7yrp8NQHI7UqqXzUcoGl54euXXLAxzA2Kc0DkCxhRafojRnbqUpWgZWCIqO/+Ik
e2P4EkOydZgDtZCHHBty6JZheT9Gf4vAix4S+I3yrbyKHFB+mGjFInG00PRIdf1Y
mP9svdC6LJiVF9BWZOFd4C51wa8/Ny4nUssUAC3YiIJ9xfwVOeV/ayrtcmIVL/TZ
iG2p3yJx1864pa4BpHgzfpnxbTQvObBaItNXuuCYdZqLvVIVP8QE3/JHbm+AWswD
2mIJ7uMmLcfsEgbvHQSzBOm8tNEBeLMmplLFbtFSR1JhTHkFzTtlN6+XInJtUs+z
k5gYNP6nbaJij7sVfr53+8zL6PxQ6xoPkAiG76mmrk9iq6lXnOrFfvS8xSr77iqK
heMsZtKKPq3BabZEsRUYCBvmvLQ7s0OM3VBSOZIMe4uOxsqTFXvAarf7oM5CJnUe
RIK9Dh7d5OikalCBRC4jeb9pWNd4Jow9/mmqI1Z5YtrMd5ux56JM7PQsXD1+JuZ+
3+5pRVdvbYuT3N0a+yfQ4To25IDqRg2mhlgAkgxb0Kc+rjrYpbsRb2qTYUkK0VJn
Il4/m5lHEsnXqXNhrTMCsvNEVABeseITc8Gh6ocNxg0Xd4b4k4RrllS223P+xbaa
I6cdJ2HYMl7nuRVIjgKffoK1qg8S0+p/1PoejE/sh418v0HMwE5c6beyj5UOkkvQ
IeWnca30NZy8O6mzj1ULf2PXgEJci5uUy4eb4Xl5FbL1gXvLzeMzY0GyxaUTQTj5
V+THWlmOv7lur8yGTBzqLYGFCgxSPxlThKoQcDrEPY28ugHC8P8hdHOQJ/pl+JBe
AiT0G5xwnDyBp9MTncY6OFZ8ziPFSRYGkbV6GxDNYtKTm6c07RdX3CSkNYBsoNGT
s5phiQl4JeFndMRy4Ecf4KRgRhw+pYJgRg1gAdiVjo4fET5R0ZQ35k9LzuVCkRgC
1iGY8EreYIVxgwxwLJyQ7WmFOBybUaRwGA6l993eav/hW8I96/YfT3PDzIMJggn7
7KMt7mjaB6vjYbnzOksndJXLOST1KhPm5vDAtQfEPO22xHajBpt3RnI52FH3dps5
MtjGSw+ebMU6dWZLL3GsebTqMg+0+CboZ/1Z6QlnZPSTWZjEayphH+k59aV6zIv+
4JdfapcEb8iNeymTK8TtSKUIA//DpSkwZvD6B4nLA2bLrGGHtPOja9Lk13FcjHL6
rA7Dxo5TE1Meqm33t/7e5izPMAS2X9h83d6XCnnmCSDURS59CgXmJiXi6gEBBnTK
RO4fHl9vM1shpPXlv2AmjZktflnauuUtnuAOenfqNflu563XgkqDSgMvn/ytchai
VQv0d9vk094K9HCxsXCYLhshEb69JP8NWPf6L3c14B6oyTkXHSCHPca5JD8vUyyX
dpN2n3rkjsu5HZq9y7zsEKKGe2SEP84rvhBeCIfiJDGjYaQIn94yx7BhuXQyVOVp
flBLCL52bb0nRjGBlg9dCz41eXPfFOT4wcX2z+8T/i0J3IwBheFrA2driL4Y2ga0
uOKHU9m0MIDx0loO1G4ZPNRQeJxZoYASClIiKJtQZKEY8cUFzbTcjIb6pQHA8Puf
3W7UTpsj9y8z8kfeGyHFyND10+mXngsaDPznBTPQ5HbFgWRiU4Pf8jTEcdpesyK4
/OBOpRVSKU1hSNl/CHN7eWsP3OZ713c6KalZXZD4cdqQ9xHNkzRnniKz/wlXVyFu
mY8sO8ZUY+ohxV3nb3O6DazW1gaaN4PGw09gK9qa01uRWEic37Me19nA/jXn9BXv
Qrubj48U7HyUPvk9QHlQlEgA+K1IGsl2RABlpjzT/G5kL079g/1AbXmobmWCuGcX
cDj4+GY3LMUe7Zwq0QtKuKTo2U03wRH5K9KplOA63Ybs43g9J4QqdoHnXf9jcsQm
u8Z95O2HBEnUu87XouW0lUOqoBbHop70OFarlSj0mXtehG18Ou36+QrchTlRYgxx
y7fmc+vA5SVq+y1GxUCqVJH4rO4pRkf54T+w3F30CbfKU5QZtWppThSgbue94OZ7
kFpHjlNfR0JMyWNs9C2BkwW6euIeLxEzS0a81g6CpJfIYvaWj0cPxU8mC8Gv2xES
7HgHnA9mnglJl42Bt8+Brss/HT3AV1ll8qa30xyTADKol0TADcSMUdAc10sbRvuQ
l3OGrt1K7gGOBYTlcRDP8hy+NuhcJEWwz2z0ZuBX3CmWg+CIzDoVGbEnwwEK/qL2
Hfq2Z9rqkPN8kStz6xJOl/W7fXxyYx0Y498otKyDuRSuF41ELokXs2UbtWngFyW+
OpQOMp58M2ICD4aKzS8gAgqfWGPduORBSno+coOhmutw1zC4nCodFRyNovOOE2iD
0qpYMtzITWv7elpJm+ijtt03HUZclqi3YE0wXCUQxIy+hrokrlb6O3tEgrL4Ni4V
VVebii0Z21mvo/GpbwroUvMNXQRdd8Hms4cqGWTSZ53c94GLzRe5R7XtuYJOztyh
PV+jMoU0c9AM26B3GBN90hu/meztIC9u7DnU7T8P55aMSnHqueQgjCqTJiACMedB
aYaXU5vOSflYjgQdZuovgWtgTClE44YfUV5UpdMPndyLRGuSiD5jxhMO4s9sjvLb
P7eIo0dtimrLHFzwd9vTwwZfkf6ahTlYlHAwMHElwNNGb2LpAqQ1AUrkebMaWlv8
8Dm/5cizgDjE0U3MYs+9CechO5dsVHlSBko91P/iSiwMOyBXXcrBBhTyx5J5EzwF
GZ/XYzd/R1ZYdc1+lKVhpjM9sNYlWVdUzPRKmMNbiO9ra0a87ExG9cWOC6oFZrLX
s6ZZuwh3E5J0F8XOzR80OVp8CLFCkIJVnQiiW/m1qe+6efqvkSLfJvSEeh36ES5X
7jZb3Wlo1ZvFOQ1Vm+QwGEsdW7leERKcoJXIpF5uVPVutTkhye7L8JAZ+KYnbx1r
X5QpNBA3uzMpcBnKpTyIz+WHR8a87aXj0roWopd0cwkRNSYcg2DXvdqpKzRm7NcU
CQAiCIQc2V8NfIdWa6yIgbNMPX2ylv6Q5IDeGlZy0KEdIh27dj8tm2eiS3B0EQo+
MfHIg0axXTMjHWEAAGd3hEnODHOL98E8/s6ByaiZHjzmYptE6bNi7lKzsWE3T7Uq
aEFGD38cwclkgp2sdN45GVKw/p8pc6w7l501EwGiYgmmJfbsPCmYAV4cfaPHRSok
wPBe6hwPYFs9CWucNWWG5RM8FHA/0NEIUYvQw3wIqFnEAW1KF/uFDyavgsFTokGT
DngxyVS3cpn/TR6VvsYAwxlqJplgTSP6ffYVPSmtSw0sT2Y4M9JQJNvsQanZ4BSZ
2Ce19tHwNcB+PNkzME35nBWyyae+igxP5R0MHGd+0iI=
`pragma protect end_protected
