`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qFl1Hpk1iqNL7/wssvnRkaLj4HntHy87s8UhIO1RYQM60Xl19fJRJoahaPgNtpkH
wn07PJOp86+ZElhcqfZ+SmjFpR1FWCBPr9oK69cyIvlPqFMWjctZtbVWV4rn7HyA
fSi6nbxdtKmFxiSfqZtEy0Jin2G5c+E/Shbkm5cY15E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 109136)
LoWjUNmKOGBz0nAXpki7oQGvfegA50XqHzISycpIo2wOAdacJ8GAuExdVYG/zyHR
tn/v5/xxHOU4scib7k46HZEcgLrxvG1yP2XDipEY+dZnFVj2jLdgkvbWjXhxrXhz
YfT5Edox/RI7Y+DLkV4LPt4HDWlfzu7+vzbUBPbwescbqMXZFkfTRQk5/ox0uAgP
xGn6ZljhfhOkMwHPbH/kv/8uiIKw6M76X/I72ncGyqgLdjSA4uropcEc17X3rcSq
UwI1NnlfPpRf6QM/mJYhv6eMko24fb+h+2HsKhOCJfoOUhQxMADxyeU05PM0cmBv
O1Z1PQIosfxe3X21BX4VgqXB0CJYZQHIDz5V9nKuxCOcZ1zcZBOoqoECeYlXIxym
/TiYY4E0SzIju9umlAnzRMMAIPyNQGBB8YScy73siZ1GgkoQ0bXFS787T4stARlx
OPH6S6X4Uk9yREGDRDcPJe7GNmr8hy00kpWJExkEMYZ9IZUDBvRvxedyRTi6tUvU
jbkumbVZ72yYsOwNdIrDGbOEPMg+SzilAlfAVrBLQITZdqmE4T+rPOfjpq1yVFDc
TtHHIu3yPzpvcgBMIQ4TBY45W8dydQBlYYNORMBTU2TEhwINHB2tH1nQwnyr4wW0
AQfGSfpzxm9mcuVoCZiDtsXiT7jYaerFAA47kjqcUWslNQ40slHBG2HEPuWKq80P
pJK9Il+0L9R4p4hjDuh96PiqWQcfSddfROF0hRyDlsOg9ZOcp8WXYCzNvRo3AgIj
GXYTlL9YsTVxklXBTp8TAFfR+PzyGWxZOnB5Ebb3XGYdItA1LgLVJJCD2JF+WTFf
0Koq94OdE69za/Z4c0jtUucKZhpOodWwBI24PN0BbD1egpoubpTu/tEp9FYfYaON
NIPZKslS824fHridBp0sgSscj7BkdlQLBrR4pJILBy9Y4eNNNC0WQEt3L2aTdjA6
SzJit1sVlyk5TqXalu8J8KDzXGXRmiSOfdef0Bm8R/+n0/nic/THR3//lLXrZTOr
VgOu1HB2YqCw4dsz3gi9pXP3n4rJ4opRpfVNXwTpQzGtgoOp7itlXS9WEzhRdzEm
t3EhGMDl0AFGKbLIECm8L7D4yFNstcg9nQJkDY0zcishWwhGc7pVTnabh2uPi/rT
0n1Hp2PAZ/cGl9+wY1nvyvyEV7nGRlYbtYfCfa4W4LYgqn7hpa2qMRJO12XWLioQ
hGM51RteZjOfycxDIINtK11BNepuDsaiinqUQoR6mlOGLT42YEXp/Dl+WRA9+zJV
YGVwSz+cvRUaJwRLZuZhLOObmivUpCbmDZG33w3ODTDgb9ULtx6wCbq1W2KhpPpv
IdOk4S2uiV/WkiTno5nwsjddu3pr7tOV8uaQ2RAR9iJfd8WKl0beNJv50uY+3K1D
rt4nSSXnyD6+tDv4xp9MJnbwMQ89EExS8Fb5VIxlEFs4unb8Vg5ViUNVtUvyVC6V
x/Jexc8DxDNRCWB4vyRrzhA+/XLOiZRSMQdhiTKKSRYphgCU86Rjduc0ihifKQ6y
EJVVUklNevwldiarf4AfaZ7RqRrYatN7xJVgCjUOai5kDUnbLadTrht9kkcUz590
RjBKmscdXYGJb8Nknmw41HozoCYzK37wp/u5zNaJbKlqvpjopt6l39vktfk7Izyt
Lh4pO/uNCMQjI1SMkoBKURpi2t0GQIqlzz2HyKq5cm2/Ln6v6qZDjQdWNulrRWJR
bDR4mc4K1A3cKFEqRfTJCs/EuaAjSLg2BWbdbN5NM/N2l/I89IgwoJ4C6qtLFR3N
4kWz5qCDekBcfp3WG+xQVXuJeJSvvqNr500bSQQ5KiD6/N/QhADwhsHursVXCkVN
sFZCPo/UP2nNQqutcj+UPacu6dpzChexRSracRFQJ5+GI6kD88tEcA3GwiBHlDLb
m9MMIzsuV8046aU2+JN9vAIkEMREjPio8VLQ8aBYymJGiVv7hnQ3uUbgXnc6oZVe
VV14g84e7l3GrYLksBy+tE8Qn79/eJiYI50NugilM5frulwqqTEZ4Y1QXflXdPnO
6zgFo7Eh6JeZTQNuEGVs+RYa2SbqxccfYJOxLxZrd6MqhTARIaH5twggyhFg8qf6
fq0fFj0NSuzBq2iiFySyApc7lpvaIoASYkNqesyKXsbchLKTv8MHZ/Let1oyyO6N
9Fy96IjcsnFZdsOAkk38FrVRFUEsygdPPAU4q2e43U23K5L55CxpcefbU8bOlzw3
ZPVXTmfxO52jHmFtny0BOmi3zXOjp1RzItLr+DoUsgeBoH09RklA0L2QcjyJt00P
pfYs/q1idOfZ4b46J9EURDuxKcgLc5D/PAPbyWGUEMl/9P/HJVbbWf0BdvdoZxCU
6ue/C0QBNRa3jV7KoKWClblsuRYOA1vxiZCi61MJkxLM6bsEvlOf+Ch9xBP8zjVZ
Uhq0e1mLtBBH7LAltQYFbP9VnYx0jGAYl3mpw5nVeZv4FKr3ekIhdnVb13GfozQn
jNoIindOKVrNV8LJzNkgvxChmx7KKcx5HQYPh0EyXyfAzjjz+ttDkE+RmZbQgPB1
wkqZ6nL2P5B1FYkoijB3UaONaDQWmlCbZrj9qoYay1KtCFXhkCED7zWP9nE/daSd
3meH+91kzqkCrbAW+lEiezI7PkG0GPCNZYltow/CnWhspJN38qOyz1wXuv+Quoda
JHkxoAYKNnoyyf022qNjGMFz5Ru/vnWB2ynz3BOafuwYMbFnkyTFKUSCVvj+XFAs
VGzKbDyMBuVG9PPYmWv4x526hiMJ8eYuaqCRoVhgwa2VuIGgx9eNPgTuueINReNk
thlzZMTHgm5aHnZF3GqYc+HhofK7P5BUFJww9D9L6OuYuzeKXCT+A08ifVOOBwL3
ZmExYBtY9qCrWUxJimqjV/51+NR0rSjXM6AzfxxJgygxGGY2ImLafiAzEMNxOzV8
GNKSjAR3Qx3f5lH2gCQ6DUigriTTTnKLcWlNkUA1r4NVYruLzguRApMlcou/L5Fg
APcHYdxQljk1TRWH1eyWNZYw8HJdYu3zY5Td7iJ27qzOOTZJmX+DhF8pji6Kixny
8x14onI9v99dAPnSL6sJ5v0Wsiuoyo89AZQt0Mk8bwsvmD4C8HV/bfO9cqq2KnKg
JTQRMcpbmE4wdCb37CEk+DyqB45qkvkIBTXO8Qq+hkbr6JFeN2xzJ0w6W3MVe3dd
BpC/Gn+5h092pfSHRCQnq5r9h6JBG543N//m1+XGSULH93X24y0i/IX6dESZtfN5
PeH/xCTbpFLv6bRDlE0nWmO+4zi/teYDmrQ0j/fQXBYeZuWfYXcq87F04fNdQOxY
xcgdRpeVtEXND4drIXW6+HOZS6kYUn7PWK1P32VNFnktC8/5GNBC+FD5/4a7urp1
ME2qWzHPpsTNRvl7BAFwReANAghznGPM57T9xwNxbzbTmABJz3mgnYO9aJ3J8GOE
ugngnlVkNiddA7DoRdYgtyA2Me3R0D8HY/gw5G0GlmeR3qo1eETPd949Ej8S1Mwx
K5P5FyJiaNIsnujqehS1dbvfXWpuyqAkOekammFgxISzoLdpXLVQIyDO1NsvFI0N
XQD/wefxUztsJWsB7nSX7azwHOGKT6K4VumZOAaYiFynt+cTUaQii3N+HWI8G3R4
xkrYrqiZZTNwOe9k/Wa75Y/RYsVGKq/2fcFsmiXCE31nfV/67iqhMiM6TFLNwv7N
s+zBEJAYM9XsML/myOgd+lkpj9ikiMmpkA3svb+uCrt34Iqgtfw/BhqmJvoUzywj
VKP0hJy3NPOyNSArrol9Yj1Hq0+rVH6/I1Uxbt+6V9R+lbqtCc9X4wkvvAAJZn6Y
dd+eG5OvyX9G2QIVyvVplnr4GI3thR3m/9yTLbtxdc0p44Yc1e+l8HyeUIYyJHmb
i+uROx8kqRlNJMWw8F75p4Fa7Zaut3s4arhpSwpi0jGyiuAzoCMqfa4vy7YCEOtt
/8pVrFXi015RcTahYA3CaP5p3WZeHr9p/PjTtR5iwWLVXQUVqat0VshX2kq1/Xa8
b8viLO7eRoSkqbfBz/Y9safamw9/gZgKloN4h+HhQnoj5B5j7415D2xFjaBLCwHp
yBzqp/CKxzUQ+xSV+zi3sJSTtMKGQd3twhVPnikAZDemO4euenumkP1Nen8IEsYV
LAgwc1Gs41H4w83BCmDQIwzZcTQuwIig0p1reMNyCTXE2NC9R6EbqhQW7YCsRLaE
pK0vSAoraFWrRioHwdLOtMSXZE2oY4ZR09uSNwKtuQ8/8fxR0YWt17uYpNo52KI1
PwW40VBo9s8s+WYVRcrDP32W/CEvuy7on7zT4w74bYbl/CEgCRxDWXygIeoUrM3V
qvy+M+zyMH2hmL1MDJuuvShFdF5RxWDsxxfZVW+Rv0Ibkfh3wOGp+16IQMPTRn3e
ohNc0Ncb03gyooceavDN2VAMZBSgJd63IUjCFx2MhSocKItW6tOE4AJKqqBcHvNQ
YUNhPOsEZ+D7yS9JAhKhxhQYdvTJr91vhfqTWTnTw/TTdsBYG19A6sTWDk+Vv78v
VJ+5QKSHrh2UvN3t+zFQG6TSFD4sfBZ5jrrkXqXiXm+g3lvI++d6edsIZUH18iJH
TaAXbAIGqVaOiur9OT748JjYciehShVQG1Jnxk+HSfPr7yvAo3f+nETFJ9FJ9bVB
BRb3a1ZelOLNiCqf7wJl5/w3FrvAKug3mWiS15ZhZvuT03z0fdowbM3tV7HM3AHU
wjTsQgUKVPPp0/G2a9pVy6zOg1dsvAsqU0vTE9hdQxZ7/QrQBs/NKZur7TKVewyT
N9bgnWOgNImjhM2dwq7sVuLzKT7DKtAes0raMuRgwjDEjD5GMuivp5uglqlSKyM+
PwhdZFI3UyGV06CeGgXc0XXiAOoJr/Fq37BDBbxmbaYzzf2GVU8dCkGbBoZ2fIEI
6+BdK3Ebv/vJROogkTrsULGwWdQb/trr8cAoLOOwiIhBVxqXj5Bg7Z7UXpoCeFS8
+xujTOwuGwn8QOQG66j1h0kx9nliP0Qs1nR430Ixvw0b5rf3teYGSx+N7kP01aaj
7XgerU4KtWrbSqawjZPqk2lQXs4om6P3QZhhFCAdq5NpZ4xU94u4lcDd/IhrK2Jq
uLV43psg1FBTJQFgzQCCf/E/hyWFpdtrnf19/y8PAH5vmrreLZ09ecylxturvf56
bUuW6ofN0gVtvjTaSANI/QMQPvii8QfXN7qGJE0VNJwSpVwJHghk9IbIrbpEKKh/
7HwPJBuAl4YBzCdB/+uJDRZv+1BiNOWppl/zxPQvE5vDTf71SBc/cYklyxfzU/T/
2F2yAKZQb+nCD8Y4OASYZhUUa7cy7n1wbHTSsSX2ra4eDgngHcA3aX22Ygt2Vzoq
VD4nlifLnOa5nuoiDPKcFlC/aBgSxsRoHvIe5JoZ5He17QZgtMhe5RxgoNOXQfMl
1gjt3k8Y2NHOnZ++wAAXVdEAXtJzR/97vjznva7cwIXGX8FM5anIxxcSigz1S3Zc
ZnhViWfeaFsdS3mPj/ap4Y/l8rHXnse1QKjbpZATkrqivvTiWg/zZEaukNuG5Jjf
Pmb/9gd2VEj3JFxyjyMIjgJ04Ekz/Ibot/V5n/3HP82QCO5PQkYfJwgvYo9VpZCp
tiKWPK4b6Gmgo/mNT8j/LVKqEy9OvDcIk7mDVs1ILJaYUaYImewWAa3Y88fAH7Zx
c1qzAfTJccLMtlvebfZUXY1B4k1yWrECMBRI6I5sO03KDMKvAugQIcAY+y4WM/Y1
lmebgKJ8RGYjzC5fLTm5kvrFGUVgSLkR1h0NEtyWGlSnzObMO8ibrW1w1IzNjno4
wCGvQ+UXiYprQSDZYNLWbfsrYa8cRm6sVyum4db9J/sZ/zVbJCF09ipdqcGS9BsZ
+dN13XS97Cd+Vx7rkwc43NM5Pt1FEgR7k4nHszBsL0PMDtkYf2IoztRnIVtGDjmF
NUbGy9obxOZPkWIhSiImRalWCz3c2j6ApFRN2aOboCyX4/DmCsgDXoSXy8bukUqu
zfoItg+swt5KjByMMkb3RsfgaLqzVOWNvz/YiSjhCJZhOKRNXeuUDqI6L+eT52pd
vLGXZsCFBVTIfuHxlPP8Pe5dfwv/M7QtnQxPo01ituw7U8L5BQY7XP+MmbUSK+Wd
GfdjazVRLlkqb+60QKdloNsBN9m2OLdFKXYMJmnJVdGqqPji4/UXpzhzCcK//Ms0
jtjT+2rbHWhCKRmFBI3cvFhg7nMXZI11GKWstlHFbkpXjeqPRvYnjZeVshUUC/cJ
VLKYllQpMi4co+PO0pljZ2XbHU+N6WFsq9vpnUTyo/ItHDqH2nftAkwNvbJNVU/f
G3iujrzm/id+VRK/MZEp2BGpELhiw8GvB/j6aL8ywec9kxwfr5ySkzAxuxjg38YO
WwbNc0F83V4ispQjZgDyuaSUd2684xUqhmjciXIq//AigibPlOAbRmRD/xnqPZ0Q
7QobimcuKRmg+8Zf/zjRmmh6S7KO6IeXIpblnt3ZHcascl5Eq+URQ1iRTgK9yyLE
2CIfgnmFuYmiktvCg1YiRgnesKB3JnO8gYnjqizPUy3hiwWpYfYELAxlHR0DJSbh
L0vZzDYXdJ7IV5xPC2aZGt/dD39TRq2dNmqfcBpeFyRc8S4OvYZAahghfdhOAqSN
vDJXnCssqmwyES/F+meRcWr4Ald8nw4OxhqFbA1Plmx+fLqKGJ0Bio5m62bgy6uf
FYGWq4hy2+YSsfZZ2m3/nLINjD312D3laghjywkIVsvRInCO4Li4FVJ7plgH2aA/
SQ0E5qGN3N21PnMKRONYr/qUHqz5zBBXEDW82hGHm8q3SW8TMzvw6bERcnn6Ph2A
eZUeUjmyJSX2WmakWtp5FgzceS0X20f0HxITT/m38eyLb44DNFutvnNY9SXb75IA
YPEEVX/ZrNUUUbbcYAcl3m2fQj5s4QAJWjfsGydhjmJNTSXrIF/Ye5ILRGiuZVsC
ybTelFpxTYlTL2ub9FazpXEvelV6REXPmoN32O6QIj412GSqOj/+bhbAP0wMioHu
Da1HFtZhK8M3VXL0XaTwn1IFaeSx1yW0S55/pqT3kahUMPC/H1cQO4vuOL7goIMw
QGPvfIggvv51sYYR/LcVCxfLf0/A8A56CyhZ6+Jera0q5m8GFPedHUS21zeByTuu
IZEhusTCNrgZLRtnrtUoDnFphTk3ObpeFStq2Zu6t1DRIHsTbrkyUhz6kNYkhm26
/kEthh3sV+74kGNS/ClEeo+zJr9PWiCCG/4GZw6vKudewIAtlu+agjSABknxhTm8
YQr7o8jAxXoOObM938V07RrLBDjcv8cHfuvp8N5PXssxaQSGQsMt/sZVpxwWo5cv
jN2deag4iUO2pa4ZHtL3YGznxJTD7oYu2pg3KcGMQ6tU52/kPP943X84v4AEkTaU
Q2RHJwi51rR/HBzMYtaxwVI7eVwDTWcYavOEUd35rnDPQC/B3m4B6ZdOaAr7U82H
v9fG4+TwevGTnOhBGWbAXIaMEf5dZNe+ghaeEOPMynqrBLQ1z3nUh8/fdM+Z05X1
W8TIvYF2qF+ogCrS+QoPhjnUj43AGYzkF3zFy47P5+Hc0Gb0xyfVBjJATqER2yIY
OuTBcmmrYv0XvpYd3/pwvTB1h3J04pP3NE5OTel//and9u3SkBuqPFcrVBoc6dEt
5cAwhRwphzqZuTzSMjOn6FyBNlSa70AVIq0NocVA2pAiUfnD2tsdT+EtmtXHrVj6
gVqffjLTaK2MC8DyXJFIo7NW0A//0IJEnfRYXFkSjkZXnLcHifX1OIyknff0TVC6
yU8ejQWaR2uErSEOYv9YVw18Wak5ud6tb/+oFhUmapX7xlSMZWH+6ab+EnYd4IFu
AYPc1ElxHcsq/4DjeF3ZF+WJjNDOgLmJFF1ylIxhIBL+2HA63OayBVs5dfLj2uVT
FD4odMj+zvZvmeYyI7Ve9lDl71LECwiOdxc1FxV7GkIYup/kZAT4q9GAt6b3yGKR
zbPpHXmJX/zzo9Tg/kXgaGhuE1UE5obCs1lYTaqMcO8kvadVLey7TVOeCR3B7hpK
P3rqFDuafKYRf8iwRxWhSpGsB25I8Zl7NIIU8kalgQv1PwY9f+crgBd+5yRj9YOz
HJRUTKbJHXeCiYCjITWLytu6flITuywV/uGDqptILdUgB/vFZ/6Cw8OYfdrUg5Of
gQ7ZPGSm3KLnkmC/JM/OiZexLzopY5ANhVR3zc+yP9xaZF2MBBrYbA0ookqV2piR
kMUWYUkNfDyAvOcVeB4qE2cqbRbtcrABnzkP3eG3DFMUfc4ie4pk+Hpeo1p0akuj
yZSulbLQLNFdsnHpjiqsalvz2r2oQTqgWcaOp+yJf5ngn++Pmrt/c4kvwuyr8baK
raovKZklcYiAx4Q3vL/cIAEL7nipr815aZL4HhwSPHjwfRNZKtm4zYLs/n3UUNfs
bxxWb/QRDJYOmPalsgPKZlmIbHPHzg2+c2VBjWDJ9Hsl7yaUhfhUD0qh51+U7TJd
e3HdATk2L4m3ucfb431FLD6a4PKNCFJT/nmKbBeQr4Ce8r3N3JqRO7MUk/WgRINT
fbS62bFA7wRbXYKkgclrJsowTILeeOAHY7Fm7E13wy3t9o4QAjKeUb+gxdCvKl4o
jAPDq8yb/eaqh4ykUuVmL3jVabyTfeKiwV5MOMVzODY1SKwS+88lSn6jclpWxWRM
WDbqYTJxAzNmBj5aBipYhA/P0LB9qa9N1JZ354KuVpQ++0VzMF6V0EE1PS+BOdac
Ro/hWc9Yt5B6zbzOvbGBn0DyOSz9Q+IOsmcAjfzoRKjSZ20SnOLmLC6zY1YvKvBG
dOJ+IC3h/JMVeGOsPIJDBHqXtKlU5hCEQb3W6F9zK0Rh2SsjBgjOipJ/ktCDBeFi
sZvwDWtMtbzP+VbcB3st+vPKt3TrG1Yp6N1IbWYZ/LM2mzX78fbsY9/6/Bwx1sQc
CcZqsF5gopIWLqFY1UwJGX75C0aDUk07dMKxM7nAq/DGPQM4RyFosBIrZ0KtOQRO
MTrQyx8qEIpqLPmvOscuK0GHY6oQmRdcqFcEULSem045+76I8gAlW5ccFST1xMmz
fIAoA4XXiEJkT8XjW4yt1VhiSQskg8lu/eIA6EK2fboXOx3zkuMJs6GUbjkL77k2
kQHj39UrUrIK5kXkOiv7/ORSR/bIbxZfKTryCdyvooe2QXjtxnMEZpPnaPOng7C9
q4yPLpg/V7S/BVE2dDpDdONrUry/puznH9/u6OZGdZ9xPj0ynp+WtcugHwdCs9H/
7FlezSsrL+4QlCVa+vVkaxc2r9vjAuq8bZ3w2J14ofh1p0+po31HsIwVR1SrQY+v
bxEqsjXjTlT8D3jzGdWGcu2dBn6vPNAmkS+ETF1QiRizVu8IXkEQppNdT8vfU2Hl
QK11+sLmoBy1ZYwXsu9Ub2WbQ0SMprn7nFSR+aconCrILQVYss+KLj/0WtqByrL2
pxhn4d/uZ8Srl3wKytnAxNlai8C6j9JJHkrsTB9rDAJa611SkP2FSYOFWUO+kb1x
7VdJDnYc3DE6sKCgxVk8fA8sOEpkRyp8lkr+DETUU+YfaUuBFVP/OgvIhMqjkQpe
ctJmwBb8zd3rw6N/Q9wmhnaAR/uDNAitylzueVllJ8oEPdw5u/9waHo3a3thIUiU
PSCTxk2n9ga683Wki8iKvIYkN2z/e0STeSZT8Zvg5UVLB1LqKxTegRwUkVz27N/H
FbdnSXcqCghKPrIijShG/Nadl0HFhIAPsrQBcJGWmKEzqNvKgnqnPpAIr64uKOac
U79UZCpTacLtCj+SImSpLKJlRue5FQpLuLB3FzmLFXy8rWfOx7hxrvwu45ui0aLN
+J4Ic2lH5PruPfjOjPiaggp1orQblqO7jxbrS8tf9JyN8xJ2SHC0dHF4UYmz1GAN
uyWQYWS17wngfWz27xDtDMUTptUdHLO+edLKiJepbU0CPQil6kSyOt6+1sdkbCxz
1rktP0xwlyq+/KAjNhCptB2lqqZVUR6SgbdgXzs6R+m3/5nMxJNvcboYVnvdgvAe
2gwHzDmKg7dIhKnE4/EL5YSv8dsvlh5zoP+J+IV/I5I1Je/1PmZe+RhO4a1GYAPE
HdBVfDWJKbLgw1UkrYWr5NJuqe+Bn4oG1Q0ithR/fMLZB+H2NpO5td0o0EFz7wrL
WOuLyx1uR8WsiWQSOALGcs+z4rafgcAAR1f6BZsTFIbQDcCakonaKXKcBMsuo9tN
c1uuM9NnBjo2JqWDgbnFZTpNPC79C/lpxaoYyT6NPU0sS8Qlwvtank5FML3fsIMQ
xwx+FTfMdunK6sEGY8aG393wBiRulytF2vGEpJJGX+21aH32l1geBd7elGeqVrfv
PytgcKF55WwaPkjzNiPi+S5PQWXYcl0mp++r+OFkdb/Rmr/3dXdQEwHAVRS0hRXc
KFoAFaaK0/pGBJtTdi/GtM7T0f7+/0/lhMwxQARILhoVRoTHcm15mleTtxapRBC8
3hT3hNEyWIKClYCiglHHMSMOdOqahBguHS1R6NxwYtaJ//4ts3C7G5fOxZjuqIDc
xbU+dYPHD6yxWshdQPjFo0yL5G8cf/Hb0Nz4bQuuHCDWAItKtWG9BDrPLzO6N/Nd
D0bsUOk51c9zN8Ugup4w9quOJZefgV9y9/710c5g9DRViQbCPHHZyBusZm6SJBK9
fBCzBE5HJOMAc4ol6stZD7GdqdusfoVRX7urct2G7v3vxQzvsHFTTlfnNnQvkooG
sPA0LjlcHhcWOWT/h10our6cTyvGBVDbL8SlohDCxlNKvV1DbijbHLqT6/5XvoQ6
YmlNcRf9WiVY5Xo5aVOqn8RchMHI/lfSvzRpWZvNuwox+GWo7Y70R21bozdX3mF2
8zNIZg8Ji258kZ7Y0jw4jAaaCcM7zQO54RWcRi04iuV/gGSR1S8S4/1Z5ymlbHrE
dDaqKLKbmFEuI/aBIT5ZnvAMNkDRU0xVakhGfBokl8VNGzsyAHl3uM6F/GiEJxjQ
EESXcmck4ViNL7AM9l20StuPYdwKAcJG++U/3fmgDJgrX9Wq0BKdNB7bnmL6SvnC
X3wahYhZ1glnZ+KMi8UhXYp2lClIRzTz1BjCTqV9D0zlV3bW+0c8cWNQLm6xlDVE
by5xakJ9IfMxyf/2U/HF5gACDE1v/ZiXK6o5uidWiBaOZpOt0mPcNyCUDuceMl5Q
2Pi2mmE63L5ACN58Awy9n8avgKc01xIV5OwiDPjW72kPgM8jj0N1OUZQe5OiNEyf
7AnnnQENDFqeyD/7n2XHZ9za9DPMP6Oy8KGo1NSoKWpovhhkk7AjONbWLL4+hjAg
myaVZVvIxU+SdR/Xi74A60UGrsOgU2cMqthllKec3OlGj9v6tQhdH4/2F6VBuflB
3aIHA9Y70BEcGboYBN9exqtcAlRwS+5DhZ9KdMH4FgEVp9thIIxrchTldYSp0m8Z
NWx7+cqVbF4F2SSl+ULADmakNvegwD+r2AuIulm+BBYdeGi4OQfwsFCjuMYi2dcI
jr5+DjAYBydwvNKkcxlD2bIJ1RuKkLxorYDgX637AzMpj6UNdk5ppB7sdC2jM6IS
MNltGWEpQtzOy0DkNhKmhSZKhkm9exv7+buzEtMb2PtA0cpdBW/ypVDfP5kpYs5Y
rLpraKDEne3vsut9MpDA1GU0+Yfk+P5eMDuo+f9XfR6w7stY69fmHHAiazzoAR60
ljIA+E+NT9effWOxNm0BaDUBbU3gMBcoeO6mFiZrrSWahXVHAYWF75J53RarMy16
aDQ3s+E4jpwpsE6gPrvqV6EcwGyR1GUv6FnIqz2c7itCc3wIDCR88JHM/50zyJdb
TI/EbS/KBBE3l6pleJlWMbdeFBX4q29LwNwP6LdbMcsr6BYWTM4VXhunK994eGBP
DlWgsQuoa73DhL/CVoTX+abK4lkVoNP2O4LRW+M5sixdpxPalL0MUAiTETyJnzU5
lyEjRX26QhHcyHoWgeRR63QH4yXFyUDPhDeds8GZIisjwqxdSivDG7yy7j0+OSMV
ZF3jLsn6e1kHwzrsgRnsEsyb3C9aSAUC4emgFJjxEuJOaSXd8SWlB/AOu6zczU4y
mZ1qNzE6mE4TYRUqy3Ph67nb1KlVJ0MABUDl7iain+YRLMrO6O1j9Nx7E8Ue7NFd
1JGSy+j9U835PuuYLm6//ocygPSkKpm/bMRBCQGhesWMmYkJzTeX9jM5ZeQCk8K8
TnAZAXe8FDUu/jf+yEiwrCAVjLrOG61yGYdWsfo+s4M/PgodTpyP5VatQaCQNZV3
5OGfEpJK3WLmbJ9i2oX4MD1Dl9ZeNM6FQO7tweAyXFjJBiM7odyYXvHP7M0I5h+K
AJHrLqmGY17DLV2HhLYZg5f/+i/7b/s2Gi+KPXl5vAqkOh5QeDja4Tnm9hoJ8Bn3
cZl9lxMQy+jERqokqUTBFRrSE7v38K7ZzPukvkW2ctgVWL26TMVUtNySYo8iIQZP
UMgQ5SQzuBoZ/bwkyFjpMMKmG41LT21fjUnq36CuEpNSpXUDXMNsmkFpg+lka7cG
ch5xqvyPUqq47YF0aKJwGaXvmMquU2PWM9+uBYVZ3r2Kr10oeLvpH7nSKLx4LwXo
Z4atCqe9sdFYdZdtkq1JLJ7+uX0CTRGQTugj0imRhhWiuWnpvhCTKdevOPeuZMPO
kaOJPvhvvRJLnAtgFp4ZXjTLbmydebgrVFsP8evqr2RMFrRW8HcgaBr+edArNXgt
z1HsvCh9+4n/ZAla0iWWQdCxhgNDLcQnenlrCrljSDtY2yHn6lVLgRXhTQGExahp
RlUTPcOqk0HeEaaIpFgQ/UBCkM+pwXwa1m9iUEIC7o5Ito8hRDwCHKx1SU9WfLi7
LhaPH3OI3yuhKpWpszHmI8qhyK9FPuDVPv9Rp7V1ewSOOC0ONQeWTW8M7Y00aIBj
J633veJwFFHN4M/Y62FGnVKzQRDoWByno+hKlrCFN2rm0P10ZTXePrCMsBqqGl8M
mWKoLbzUFgrMdn7OJ/EFBjzz5zAttGgEg813QL4y/lvi8NFUMbDtg/7jjSakUzG6
lYa87BWflUAsE6JksENm+chEYk+VRQD4urvc9k3oUjJT0D3N09+WPNE+qe2aYMDK
b4pzFq0Rb5fEMrAeHS4VllxQL8Z/J1oAn4/6uAJIcgy3vpaKdYW+Znp4qGd0Q4Yv
mmi7yysr5Qjur/+SzwXEPwZveQQeHkG2UQo5IOXgp8CduK7ER1yhDiEQEseIgwTp
O5eTBobqXxjz0oKUHlVTRyXKBF9N+OIZ0mizWKHNMqL0eaIIq6yG6ItX4CcGxwVd
MPWjhHTToqAeOU0rPDpDniyFlYxhX6gqyYCBzzu4oNZKMfgsFvHifNiSzK2QPSvh
5/DB0FiWStqn4nQYw3evPXLzMqXMqkHvsZlYW65IwQc4T7X/K6q49lXiD3Iz6EKL
7E6kXDFwuis5J+6yfRTcqJ5kUKEuLY8QQxmmHm+qTRLdeAHM/1Yzp48YdGwyKNdB
PVV86Ec68rTM3ZEaRmDk9BYDoI+Q43pigJNgAu0VeoOFxe9WbZo5+1dOYXOkn71e
yw/TpNPQxzzJJEdrsyL56Qglsgj/T2Fx/7jp8ErC0jMlgx/yuiqcIwFL1yx0wObp
ZJMYSnjO2mgh17q1BSHyUSiofIRJ4V6M0MNzDlm4g0rRiuZQMVYN3nmVBsmQ0Dg+
PMxtidLcAm0KkNY+Sph8WOczXWunD0RKajHLdQXH7/oFVlbscOuWQbVTTNeql7/E
WYsX6WtorXcwdRB0AEIrxZSZ9tuAmNkxRgKya8fKJ2xdOZCbSzwOocia9X9baBr3
RFU5onof95rGRwqugjtaiNfKzMDFs2GeZZIg7H3YzRKsSz8axDv+dPZcW0QWiHtT
wvQ2v/waz3BJw5TVMv1frlWtU7zRKqS3V8HqL992k1svWyntcF6YVoUcLndZ4AlA
UZYBKq+yHH9n7uaqiS+rZhugr4Cuegwd0eN09a9jGomULPMX5RDRxqlKXlbHlcOR
oB0UfOfRBYpBmE0etzSo+I+sjYIsNzarkM4tQRWNoomxwizL/8WFEiMvJM1x/Oe7
IWajabGccsh07skMLAQthcdUX8R6JBnsKdnxQG0On8pouvsW0IrqqHgja9Pg3otV
tSLH6CSxCN95LiLnd/irSS2QCZ8c/MT2S9WnHNk3FJZA1KWKrrhwZfkoRZbTLNCS
JJewwfdcTWsWYfOnaIiBKwiCaKAirwP8GIZ/y5ZABWMERuarjBV4BGGgxLe6S8A0
/WgSRGp0yH6epIREKPU8hwk7SFlAcx6LwfXzX+IIc5yg/fkZO+FJW56HxxgHh15u
SJVFAWHW+JPMrGfCg/sFpqi8evMv43VJYuNUJhS+U62yK+ooc7eXeGRF6N4xqu0L
Qf8w8W+Ca7hZceWmOeoAFrol140KLL07t7FPTfRK8JgRDZQk59XPxUAPE3nUpvrn
tJX7tFl88dRntaKR3LX2dlHKT+v6ktyObQFV9/BvS9eT8+4EYdn/4HSzJjAzaCGL
Zc1MIe7c6fnmP6DFd/l5+oHPjIfdtc5A4zdgzWSUa9QeWn/YWzjIL9MYkuak7zAY
8NajG+kdLo3Av08tpNvJ7n1qdqakz/wAhDTShGQYS5K5gnN04RsuE58vsQfeUDia
ZWcsHk7EYcbgw86THLeNjEO5ecdp5viscxW4fRUIa6pXYTGhuRyDwi8eLyk+RidG
5QBwFj6WHoFeynmvNPrm3XjHUIjDHQeJO5zGezgGO8YVD3mGE4MFKnOGLL7EClG6
p5FMmQ4M6SzQqryZb11IP30aq4CGlnm3KVzkXlRtEVCb4/6qC/UkaVO14mbtL9ZG
Nrp7viEZ9ZcXqESAFjeTDBJzV4HLZk5L3HxYrCBIt9AD9lnaTshJeR0IcIarkbv2
Mgj888fomRFl1q55iAXDSZe14ZhiO4Cw7ld9kQk4/ar+NLCWcu8KgyoJZkHCwN32
33/nZLcJtgdmCpfZ94jnIFNeYOzJg+x1JqxYQn9LENxShhwHo3OE6QcPuDLkHgo3
dEegbqmoALskay/IqBOlt6oNKfIIbhJVmSXWI10r5pj67xtnTzjCuA2ni10dZXye
y1MD5X4wkQ1lQ5HKgkkSi5UMXeFG/tY3q9JIL0WKj3mfReG5JAMRX9pCruAYx+ku
6LbDpBfrBH5gktofK5cqtV/M2YGXRCy8OTKw+86726UwO9jaF39VVr6LBhVafe/g
vniKUFgJ3kUvIf5uN51OYjnLDGmQhqqfzZWInvn1JTyrgw/Qm6hjJXyUY+7gh6ug
0417Exafz2+04+xzlplysM+mIGtQlHnOSbUdm/FUBAbev4m7kVcwRQ5Jyo1v9lrD
tge4bHaDQ/f6dpmG0ynBsRR+CmneGY9GlJ4X4y4ZHcG+eWTYrSzp+zjTCbgNRRpe
sjRCZ+B2zWhW6rCaS4tXcfLzMWLnhwS1peLfilJbhQ6/kWGzXYuJ1J100ACb9Fxd
oC9av5k97m8gmQq4RXPrrYSW4y86hMzGKm954kn3xybTR+g5DUnhdwi0Q7I1P7Sn
9/M2yE1rgHgQcw1LsZNkesF2DYcnwCvi3adp4XPmH3oCukSgVV1DckRP8prxlzuL
vEVEik7kIobYs0VkwHr8PgykuVERnxOXFs1DU0ddsuNUcuOzowkkrfRO0axpmCOT
no4AF/pzbjI6Nzp5yW6AX8d04ZBWP6w9RMTBXxdST272odaeKsBLOfiimntNj0A0
fGJGHXl+SLwDUn/Yi6JmOlhrtH7JAVJ0cK8362y/nUZplNl0g+E5yRqidMjJGb8R
kCeWN7XOuBHH0kbdN7EL717JF3KZfXYEJXWLhttDAJp7rKHF4TrK/JB5BYQC+gOS
BqBb6Fu5vWLFcTd6RL/iSoKqSKJeyyhFkgTx6p2I6zgRaVSiLptT1NxvwUIUQBez
4M3Es8H8/pnxzKqPhTU4rcwUAKVpSRXQfs+5Sg+WdPkhem8sBFY12Tcep8vTV6H7
zuoQp7rRidchUIyC3ui/Gd51/AOQPJB/xPK/oaLDtleMD0zvoM291IrfMT1cyhT6
MAurrSEAVDYnSrwlgGT2DORXex9LkeoAS19qeiRdLPHk32QotTUqlkhz+8BpLKfY
TfFT7M8ulcmBupqxFaCMpPjkW54zfyR3dYzCQCeeAS+rWc1YbLxdOyCTSrkMrkW3
XS9roJ3P3GdjehzX13yhPKwn/xDq4aBZ2POGa1GNadpBv2gN3esArLZ3hSkgCLQf
eM6tvcgoOqKZZzcCbImlbriz0dky7xRamufzvY+Gn8Mpko4xWKb07tpJl/6MQ1jP
rorOY9awCuRRM4p1ty4Oi+XH0okvySPxQA8XWJmWGnQJWzj0pPLNGk31kKHdEyam
+KQZ0XNXC5z3QK/0x/Mhn5dwzrRxdIb04YdBOU5a1toWzxaGbdW+J75v+R4ilffH
oH2o8haGlea9pdnYO9/qHIaZ0TrO1nkoWI7go9UNmyupdlQs5dUWBc8fdpGXSD9u
BgkHLLBGH9YxA1CIEoYecytJj726DoN2NSJItjORxIkM72t81Ncik6z8PUK+A93x
hDaN7BrZ18N1pcMOQbHLLuVyGGUb3KEiMnlZU0SigClTHjz8Hz2+7fkXHIRz1dVS
7A1f3NK2R1vmUvEBA9Zg1oxARE9BMlhTb0WOw8hfNg0eZb/hQZNTJgW4wyQUYKC1
KYiJB+gkdf6D6M4vEAp0dOGsmdGONRS4w9E0G//pkBhPdluMobt/INJ7S5xUXcI+
InUnGvHyZTbuyV+uiYP4MKdrnCaOrJzRjBYEDobNVsAuw7AGI4WD72QcystPWy7z
wPPaQfc/RcJ5pQ0zVnITpyht5wx2u6HspxUqDi592pC/yr2Y2MYh/fyVIXDnFL37
OCIS4zcvy9DVu2wChDyEOpE8r80n1QQClx6yq6i4quEt+bPEJpZojEIF1txl3ylc
q4VnL4mJ6o0qg0yULgBnZKIgB7yzi3vxqpfUlkLtR9zMkug4qQCk00rbTNC3bTA5
3mGfFsDFasmrGWSrGLYZwR8sdqjTdDE9AMlq8XiSoGEXV7vBvC46iwMaIOM2mFQ9
060dorKBvQkEkRoH2ly3btFhTn5elhYnOGnIitpbOsQvmzHdxVr9thJY2yOhO06A
AHyokIsUeIpnlZRrfi3b+bditfNILlMWnhkVok61nyiXGx5ZhvfBg3ih2Qc8aOJ4
EzGb2vE1/YI833psYeJiubjST0PvTFEcI9Y6ZwcHiQrgL1Oz/fDjqPS4XdR+shUt
yILwds2J6MwK6R5L2eIhcjg4c3iED9TG+9bNd1xdMCM3Uvqac/pwSkPG5FgZAa5N
0DSowUu8CkDwJCHxzVI0NXcR7trPKGWOwEUt9wRnx6SYFDJpY667KBJmOvK+BzWs
hxhOlXCMskEnZbwH4Qy9PVTRvGAWEaAAdPYEHo3p3lv+XROuc803oF9n+mcCRKg1
ugpDOlWQjlqACtdKqTlDN6v5vBDsce9Ytx5T4iD/G2rSEghrR+AEfCgxVSznRA3f
BVMML+5B9r5+t3Xd4aG75FFe055AOnhx/OccXoW01KBnvha1Jv3t9qJfDWRzt4lX
TwiUmg55IvtSYaMlBMhtMuJPoLUyfkhwZxjdh38OMMONd37oYDdNE43QQbu7zuv+
gC6gNm2GLxP42DhMymWNskj1f6N5dGiBB42Yx3PniA1A8JiFHXJskqfKvG/HSSPD
f6Ws4a1jDmASb65VpUJKY9DB0WaK4tgJ3kD05nuoeEjCyYfG7LlFn3PY7sREisFT
0tLX/vFtpU/4hJF/pDUMl8JemRuKcSPQ3tJMYeJl/N9k3BLMCPgMO4elNYoPggJZ
SxJftI4euJh3SEC7fVcYwHY7/JBdBAzOrYucv0cI8FYG76Yy/fE4AVGQ6K8v90oD
iKAa8SsSe7+BnjwkFEcsTKfl7V6Q80BjNYPvwE++hQ8j1PRoZ/r/b30kC7sGl0Cl
VlHP5FfeyU43oJKuecWHHPZVw4Z2vu5vQ5RRvptoNpR7vQLcMtHdPuwbHiONPLft
WhJNuVo95kPHbRs29kjxe/b2loaZ+Rc2vL7jYVKr56UIfzE+P33MHxMX17kdO9yl
li2crTyZEzFNhdvfWxn6rioMvF4VdMtmmNPSz40ORoR4qQ/W2lvbOIzczFEWls9X
NU/9K7aRXmP4lvmUrGHRSIpeMGA5nZ6kJRywqASYEo9h/YmDmkvo6sN1UwkNuMwv
46LvMm51iusQhjsrGR/vP0Q6PJNs9AmFtPWrVhSgIAzUgmz8oYWmfMXDhFp3Qn+p
qsfpl+SQHjH8zAMWbEetXeAnQZetxUqInBIiduJo1qm7h+1awYIGYErt6hdVLykK
8v1IOqhxwPNn41CoTVKaTHPc8qEKn/+Ni8zpEJfcHt7g3UwOvPIXIhulLoL9VSqj
AP5WeMXFqzyy3qi/oEOLL5nijuaPR2RtbSaGqm5vyBVDX+jgx0JnZ5Ds2EJEr8+V
ILzFH4qWKeSle2Nvqaa2fXpy6dNNLqG+2ptH0OzgxRv8nLdrYan93yrI5OZY2+f2
kWfRhgOZgqWKrwZuxOQkH2UA3An/GXB8R2Bj1M5stEGEtxERIT8nKetTwMz05r91
MYFDoruW6ysKDnkq4aSh/RPHhz6YuEZ6ehJjJ+te7lM8PjY1+d2NeERwSJHQZ1B1
agQZzxTCoBXCRcHxPyn1GGmLLhPX75YUHW2btL6QTXh70s5tM/LqqLGSohu9ymuW
bma7bq030lpuUKwLAKDtJ/IIAwzVYiBr8PZLjOfccjnG0Fvc5reVCNa4pE09W5YO
nJ1L8IMr/hHkc7rS/1VUATGYPfynPR9uN4vBMxSPFqG301d3d1j8HUYl8ryXK0Ys
lBCEfBl18og2TbXX1axafRklLlCvgEICnRBRTSjLCL8Wclz9x6I1UOpNeDfU6XYk
OD+9Eie6Ue0Qj5mmIzoJ9hBejmeUVjSk30LO4dsY2/awtq5EJLrNsQx1CXl7CWJc
+WosLRVJwrn6LyRIaYggxGs56Y6gI0maIxwqUl2KatXW/HVpDgYni4exHOlREfPt
s9j3qSBKIHiWEBwPfzV4FsqZJXhb+wUT4luCVojigwgwWrawMxKQ5ntzfvr+ZXWC
p1kp5MVK2Gj0nxrM9zlmY+6I0JNz1hzWjcdSV2NWrbw7A5AZwBL1xZg9qdocdqP5
usa/ZXocAq6HnwZbnua1lwfSilZNjKYs1bStWx2ptSzw6lYbhLvdRTuDgG0kOBV1
AXUb/OOgMU14oFIHERYuGvUWhNS40Tu073hhAybyGvf91NJZZ3Pn2P/rIKtaLSi9
PwVQraBt5kP37uVqvyutI8402ltdMVxUU0nRytL51GZRJWGEx+fQTBMst/lhtIqg
IAlqadrSCpnuhggmk2VfnMiVkgDX86RMKqc2N+0b8lgue2IO6qwoSK5VAOYIeVT2
cxeeNrzG4lZ87RULUE5Ptk6us3HQr8uq8BxaVfUeGEsJGPcisK7wtztGqMVA95WU
VhQ5e20dLuU1IypFTboCRBHrvpR+id7z7BeEAfKp2pdGzdIFveNSXJJRsMfVF3mX
/UK6LHj6zexSMmjqHF7s+Xw4HD+lv5Icz9/RdlGaLJYUnnC15Tg8JOF0xCXRb00q
G5vg2ByqITgZOXrsWsINo4LA0O71jTSwqX/8fETnXyjSoP0eB0tUiEVBvNZYa750
si0/XuY09iO1oEzNsaudn5uosGxDRM91zw+Av/V+Dslr5UgBBrRfQJCK6CkMQocs
cUw7BJ6bwz0IX/kFKCzFxJo+mqv+wQbX9Rdhrwu21GafGZKUXal7juAJ1FqYaH+/
M5FHtrCNyk74Pqd8d1pKlF4GDUpAB8YKgzIjiitKH4KYlLeXGg6FnIa8XiUMUCl3
EsyeTS2Tt6Exm6ih2fmlBL6JrU4pVX9RvWQojNDHsjeIMu9Zn85uo3lnbXbqrPvX
dYqOmtMepExIBzdYO0Poj91z7CCEHB+z5GBkT5BZFJ3XARkyArqB06ZLcWMRxBPt
EAZlSFZjn+t1lsMxgvz7Z2AEVq12C9gsTZMJN7RmDojkJEMfDZ2Txs19ACWi42tN
mwVjfI/RR28MVIHDh5jWy292rPQXzgbyLNBzuXijvDtDM75ZnxSkJZKO+NhSLK+t
o2SIrCtfotohzwqb3fp9eRVIoiPsTKrbLQ5ioiewRPX5BI3HZRWdGgxs89l+jsfm
dFYF1tx1xMlgVuUt4oFOtHzGGJn1tfaDvzfu6sf4c6rmU5SutF5goO9Y2COIti3+
YQtOPwsX3aSbrp9y0OJc956xtT6wMDOXfRMC+15Gm6Qf/l5JL+a4kCPbhzbaywaV
7FGEfscRefq3tlebQYrxPIHTiVELNgLIKZmv8Gb1arF7+6wMsKQFlrShw5q/fvlN
796+WVsdB/U1SkZWusW5jj/AVQNjrt5p170rn8y5XAdVSsbJPrBRofJtNGwHSdUo
4qEHXaA1i3u2uUr6Mk6W0AfVs70XvAKIFNNwKb+vH8xycqnYcQ1diJaby4ioF42/
ihjLHAtohSxpEr0r30I9QcusU7nnP6HUorYYUoFn1QyJqqXhYUbQWrrzbmV+LjFI
/CW3jhNNOZVFQwhTDrIpqctS5978Cv+DSIDoXzlSQ7KhFIZZcaPWYs5GAsg+YhMI
xuzEFdfShFFLYtm2V54oUk3JnC35bGLjxkI2tsj1Xqwg5ZjV2+Sq0rDNCqk8aquW
Y5bDpnlaWrmPDO5AGwwFl0jDL65hW7ckduCePwR/MtXb4vmRiG0+wny94fwpcqsH
8rR71B4k/p2d0AY0HhCpCTZMzWmdUQx2+qOjOQ+YerTLKHuJgDmTb5dIIS/NZQf7
0T3PLjY84ypKtLnbRWf9QVJMNDRa2yztJC3JxCO3gytK74VP1Yk3uBXBXJiEJnLC
7iqG6mis8+nO2lQ9KMbfxgs3SdKWFC0BoDr8aU512H6PQKoLtlkzsgfKE8IOXKAo
pkcH0R6z/w9pzxG0iITiSzg1h/yfmRR/AhtK+dyc8cq74rIOwINyNelzbqjKuebo
Udoaj+tzs6Ey4JdFqBvITcAxSwqdftFhoOVW3X12v/bCVnTxcRiEsYmWZSMoSYdg
AU7G6jrfNmctbwDvxsAJ3YUpmLlxUWUjEdxOPRidwLyuc9CN33L/5SWkgFVCXnr3
o5WYTb97RRnyCf7lJ0BDxNJsvZ5GXHIep+EVinYSCAjIXGSvY6RsnLc33MTTIR+m
53SAnJOG/T8zx/lO/Y9EvNtm3SFHCc+9lynmp66ruz1o5Tlse+zDyth2OD594EYT
Sh6Qv3G3/EJCBOismnX/KZXaXgpdicHcSgEKp37moapES5zMnNcBD3BBb9Yul2NS
0+rWINJRDmJUyx/vgBy3wfIvNNVCE/PQKsxxh2e4j8Nwn6b0+irTgNzqlnI1mw7L
aJzt7BTVL5QTWZ8SjzsOWCyZqJek8BrSrMmGSsjy4tCO9rITZvwlBNpjnbXPGz9v
2JnZUu7snh/ig+zDYyQlaA4qSlDLVv9U7USmUO0erhCZ4nS2RNQmxGP+HrJ7lZfk
5e2Nm/Xx4EgAwambEFSzL66r/5Fp3UJ1dKk9tYf8LQoXo6CgTYbtuLgCEEoZENgP
qefJz+ZcRQ92cGaQg+xskON4aGss7ymLrw7ksXWKdmuraBDDaEt7+k8ZQO0HB5xc
352qg4GKkX1SCNQca/dfWBmf/OKdlymIKrsmMnURLBJXGFm7rbdOe1QG0YhDL18x
YEtToJfU2ELFCi7jfqqw5FdwnkHasPFXD170/6arBrmfdLBX+aDfW+iUtYdmL77D
kMi6kMNjr9PwfOETsm7PU6Yoj4BWEtgpygb08Z5+HxRHMIH/HJyzUazl5AAHSVfs
RbdU2vrhNiW8sS3pGXex9PQRqYd4Q8wMkHsiHQF31aSTmy8uK3FcmgAjz0x8j0ij
yiclC19EIvrzOEG5D/0kpIQjmqLK1t+j7NlMdJEKaRougAM+mnmDyFGs7SW3fDQU
16z0lk7Cy4B4hS3jLLt0BAcA7b1BYeSLYtuqUFV/co5eQKCVHp7XP025H0JZK7+U
CMfRP4h6d6dTHxbvOWRRVnIBK2ZRjYajzaWQ7Hp+TFwUiD5jlUwUxdgDhM0v5L+8
/mMUZWvVkGLzathG7kN55X+CfJTV+1a2q4EyTnQJMM5B9QwuoiEPy3vdrvS6vRYK
HXZB4BpILYPLPAgcCkOqpzUvcEngSY65MzZEQZWR798DMb4qj1exwACA5eXJ3rkp
TevSo//pGY/uKQ4c9OLO+Us/5blus3drVefXU7Gg4e1XYJC/BgraTSh2buJEeoUY
WlrkBGCUPoLIgCQb+1EtBz/12lDPVwD1oPYA6/pdWMDhLdcaTkSYpHYbhZOajn8X
h6KhrW/A3T8zIdkypj+4Z7b+BlCcf+de95rvBy3XjB+2CXK4tN73y3I73ZGK7jVx
Yj9tfyuPxeDRRn9BK+R4umgQ5DQ0AC7VVlR4HpHH4cE56ZVXm4WHsODjK+OFEjPq
2DhNbHumBzI0XIb7SZjyx77ZX0tmleNjIPwu91//fBM+xbpixXjJiw34tPb0dQF4
tjaddHyTGd7O3p5qrY2FJAE7u816brOQEah0P06Z9BZsJO7piP52H5IAYedkOkIR
IA0qEjsLIba1opP/zLwOPo71rI4A2iWPd74Yiva0Y9RCV1TwYpfj3DrFicFvp/zP
O8TC8+IHzcSYddvvgZx5OXV7UoClqhaVgg1D8wQtpW/6PXJTrDz2bdVewzPNHqqS
ONl81SZTB0+HkMSBDkf1QxwqRvt3BO2BKJcg4EXCujprmzaNxNdzdZTgw214E/UD
uHGUShRKwGc2FuJe6eccWazhuarDI2UCgGOTCq5cf+3RWS7nJ6TNSW+CHyTVMIwQ
+Rx8YK+mrfcOb1uSrN0OX1nf6H7mEnhHe56hC6Y2LpDX30mgeN6V6D9B8tVqh9oN
9Gc8ld2gn+gt1XIGW0fgkvPl30eEghOd+srD3nXgewnUhwwlmUYzOF2yyiOgMTlN
tPOKk92MKa/EMxbAYKO8IZ4sjGwDGz+Hei6EU8IemlGbu2B/6qfa+FoYf+awjHKI
I471qHZHGuUrcTPiM89ftLdhRZwfZ2lveBNyZ/ncgFsRM6RgPozHeYqF/vNvTiew
sta8XVRNHvQF053RuJomyuSE6Gg2BrKwj/FnR4LVlIjVSBCwStUfjJax+2c2hCTo
d1TuFTI8uC5Zzp6qFj3IjF6op3c8ZuU/h9x3CH6LeKr9ZDAlGdfu0x/6o91+x2SO
Nw42C7U6UzhlY+2/4VLSUDM4kyLT0EpLzc+8VzOrK4dHpLlAXj2rUrvneCfGcz+M
Ng4u7uFBmxcdnb3K1c5nczNZ3QAWxja86YoQvdZe+pf7APjgF4he08VhGo1tmBja
3SG85p0uleOWau4KYzvKUaeVvnSV8r4l9QldmZtcceXM8Z7oOFCTexY4Z+48PAJC
O0zk9B/a8wu2z7DE9DNDysxFnEdc4gdakQnx3u/2Auh8FJgL4B6CLghOFhO1PSXC
5HjzE/qPtFXS1f/sWrRY5f/LLxO7OiYGE3VCd13Y4e2vGTqaKqzJnrT2Vu60GNLL
h4/5GJ7JndN4+5sUD5w9IgLqrvQ+gLy+XYUM5F9gHppf4SPoraiakqKFza+8XHFT
SPdMZU50Ux+Nn+QhZWjXNnNFVkpR86hdx8ZbTze4O4rWbmlQ/7n6oTLOW9JSPKlR
jpVU3Ydrlfx6vUPlPJM/4pzGPIMm92n4676WBJGT0fdnJAAXxj9PTUCG0XNkyBim
SGeFO9SgnUuTQONnlYAS/OKvJ6saqsjOb5ny2t9kxLik0X/G6W2qwtz4H8g+49pa
jLChxwaM8JnXWDitvYqzpls74ho7N4EWoiQU1jQYS2uLhwagGFnaBu0BJujbrHRH
7GG3ZCHjHcHCks09DEsxpj3fa5GKbxx09tcWXSUuUYfSoaWQkynejfs/eBzHkuxV
u+QfVaTZt/RCX1uUWhNmOUBE8gfWg/A7JVS8EfyFXm1GlwVmCdY8DvtmCK4kzJko
zP1lEEH6OkONKFbdyBF0KnYeAW8IHzZrwdgyd6aZGHarnPjxIrJMrswu+NyniFbL
SvxykU2+ULQnC0bLcVNBuzU+Xnt53IK0lvJPDj+xRzi6rIqqG5HqbLjCaH3Kl4yQ
iTYyqFGABqFXWh3WMjtFhNo9A+1PkrbJUeP0TX8H7BNDgm4JZlycXcHzs4FXIOlw
RQpCGz18TrtDazLN6gDvIMWQRnueydL243jdHZYVdJ80Rr7hIhjMO5qEDx8oq8Qf
D/kTEC34iWPEeb85EB/hJ78DHkueTVceOggv8CYsXXI/u/J4YpyfsY/ywsql45ik
jF9MLQKx0+3BWaxTSw6WusmNZb0aRlLB9TpHhcRBipXRVrdu7TEg2wscIv73y5Tg
RaCQahzIEmOOTP8wJOp6qI+tbu0Acd9hsEq36nSxoNL86wE0GGMocRrS0ySZPA0k
fsiTGDEYPts9+VrwuRa4hSDNYY2dJxSEVK4m0z2Vr1iaH95UiUFYULcwcr+pA9qN
0UXlZ05oUiwCFHLUHskRaDLVPmj9qYFNELzj+j40Knr4yJVX0BeHpUgA1NfPhP28
RtspdD8dT7pu722azIQMWd0QOfMTTECKVB8ozQWgQ/T7mhoL3+NtWYIRcQPjP+6d
DOxrNFmCj8p7fmMCN8TN2xHksb2o15i8OkKmcbXtEEhyTku/MLD/jjSP6y+jiKrC
CcE0z94a2FJrnNvtmKbKht8bDLfRo/UDdYRmbfYDWX63nqiT8NHighhJXgNOYQcp
bzJ7K2Ar5dSgnNtZVLPtslNutdZvd/Hz9RdRVbB00hYOe4pab8iWwlE0EEX1BLVS
ywcRwX1xWTWlgfoQu3u07HP7MAe9AfBH86PGhM7ctZnDLzeJzhcwynF+ANe39sHD
St3vrx81Ru0Z2jgd16RMVt/DWisQJbLFHjziM/LHYI5MbeRXoUBvBbYlNAMmO+ar
I7MiqeLISdyEUsl3N26HFXLWU0xf+uNCufYbMMQXFth/bg/IrxqVItiN3kPubOFn
DCuJRxdaRCQ984v9+8IZRXW1IOBTI80UWoq0qaWzxliERJXm/q34k3V2RZmqmN8A
aWfz9h4KbTbZBxrUbZjlfZV8/FFr3oJaXx9qQI1D/+AuA+OWOf/XBVcRKI6Xi5js
I+m5caOim98dVllFV6YpcX43uOqMFW9KdLEur7827Obt8DUNXKP+gIFgKLkhaOos
PVF06YuARMZVFf0P+DDd7KqQo81dxv1U5hH/SnxFAd0MwdMNqnfQ/zsjP3dmpxzJ
QU6x/CdtrcpSCfbnCFWPMfwfm2XT2Or1MNpmAUSczEoeEdyh90pZC787fj03yR/4
cBa0cwlQSsG1Ejz0HGb61p7WrX5RM0kk3fLfHTqjVX7q0pUfrSRDGlmxoFjAxlJW
WCMaI2wuRK3rWnOsLxzO87BJ8oI1IYD8Dycg2uJUkXO9yzMt92wLtOw4gIfYfHo8
QFnxZzgeG9PKJDTTHtO323ItQ3htY49i5Eww2rDfPHPldjkCHohXlm/mWm64d0iM
ir7HfQc/YfvhCTK+/BggnVcJWQ5wbYIB04NYhp9B+EO4v2VLHsoB9nTyStj+hwMH
Z2u/qGlCVZx/rnNWfum9FrUHU5S9GWcWLWE++6rOiXEm8za6IOHwxT8OtjXBYdJM
xysRyWI1jIzikzboYlIGyQz6ZEFY17R5Akln+rJJdieiKFNIpjsMuYqdYBbdhr0T
9DbFncg+nO6aJq6CYe6Al+tD4L1BFmm0AjT4ksaqqSwnAkUs+boWk4tsv/8DvJj0
cIF/OYZqGPi0qkAFTn97t/rfGr7zJu4GeiMtTs55D6DY7dRBXfbWrB/a5nT10zrR
gHjZ8x+v0c+AxHGgGs/4McQl4c3MCnV9iSyiFxag+TZIcPHich2IKWNUtHyfLd4f
9P8neN57o+4J/j2RNMfMANvc4MmuIW85PdvJo0TS+rX7RWlr9lcThERbhoPkntoS
jq77IvpPKejXrZn3L0EW1oHLCrNIFNJkdmjWXW8cNC4FnY1hG7q8z8KpFTUOSvr9
fP5vFolG2wQovhUPou9BaZJCmTRLKVamxdEsBNev6QQEqLeuk8l1fqqnAh6pzKnH
F57UHwMl6fSE3MdjNSepCEZo/XCXO0oXZmkYrLu7TlHEX1alm/J5kGQsbu4FLAx3
nPuZwGmJ6CQltlbyqClF5V1YaXSIbuvF0TOgaTkAm/TrrssHsHpey27PgmWx1WRp
udR8rcv9Ci57LS1Dl/+0RAYqZpFNAo6tmjgEdAxhLWTgfsYBdWv7bEPRhURr7e3x
JxS3ha4cSchDTthPyTjKlXlswVVb0j9MQWBt1oAa6RikFBFkPDXBp/ctcn2lRnbV
FJrXXZgrlamkQCRvs/VEgsyp18pXQf/9oZ5jnZ3SMgzcoXGXUaQEBwwkZWDYG5ir
KVch2JdwLfNh117E42OmLS6USL0fAyp92iFqR1RBbGOdQM08xvORHkZLKXe9TNtR
ZWYqfne98voI0pJcWSiHksmIsmfPF1nOBLmheSa/Q+UkAx2UNooLFLBTdFEJSXlY
1A35cWp/kE/V/TtkPVKhCuLLugVnT6CkGrAepo1tnxTS6gw8PMR86W7TH3CrGmS7
8IrSSG9QxbEyDGq3sBkYPrshcvGqG5D6bGhi6CCWuO3MZ5o8OpvHgCZjNVmVWOOV
icFAmRRoTIUMK7hM8cuU84CYVWPSdyECqfLE0hENvFV4quHMDisitSBYWe0Me56u
MfLYVjvtYWuSXziGZBlGzwlzI8Lm4s/lQAAkvRJxR1QZGQ7fmwS9CtNbi4yE4nXz
dIN+EDD6FWG0qSTlcMdkNuPMJxbPcJc/6GWGek4EIzyNb+bh5pn7NxL434EWY5YN
WI0+dERLylAJZxcNlF1NkAq4Rqil1cm6zs6O0S7dptxVIFEMwALLuLEO/bBukQcj
wP7rWy/Avp5t5Czjv5FcHd6gkSuSBkathcC9JKm8K2RizFn+v9rY/BCqmFUfoQYx
kBlgxI4vXwkuoxC8oz46nJ3PCeG9w8TSfGk6jE66hflXalPS8ph6PAcLejl6Oq1c
wAg7mZzuYD2CLJvyuqNVBB7dJGnd9e8MLwS+dRNsP8cBTfsjVN67hixxKpRQ3rhu
TFJSwVWlvuW4EV142WrdRvTFAQCOpAguXyE+I4JSdSpL2Facofmbofz06QBQ2FUa
gEIGYGVSb1TA1JlbfDosHyOC/DL0PCT3ZHvQRexR12VVHJBNbbeS9YzjDKdAnyO+
qBhzFqcG+DvknPNCklRItg2jCWE8BG7ZQWrWKDY6tfUd8CTJw6VON44I/xdZOjcq
OKeo3eQtStUjX6MZevVJxUKqimWRUbiC6NMothbMmwpOfTViLZp54v3jMG2VukDT
vr0D32XetqCB3343oZYLC1UYg4t0ihZvA1lm/AXkHHH8ab/mJmnaW+KAC+F7boge
dLCzLuMjqLE1Rhsy+5uABjh+g8e+oU7uv6GJKe+ugPl3JJVniXmF3SL+IzwNwppA
e2r2oL5QU4tpLJ2103TUTsQSAXbyevNAu4Kkt7qKosE+LYsZlXh0cE2xXLml7NyV
zEB+cdXs4IBjqF+oiqKYk1HmNb1eGASfRvrSyzWCLZHbCTbz8v6yB4f4PxPKfMsm
ehru2+NjUBpEFVub22fTRylRgva6p/NGUFldmsR/q77Z3wk/o0pC++SmiPYkabX0
8JgKlPKpD/Y1T/NVie+DMPNsAVBQ5QYeeAw5fls+NcNS1MZUkvHJxPO3BQvOFdIX
CCdnWXF8O8JBbihr52IdNQSW2xCRIGVBuWdW4DW/lxwYgql8oM36rS+iFbTuxZ6w
quv1DBKN6vm/0XnI9PvfK+y/VjlnT7dvJSZVAbgCCkw03GB/nFJy3BiF+08+UawI
bXpoewqUDWxnCa/Qx+y1CMlZ6B7MLyr7oQv5jFT1NvBQQdjl0tGFL5cji4RIWNJL
hZ1lBk3tWdLckSYKs1ke5+t6WXWfCMEbYY4CyEZtb6ohCXJxhIUBNk6omPsIOgQT
+/8aJTvZOO3Wr/Px7KUZS0bAXlS6G13sPt0kv5zlU5uN8/uz0OLdWhhZKgNkCUOc
FP5dd6pDULRApRBJS5CyIL8cRIfZ8PAFE4T07eKz0SehsU+n0cYsFViDoQC6ZoYI
Ao1l1X1q5daxtm8hbZif99EnWzJt2Z4wHl/y9LcqfJ9JJTr69G9L8jG9iTwL7kiE
F9ApzBnj4mAFMHHlSrI737d9gbCaJa04fu80NMnjq/hOaNF+WRnxjJPTa9I2/z5g
vIGHBgldsIoQKcio9GUF1oHTKMsMiGTh3vryUcigXwh0400IeomsOSdm5X5BRLoQ
GPNp4mRMoWoGm9nq3i7HjEyOEVgYf5G06m8rN0ZRz/CLd5CjboDu/c+pLU9PP0je
L34QKMKjyjFjCUVhXSvDUvdPqJLdwI8PP4cZXjXnWACbAERH8ZrrKDrsTGsjnwLv
EspgRcixSgDmXvQvNH0mYQjsdQMDXiZ9rk7BstsrRmAT6Vlb3Lm1xFSkrq1qK/cL
mpXInXrjnlAAPotXLQo3XPwy0I1RhIGND7ZzvYnb80sWmlcF2LkKGa8XrgI0X4zk
3tB3+Pi0xZRrn6jEd4OS/L0Hb8XdKb7Tt586xv9itnBYHvdMDbsy/0iXIOUfHVW3
vRgpH68YBKm8a5Huh1ftKMRwOgVHaBqzSzB7kA1DLFInFVCPKHq5nK2/Yr79D9VB
qF7isH4mVGuaV0jKpVuHV8zhRog+dZbaDtUSV1Gz9ikXAFzfJ10cqUJPW7l1+ESQ
1rprwbxdPjoQRg8bJVfdrlGMQUQyto2HEFhVFVvoGHhr5doq1TNU2gmXsRll8gMY
vi0/BAjZg6G259ZvIBK+gd6Kn/9DHOTiOy1BSQhgySYBHhuTz7QDI0na++wDjflM
OKduZlhJ7bfu9z2TgqClPecw/IClODfA9ByqAM9PqSQn0NfcxLHVtzBs/FTuwxPO
6o/hXgPx83eza8W4rwRPlYlfA9ytXz9kkdXj6ux9MBJTxGLNwAZ8VVtMMj5btqZL
oS0sHOepOeX10sw+NggsuxLK7AMZEopZau62dqOwzq2txz6CycCAh9PSO4QLdWjH
3Hlr9uKdw+uWKyWAOD88ZHyT0o0nrNZAa88xGLTxitE+fUsdqhMGBGOcrnLRPCJw
PTpwGbZR25fQjuHzSIfW5tZxvyVJjHCi7n5u4O+toZV87V6wcCu7tEQC9lWjtERh
9W2+oEUQzzEhXQcSGyq77FHnE5rSCTFgUWFyRcfB4y2gmCJ47uYhKTbpB57Zevl/
5SCgiHxd+Y4Zib4RwQnfNhWIXJ7iKCrClFFlq7v4dCpAowrbq1njNw0gREyPC8WS
wIRZx3gA8SRhyOtJ66713NJtuvb7kBO3M7/aXEGI5m5fOZkdMRGRTmAMRhE4uEJ/
D76h9eWaJ/pYIrDjCcVo18LDNp6oAzN8LuNtAMpvvLBhhDfX3WFarWqlCYoAxe08
Rybb54gDCeY6ZgbOhXbpVBp/iAUW1w9r3wsC0uM1XtlfWDfupDri0zlueb2RwC1P
FjY0FYQFtI+YJZeyQeDG29l5Iq5JtH+hn+pgoF0WqmORhti+ay8I1JCChfenMY25
4tAPh0NZmGOjDkAyByhy3L2fLFOfk2pS9uBHcS13OLVzVsHAItWIbOtuiXO6V7HE
dPTfOs8veJPR6nkqwV4s9hC+AFbxvAzd8tC0JHt915ChbV461FI1OHqK4izSpPDx
5fdtYmxz79QiVKCYXWA4YDBVWD6FCf9QaZtunSrzI6Q55C+6Myn7VrJDzpHvEW8V
XxzJWE+dMwh3UKgoO+BmFVGSvbMcUQt0WBAeOvalMAcrQEbWOSESJ+3v0lKFlpw0
VRwmtwUB1rw+Web8b10Q62uIzT+qxbPufxEyBswNzVbPWtYOzoq6+wxp88ScfV6G
Z6p6CeIQ3DMfLx7E4pS0UCrK9LM60jlGRigwDgknEyO7gh+L9cJM7/Yu8YfuZiwq
wXAd5WZoni2I2rRtpvB4J4jN8zGY2eJ1qf6rxJepiEXh/XQcEgBtaudhFa/Z9UIy
D58SY5/u1TvyxUY2AseNmrnoFJF1U60RY1IrOHd70NHV1oZaTJXPgriQQ8xeqw5T
Bq7AeUSXcqXOvLavXdTVbGDDyspEWoFv6N3Onnk/TvtOTRDHOw2Tz3vK5fTlPmY7
n2eux9jKRnyBqMhKhnAIq7zLPDwCnWNUO9to0zSiHpQ8MfokLFQwmVfaWLyC86bx
qQTG2J8m7qfoq0csKocDpMfQSrXeEQyd9S8ZFWCCRx4bId54y9wa7gHrxYAy5Xb1
O/ycxByARy8of93ztzhURchjFS6kda1MAZRmudj/2zSCjbUQmUjPHEkzSfl1uqvU
VJ/FszQJeKxqVJdDS4eGEOXPjpXI+0f6JORqvE/ppGVT3Y8K0iG2ohgxTle/UJ9x
0IfajPXhOnd8Zk32iRV+bMuTzHLGUTGdIX++dIz1fmOMpDiz0mMGwp4gwL1tF3SW
VE/5W3l8Yzou01zhh+sJId5Sw90k0XWJLUyF9S39dgIRkEHGRAr/Gm6tuBDVo5xv
1qng0QyxBIdjyAsNC8q5fbiXDIXdLnXEJII4+h8kPsUEocT6I6sOHhMxMzX+CIaG
o9cK9F+LoezfNtFnG3TCKpf8UtL/6S8kpuu4lzLuEnjbIxPIMJTTDw2Xi8CW7+rM
HfPtw42YKjdsQBWQAWp0+Wahw4U07mxgCfjDIlVLtu7N/PdKIQZrpBTpcZPV/14i
hTBG3Ae2iIQoRIFOuY+HGLsRiLezdURfvONs8PXs5bxDtHFoD/rm4dI2koTF2IbJ
suCJ7YJaYe1xVSEyZxA6HIzebF3r6UaQKHneE8EEFTKP0axONwe32PIwfSUmpGF4
oJjrLF92skryy9esKOSDSEZWw9UnVCUOX9Y8MgXVMTGkeKHOkxblxjU/UPX5Exxy
zbVZbWA80Uug0hK3ecVflBV2OOmFp+7TrcwitoiRCaKI4VVr1Qxv8d6HlLakvmsN
sjgNbA4JIh35Nsr9AmQlCy05OuPYpkSlo+SlhWEZ2kkW3rvqe4DjV37A2G0mI4HL
eyqAspkzI8JocWBCE9gcZwXEbdfdTCVVqU7qIud9DtklHehHQrcOM/vjvWNsc+sa
pMafXVqBaDLDOmG0Qrl2cooNJUwwP3Pav69Wzv5EehXPLAujD84jd1hOWyPkgupW
PzVFD+tNLEqS0WNdZW3boVvlmAdEaNRPz0u5Yywus/xUYteaeL1Xvsas5trEIzsG
0mmLX1r99hBJSoH2GR6NH+cOmG9Ds1IaGOEt2ndmA46s8PUFGJghl3tA0/W7OnSQ
bo1RTJVYbxLt2L/Fx5kChUHnEYX53oyadTTbQub5+pb2O7ptcvWpchGosF1GNlj5
CBHfGy4EsUo582veVAuBABz90AX0etlmjEuSCKOHnysOoR6F1B5pRDss+n43YcZJ
qj2djnqbypjAkeky1M7lR5DKk7ddGX7rnbw/OO9k0GkOPYH98EFdq8nYn3bqLHOj
SLpACmTR72VNg2nFEdq2D61efHgj0kYD/L1bd+1p2vsUdsbzncoDA8ny/c0pRimL
AuQRIQxBSbmohiHv1s5P0aiPQFwfAnJQ2UfvJHkdfiHMzP9UAY+qQi4ujCgReCX9
1ckedXNnkz4IJqCeu04sBtBOTc93iOCpzXHxIu84gkK6bc/4weB+Zo25ooDV9dQ0
2BFDQRI6x0CADYOUoTglbmWSYrcoKTiuj6mgszoJ0ELED161u4xdt8Uz1k98EngW
Pi8uySscMmWVYCUWAsJQWrxv3LvRIOkL6gw6bGOoZcbs5/gPNWxxbOS3C9bFPjjY
BsbAEkamADCWTRTziu245Ua7i2H8GX67A7KDcr1p9V3Y6o5/o+qHKMa2i7Zxg5Jv
ZUPnt6+DHuSgQ1w2yXeq8j6R5eWeZevgkwN/b8gofeGiqOxSiz2mtKCcMVtpb12j
tUIcyX5t1BrW2ofgZUi0f5dX4PRD5eqYVHzqELSKvKcRc+wkuWB1Oobbr52APX/h
ev+pCHnZred0UuayvnGEc5tPpD4hTFE6avJL6ca5TeFKnFGXuQitareX+QY01qv4
5p5jjrn893FrW9J4OTou9pLidWrH1hZ8GdlZ7xplLbt+Y4nqhTr3171FVAOsL7Ph
DPYKpfAJ1QlOSLbcpoYmtiAkK646ahPyBCKBODB1LgWXcCMLkN8pwIFpGnoySAZZ
XbXm1a9vJlAM3Ja6xq7kzQgZe77rfDYkyuNnSilqvjLKVLptOROn54NCUTwKhAGT
mzKHNBKCa5OBCnzAo2yOmBgQeJYFkZ8/QZwVLKgV5YPq8dlEHFXvgs+MND0o2UCa
a0hfgnOQErwX0HEJu4KSO8YsjAPJaQ+55uzwcaxnN8/zHqr7XP6+AsQjRgwTczgA
CnRMYfuhOBUVSz4za5DYECGH/YQkZ9U3uB0kY2z0q/M5Ib5ptHJyNW8bVbBmiJRv
5vqp+Kkwc8SkOyDuj+QLC1/kecb7mCFE/ULHtebgd7suTQ7+uq0zun3eahHpBqVY
TNzgYEBcUUAt+3OVmGnP4uA998jFcXJ0nKF6IJhRPC5XCz0QIM7d3APW5snV+7Rf
gnyvZaPCELEeRgy0p+sWXDR2KNwmSCjYTRLHrM3oFgeWcOzSUpBx8g2k6IECEAPI
2viAOlfSFTHVLrmstLgO/1iUv1FC7RPvmVAkkO6wgQPZiyGnztTJwaIAM31JBMow
gNj4OLVQV9fRtiMPW8q0Urv2DscP/euOo2Nc9Vfygv6YSKavV3S8LxtaFzW8BPbc
YBK3IJYIBGwyUt3QekBT8vyjm/CBY4zooB8F4NmD7cXHq6tfI8LSZha7n+X9+jj8
oYKJNBEs0hpParH/Zk1efrWRevfKm3DQIuEEn7/fT0PdEUUYKpoqiU5kS1a+/3+Z
W6sHJL2dNeTMBISkSeEdKu26Eq7WjVrvUmJugu/mVBcSfbm8BfvxfaMrQvzOR4dq
o+++Z5clB+xxHQyQGCMF2ap4U4IGmJ+TH9/3FhzKRJZgZwe7oDZ+JSj41tBZ8Emm
gGXW2lA613H0KRmemPrR48GVI93C/yliOghlMMB1R+EglQ3DJA4bxQFi1tJKpMAw
i82HCG33uUCt5XWcjsCDiIBxWM2deVSbPgY/x1HZcTMxWoiRoNVuvnRH9cEPHSm5
SvoJZy99OP2538K4+OGwgchhFT/Y+6jyNEOS/r5yT6LeYBUzYVQXP4W0DS1p9l/e
yI1dk5YSGyLeUTEVbIpPrp01exZfxpEQU9Nvx8rD3HXrsHXiWXwMEWHe6fYqybEn
zjoWuk9FoCB6V387AF/t1zoK/CURBF4W7NWk7KZn61HVyQVGngt0B07eS447cqIz
wV5y7xyALvKF/i+JRIKDcBdElPz3m2bSKi5AiXQxG7ND7VDl5My8nopwbOPg0Z+C
9LvG2/rlFNrIW70ujOA876GGkmoC2shWTqmOibS7ApI/BBP3OmkmQAUCblzmaC/X
0cz6WOwGZoEj6JlHQ1CKq1V7FB7Kd0G7tSPFb5MM1nHuQwv5y95MHpsyaWxqMiUW
XBmdLpGyVFUz6EAehpBS9sQ9S4+vQZ4yQleuUKc6wIjZvNyhldZfYlXPA8dvX8Ku
3xYhdtLDItIpmwdNjjH8DqJVLUCLeqr7LZHdKFqzyUY3KWGk4df+cI9FWdSNQ3AJ
At0eZWJBv3qDXr94+WQOyGjgEwYuy57GBX/wHG1Nd4DprHCi2l6LLSIiZr/u2eQw
Bl0M9hKSNmuCXpt99Cqxhln9DJL/T9Db1Ytcq/xPGLyTbRUJ5CA5zmYcBOcc5+x4
kWPU/3zIwAhSfVByeCqLsQACax8fmZfE3vUqPgJNfbz+g4R0Asjtshy8cVj2Z4l1
UGb6D2r+hAyaheyxmCUHRiyCAVeMAHosL6ABAAAbh2/gbwwmjODYDCheO29HIAVI
sPnxhGTACdid5gjCAxF58WrDbVNo+V7yfu1OuKkJDGAsKYZIxuEjCXr0lCHQI+cL
H56/AmrWU0l5kFp4X5xkq5ssWcdFjyItf9iJmf3XLSTUQ4RqxYqPyaVxMvfmtHcq
fbrcHI/GPoTz9lvGwmBvwmS6sDMDQV3vOurPWGJapVHWR3gXjE8ME6NQoKnZYB70
d766BhAzQUBmXpFz+MJwhdMhHWXRtGqd6xdV0CdlIF4ruyI39uE5oBaCWtIT6soD
XVo/vq58fpkOM2cBU9VzcYvXeAwoo1X0wug0ynWKrbPYO7g9HP6EazPYCSOv5zH4
Klz6kA5Y2/vnzCeiwB+eqdWrd8uJuml343qheuZSTFQRxLuJy562IQpLRs3W0h4c
1aPmm7EruKqpXrBEwyG5wM8fEeixlvouYcaQ/7uJKieipI3JFexlJlPFsK9BK4ub
aeiruv6LZE7AvspkOKGhnVSAOW8J0I4wEyQGTFSlIfC+fWL2vhMR5owrdzmlp6me
dp7usnCesAT3rBTntHcNPj7PAXc4ajrgL4HHX71lL73mhjyZZQokBaO8WYmKXCJf
KCIAX46H5IAOfZFS4rTGHRL7OEXb3YT3SDXHiscWrT3OgO3UNYZHt6kgP7tZcBjL
z5HxbCf7J6IHSaCwbneFCcBOpsdh4KWRAQ+dtV+yE7zLziLqw6XHsfnCrQecnwj2
NL/Ic4M7Jv0/5rcAUCqf17WBeto5Rca7M1Og4se2uKqnDN5n9Y11TlYLPGuuMg+7
990l+pYxhVir8Z69cNkkGQD1iex+vIYHF4bY6NOasfEVQbzdEvGsVgDrAZWaFWhf
Rmx8CzNDmSRteXFMI/cWy2GC0b0giLg+fLGmk033nT+h/TAZ+/3y2YOpJkW4litg
oROY6iga6oUa98FzE89jhyZZN3znX2B08VIN1STx45jZMTMpnQd5yk5dWf62+eqI
P4SAFfatqFK2AgbLy7s3ly1NNq6p1B3tAmOI0gio+q1LN4hDtEcRVZWVPJpBrM31
HJSPGarHYc24AK0puDD1gNxIfC33v4VNZgEruFKFXh6RggHL3evsIH8UxVfRi6fl
QF2E7HMgajS2axPfwgECwR98DaDW/3wQ91+sFMaKa4AUWq2yrYoH/5bOKDNprfw6
x/4WYAv3+RgJ3sgb+p+Z9N/81fRsKIRGQ4TyfO7J82XzQ/uYx1ToqcDX1C0T3Rur
rCotldoYpvPWBkBe4nHchaNMGM2Wj8PtcWPZBqO/CZEbRasGwM7hN7BlbmZsD1X6
heeLHPOCG6fNwk9RX/I5kJjxYjs9ea5or+rB/soWZcWHWZUi2ACJGe7L7JpQe5f4
Yptblz+EoHLhCNuznIs0bf4NlNDCUrwZQFkx6Sh28iHmi4NOUSTsqljtJ/yfLMyK
wg5p/iiDV2gHZ3pDfcQRGpNI8bSFibQeKrmCW/Bxs3MS0J0TTUEu54cqmxMb0hEk
z869+VOlssuZ4FiXunQWkTgEC8s1CsXV/26imqONv43Ky/9FG9BDIluywKK03f7s
4B5c2pwiW6LUw6d+slbxs4hqqa5buF2+aOOzEKt7Tl6Tfbvux7d5QgU7Ezw/aCs9
DYsW0RTDoNPG8fFbtY/gL5q2s8Mt4WuK9gNui9TkyrW859wIfA8rZKWm1YfCQeOp
Z8sTbCu9tlzJJii1OWsnu74a3WguGhCf5RmJ4GRLiizzaOjfBk2tTLnz7BNn1lyg
m9DwZWqt8Or02UN3th8WC+dQJDbp2aSfRNR2VcD230Nb31NxHZGQnKvwfAwPWfmp
Uy5zHJ7xjGT4ySenL34vAfbrXGZ3PpOhsR1V5nfaSk7apdiB698TiOYku6QgH0nO
dxdHmsjwmLahwMBsmOuMlNFWJ29DtPS2OftiGHMDmsGZrOua07aTGjxcaZ1ijSZr
noXUGaKfioBKJoA1r3NVW8s0H6ss19RIRrnW2Y/ZoRu3JBk8nw3XKCGGY4Zm+kST
XWffub0c0aVbWauodHLKBdfO8EZx7tM8yH+hzgHbhgWuK3PNVXuy+2f4F5IArpyV
n9CL06c2ser7HADBoJFZxyc6crAgpS0P6Xg6+lH1XKazU1NjTTc9LuwPBhLe8KNz
q+e9o+hlZEMWq+s4F/ioBNBsFlzU7TldskIZyFyg1qJfROIjWmXmD01Y64QrxSRY
TD5a1M95QfRDaNk1+Y/06dbxKrAE+UfSQPo/sQtKDARdKVUo5EnTAdVdbwVtTnHu
9dHGj6mclYEPmyPf3O67SQC/cHnDnew2sFJgvGH00HO5AOizoz8QWPcHEkVE8QPA
XHSUBiwsEzg+d9TdD54PEE/NHXADONEbpI9ytFuj4zibjijmORtAIgLK6BpnZLZg
s4M8gRUgYaI1joZk2zv6FPQHgh2A7wMMmGxMAp8EskfDGh5Ay3pVa4iWStbzTIZQ
BhoLHgVWYkClP4o3oMZl6vqUeYh4f1bDvsaW4dNYBZjgMCQdMxjov3s/7FNY84Iu
enBpFIXMWsCKghs7qALPpmF0eJQdEVpWn/829+f6rx7kzceMVhjOZCKhG4MqMqrA
ByRVUwanjDPt333A9+zwvvkaoUvfZVI+D9TVIVWZs8HDEhlq07VB8TjIpdb1XMOQ
E6XHmnAj52Jw/nzeBDLbB044NLzPdHuqqbTGqr/YfVWmCfN1JSJ0AAifKEAVRqNY
nHTUo9ItvIBUKmk1hY5P3p7DzIxzTYQMTpNsF9kceRV8YafSdXBQCymo/qCtxdVD
EQPkoyLv/Dv0D2L+U4iXMY6uYqWbV4ytasrLbCrVCQp1UsiSjaT/sdbPItfhpm5e
T3v31nzZaRnEVHYdDdcu3QqGfX5kPwWY9wqHJcLob18KIGQltR9lYTjjjWyuceNX
MWTbGoWfMCv+pTESB5FHAdiyIu9wLM2AdDTIlhm/mXuflhO4xm06IbvygFMaBCb6
nHq0nU6Urw5EcPSaCX3wPpJXRdGi0BXM2EjXWRTsbXatvZ6lTL68JpxcsEQa9PBc
ktTwcLyc7w7TQ0/T3WOWodphLqscBgcJutCMZUDaMB+mQ+sqzubRJihxuy468AJM
NTwUJXRVRQuN9b5bKpdZBafY99aaZqgnohlgiVIKoiHnpLpibxK+gGNx/XuH89Os
GzcqCXIiG1rJluzFsyXYTi0rbiEDnGXphWAhiCUsoB5YrwawaZEoyy0O1Tl25JQX
my8HyA9Hu01FaaJLGs9IoE49NaMQl//5YCm8CIX93B3RhsgPASofhzZsR9DYwY/e
Nb5GObE3U/pSvIyYvim8Pmt8whVBFAQSUZt9z3jC0AWCCMlAlRddhI3A2FDBgRAh
0WnqzFAWDcLLaggFel1WH9YdcK3TOhefV0OE4FQKL7xIRhkksVuuHgXz/IASD9yM
5TU6g4dVVPwhp8DlD8R1nb/a0eDz3s+YPbQA3OYAaIVHMnzfntrfjla5DPxG3wU+
X2CtUgbK9g1S9XQfrJTMUbPgZM7hra6OyWWRmHyb+CTL/q70A7cm8gHSUtUNGdmZ
wAiU9P6urYynlD+zmCyuik50D5MEHZqVUFGYuI10rZ0ZI+fGUy7hE6NSTFRJlm/u
aGbDdmru9CPISkhTQGTolJbGvCoF4t52Ws5NxGj6ECwMilPxCNRSReDaEs1ZU4AM
xwC3VQ5jwjnRChlXdAeNFvVBXnnN6ZoQTsfB93X6IA2J3XnM+JR+jGp99pD/fTNJ
6F9rNcaTsdIreQnHgzPcMccZhaPXR6la6zLSNyAKXNrymVQ220P3Jx52aO266mAm
w07wRT8RmZcutoSuJSN2w/menx+hbDmuUFsbKyCdCwLnioAIAEgA/zHzJZXDC0+4
vTendtAfz9ihJXuslHXtoMn+Jkp9Eq+XwSav61YSMKwNv4gOEXR9kRWENH5rc36X
8IIfzg9BfAtUBeSzgbM/ezAA7mNEq+6JTy3ZWUCp6LNNqSPc181PnhtrDqhdrUSn
xHNKUSKSohzsc4CdMyrp059FYDNJUOkgej81Ytr9tzYyOftY/qEVt7vwmR3yHdbp
X+Kp6Z2V3r0CQOMSZC67SGPUnAiqkMAb35JEbe8DNeTt+9l3i+LbkExIehAFkYox
q+UxKcIBqTPgK6wYAJRufgFdBJ8MbimdOKSiCP4/8FHHBT1GVv8hCXdFvxcrq13u
xA79ojCZkNZakbO4PXl1h7TFMd9WCgPu+NgQ7yeDydo3U4ia80CbjCV3DENoPxiJ
fFgnR09Pf0rMPm7V25i4p5zVHb3KsV/yYfzkeep8B0xH9fAm6W52Iwz8pP/4d8f9
ljVY+0zyvyBLsstw05W0NLpgO3SZWdwkD/gCamQQ7x1M2Nu5FjQIQfoJ8+CMc7U5
clBOBTzctSVZXCefA/rQ2DtGH5A2nuzJ27EtAsH9Mh67fDZXL+k0BG5kPTgBRE7/
GOBsv68X+BDGPej0SJFCEoeawXBfjI7TTu25a4AflW+RF+RQeTR/yYuA+UoaS2fU
HxzcZmrZPQBKsrhiSaP64fukFjWfM7txxTk8xqGxBaK5hwaA4YGn4tw+Pt4RexeP
/wuubSRoxU/XjvY4xX+ytutDxXJCWlNi9vjoZvnN7i3Ca7axWu9w4ruztYg2wwsS
oXs8UIMISDHJvI7rW3JtCHFy2yzqY+MkXUjMXHVuiQerfhVaTi0DpjLYNvON7nXk
6+1C5ZiRAV7ppSOdsVY8zixwODdAvGEciwKbLWp2Ytf2+4nG3x18kGkjnw95QLF0
V6wSKvJCSCWtqHPXJk23MNbX/lkHBIWJ1Fsm5EGEsCv47jmOWpA53d8tb8Y+Cj3D
1HBR/yk9QaMxR1HAPS1CSI034/062XtVObsA3Qx4piN9g+pIjUqNRv2ZU6gSq1jO
GqhdmmFHGIPB80j+BhrOA+hXsk/WuApABqWVltmNrB5HwK7PGlFDvBqD3dAoVuj1
+VjKCn81kDccTl1gp0e2VN6UbhdT3+HvlBlRy48Iz1f2rz/6VGGajND1W0mD2lbA
CRUACdpHG5UF9sdnOOis9J5HGg28DwHvcmDYGWxRekfFxvR9nwZovbw1+ufI/TnT
+mqwIg88fwCGmi9EEgSNVwJpoYLq3K7YXF7gL0uQ+vhplsBynvmL7OzQtSi5KBBX
NAgDb0z6lb81oNtikm7LeR4R0cR6tQ2AiaK63Ps+g9Skif3Nj5ejlO9DVFSx4b9D
L957Qib8816+FtBGceG3ofNcOyIJmSAjQEx653CGM3XzEqTpYy2rQqZBp6rIMz6m
qefWcRXezyAgtKf6NlAdTcUcJnvI+9hWMz1XXcXQRLLasALkBB266DV3C4YrKlFO
KsIFRr4CC3Nq7m1TZuWqkW0itfyXzrmdR6MzCQaNzEICOdVCWcS441kUW8HmZtKY
aWI+qYDsk9imFaK+yiAObu+8orTZYQGZWt7928CZgLFAFALUPIQBVIDspnQ+LBik
95ih7NDLcfn/DQYx5uDACS7vKM7q2zmBKxPUuXgALA/sBpmVsetkwl0XniTGzDk7
aISrWZZXK/xGmuk7KDUtIWwfy5pDBk7jo7aCp02B/lXNmXjv898edH6OaxGjbFrx
cn/sqvpQnajVKIqJXvJrOAxv051wRNpTy+D3HiPv2ZwRkzMXcmOJXAPlbvdEvonv
nDjtOU2Th0w1XswupXaO1HQbGm4Q0UhlpICKoKHZEIqNOSkMPtb7vx814C/dXW9r
3tdXhbP//wJO7VBWTT414LptYa5mOZqbs7neAMZdlU3+2y7mafV0QoZ+Q94BXzuZ
2D7h7110bLbhTwmeVUZIFWvTum+MZuCr9Xh0IxK/EJA3pSNQi1GuxD5BcyE8nzl7
H43614rs3Zh5saXHo7WYw6rchePASy5p4L+dM9oCIMYa321XtCe5PqRv7rzaPF3b
2nU74dojO8MZBPOXGM6r51+6oKj9+QsLGJZdgSKEu7In2gStCad0Ed+sVxF1RtN2
3no5daRgiRpz955iwNGWFFxEhqmqKEAjDH+C7r6a4txiNYDsHxQYRZf8KxyPHSPU
r8i7545LiudWCQB1nSgF6Wvi4yA/57oSR7Ic3chYuT2DPrgWZFHFf4mLAkYgHJEL
zDlIKS7qEwqt4YyxF1R9eiOud6+8Guf2ICGLLXNN+Xh9HnFTr43S+xzQcQmNkwyj
HpPWOr0iasQk9/q4WS2hQMb5+IXlMgil74DlMsYzF/krHWdDOYaJZETUmJcjPHof
75Jc3Oqn8ILllJ989CJOprLfWfcbYSmDQzFQTrb6ZdDPsv7bzdBrm1rkkj1+g7/g
fO+t2qRaKG76hGAO0lNvcCxAFHEyA3YuB3RtELM7mvpI8+nGJd1vlYYZKg+LDJ82
krWbCHLcFu9y5oy9iZNp3mTALkBQmv5nuZwAuo0+mvdReXryl12PN2gFQeExAQNJ
QcuKduhkVArDubzu6Yg7ZRwJMKoVAY5sbA2glOfbhMg4y4MApf+qhsV7FBh2BHbH
NhmbumZy5UFwrZUMl+9CpopaQUlhM2AWXPUxWVu524lsendBIltAI0a2uqTkh+ly
dRvz+ErNq4ejPCXH5z4GFdsTVuV9+YkGrskNDFtBnTe5fjxyQl0m1GHF264CwFLq
WMln59g4cqNN+ZJ/YFJGJ0+ypUEaj4Jv1lKQ0zRfkgm5bGqMtUVmonC3pjY42NUz
+VsjLHsTXriIWg1l5epsyBeoZwfKwkLd68Zy5FF1OzOrexz1j8wPGsnAEU7DHJ4n
wWuzTP4vFbGURzkXX2c8H9MIu5enD7A6ofMvut+NAy3iI/QShViMoDpTOuAWF+51
Dc9Yqi8+o1511l1xEp7Tsg9ELWN5wHz3T0ibhvpgCIHAoxXVkiqCzDRjro/bIG07
q5Per8pGlVt662JuOtOHIZDYHgxp06zSNSs72tnnXb1L+578p/z5BtkqgQmFGc/O
8OmNFrtJIVv1JD0xeNk/UgPCqZuILp3nUVH0iDTgFRS4wtMnJ0nUUkqeeOwy1EmA
ZLcsCb2XnjJuc1Tb202bgrQGI7p2LuFgz0Cutbm49+udtDTSA0N2LJP4XrNNiDvs
0tE+0Zo7KUQRDMfWqDvL6GpoE5NL49obiq5SxEZ3ZWuV6C8IOKmW+/pAeUt4cQ1M
O0XoGO+2Oi+dp8xKMotGEbIIIVx30Nw0mCidog8HPMpie0J+jCY8+fVbYDRrq4A4
FqwUEvDIXxtGEHB2rqU/2tXNNpDhJbhHXNu0RmuAvPnV5V7fCcX/EZtcAcxL/rti
QxE8Ip34rHAofK2+3Xju/Am15xa4h60ZfYk08n/lOcdoEhwsXg+r65im0KscCRn8
5/A+xEDhGE9sur4UllRSSUDpG3Da4c6makGTBSugbM0c6gYNi6jFCEADz28PVTAM
/yJmPWXrwSt92cT02iWY4wWDTwjEmOnvDRTXy/4kBZyu5DHsNjuvLDZCqP3qaLQb
RMyw56ii6TiBOBOWtyW7xzxyKoWoUH0aIPqoe+eScVnHJaLoxIw5EhY1sbfRfz3v
4QlnRpiMrAnkdjBNA4miYGQ3PGjwE5HER1YizeO6u4eAGGem7xgOACibS4cfco7/
NFl6m1/P38aZKKnq2EOcPlpwXKfyBHI2191v8AmELv6nAeDsRtaC26J49FJ14x7H
1Q0gjiS0GJvffBKVunzPibZwDp7O/Qnc2Kzys+6PIkB9BJwf75M75zNj9H8ggJpb
SapKW2E7YuBAHu6iVqYippbXsQrONYaz9+hXUrOkbfINm7qFtzXIhwJEFI3JikFn
LmujpVJxEJ527KhTUV9n26mGhO6NsGwxjNKs6JDWvnsZgs965pI/chxTrn27FwPA
RD7hHd4uxrxjVNf5srMgS0REBvqv4j+abipEYp67K+0HK0fSfvSKweNGBBcdl2z6
41uqCWrsyfEpdWq889NXMyRvQMhwrjNUKk8DUzvwC2GF3K1t0Mtc3YCM/WYMx2/N
k2Ac41Hs9Syy/V9TSUVVY377IXBCSY7LIxazV7YI+eRyyDLvSXFjoIqKFtdah8Zt
OXaQZo1AU4tiwCjtBJvJn+m+sZj5FpV98hLqT3yawiASqRUCr2LsE1IfD3g6w+fx
aoRuoN0bL6go7RVcMbPcV5cAf8wlGUBHpSPOpA/wEgTQhS0gWSVIN2wA5rSPrbft
TAREQeNeLqI4Mv7j0tC1GLdrAvYKgJC0ILCCPb7U2t/zQsXVqxR2oP4FZaLKgkh1
bKPeycjlJtjfwj/yjqH7lsckAwhxrL51GW4IIujPaoEfwhCSTszpx3EOt9wU0EQU
j27D0dupUvd8Pkkc3+zQyZCfhLthlxMOCCcs/lP+8QWxoZpoMRGPsO2VcraPZNmX
O7RU8MkRRehSxhfNwXV0SJX+34e4MYt/NmfkaQ6JJYbmetT0SNpRmyim60eXiuo4
Pn1dJuDUIoLuue2U5OQVOnNt8M/JAPPm8HdDzOtM2Io9nnWwpkbkprWHQoXP0WUj
wZZzEd5qPxWEg6Dp2wuT8Xhbjn7uZFOKTF8uhcasI7YBCxm+lm/YEu+4rWcs8zjB
Zhfgk63d/S4Y6pZ96PioRe65fnvCtfTu5pNk873/NfaKe40Dy905ou4IIFn+PWS2
maHxHLpFL/iiXfvW8MJ4tF5mwLmMlhh0iyK2EpOZuusjv6qY22BxTIW9OuU6n4/q
ccgt1fKDiOgceEFKgkMvnfIrkmcS0pHSG0QDb47K4413XDcsfFoxWP2oUNEwEptG
2NeTzkLXK+rtx/Dg4mhOCypSAfsYFcj5vzfnakE5whUZQxCsOJXnXbs4hGsshZV2
ma/QpvUXlJvaWfpe8o0vEpfFPSfZaG0ge2DtwhNz1ACwrhXYAng1gHAxUtAGJDy5
oGNoABFYOidh4NAOJ1UBBhj/Bsbp1LwPBWSqz2gpoq09XtcfINuZLZjwReF1VrMh
mVsYIv+HKiF1q0BjgWpKDYfJy4nmu85UTgopEpmpSkHMWCrNncm7TJnfV3PLyJh1
6mQWNTUPJ+ENygclN3KVeCe1fj5owJ9CRHYj+Uyxo3r/qNpURYaq5RUAtrpKN1xT
XxrxnH38MRLIMxQi0y5t5VaWTUMdW3ZUMBzhcBBueoWAlOC0d11sDgHrPD1pCCZZ
RSpXPQ+ISMepSg+6Up4nY88s7TfwVhqGZx65czxoFa2qlZ42owKevoJJ/Jokr5m9
aOvHHoVGMDIgkQIN4iVHwcZ4xBD7NHQissU7uZfUA+ieaB+/T1Xe9F/bKfg6akK9
ti9b4s/Ovhx5UwCQyLV7RZ+lV9SYNHGlQu3FSwCX7n5Ns2nAr/rDWEJ6TFaMYViu
84d6Omp6L61oIlJoQ7WeXD8ZA/+KCi9sdNwE6qfa02u8x4K8N4oKght1dTKw6uad
p0N0AGoZ/4dJjKh05GU4X/wMs+dRo9QRF9dmMA6cEr87XCOrfTczvqX3dcYWcZLh
jI6UyGCdNn7qEYrHT72j8uSnzJykgKDbEdxe0dFrgl7AF/NeB67zV21Atmd6jzUj
uX16ExdBvD1+JzVveaDknUxqFuJpCdGf5Gm8hAZfGjp69ZRsyhjFFZkC26VTqsrK
LM1Wc5Ut7eYmnfH9bpaRLfCqz5Mq5eNQ5Ni0lXWwMZ4wTpTwzkLONC386y6XW2Mt
VOeeutCGJSowwAHz/xS+1pTFvrgS8QJaXxw3OB9d880Y9BW9oBP9azXBMQq8f6Yb
2UA4GvW7/Aeljj3GWw3YVfSy+CrTqnw0ZV2echqashGF9LKHdhar7VXHbpdnmUyu
MYv7jAUo39G+Yqr/IKYKXLO4pZc++sZsmY/OfUfv1Kmw352MuiGfE2GwRif+PYUw
7/6d1tlxidyno2FN/ZaiAM88x7E4QJg2I1nPpXdeH/rtx3hslgBDA6dx7+I+oXeY
OPJv3o4WfRRQA/za4/TrOf9XOho/s6U8wzIKAU7f/lR8jLJLCxvi6R3UR+sgn4hJ
X5HUAuXy1TAEb7IvU58aQBHAKVeYQ/EKpabJQ1NexPjaYhujSfH0GLmAL1A6ZBfa
3pj+NB54S0TBpqgIEOrWOIKEq+sw0YZzMW9CqnGCJ1OTqJcRjOSjoelDKYAOIATs
Xfj1viRjVJ+EBUSOQPuF5c6kdNUvSRgLwianZiJqiynYIRbybhVAq/jbECdeVhKs
1XK0YSKnvVZp7huPMznyXS8KkAMKpiZFC1VErQjY0smGlg1l6LLsai40eEKiHE3Q
LaF7Om30nH0kVPUizhpWiL3+01ij1JaTpHjgkfKZx2GDynOALhPs+OWMPGVb9u0+
iHv76i2ex59b2ORg1qO9qrCewESS6FoOUNl04qmqqjeNNVoOqU8DtSq+nhfDL5iO
GXbJ4Q423ijQUvYnSngZ1QhZye1zhfE4eDBe+BOvntShCVeu7gR//lIwDtECewGh
mo3mwLmIdUqW7EA/QHlpz7EStiI6+B4UCCQf9LhREnbb+7khdY7tfm90D/5r1JOk
2apH9cme2tfy9WuNjuO46WBd+8b3ceDLT1CpVJPf89oabSYFm72eGDOovVGfn0tZ
2q+IUflLx4eWHqOQOuCnKseTYOVoOAbnwWFwQOsHcHHla2c5UO/f7LEESibZYVM/
2vq/w7rXa520suDmxWtMJ5ryNpPZbXiC7XceBEmrYBH8/5gQVjXX/f/DEidqctIy
L+BueKNM2dXl8/GpaT9dB7oRFKuBu3dSe4V9HB3lHCnY7Ku/UtPWKCKPlsMo7pb6
F7izitN9d5a9LMbXOTNV0NKGMpEA1ejLgYo50mY6BcG3g+/TpSkHCgNrlrPMWFOo
Vn1vk7O5ULVhcXlNAJP6aDdtac4OgIZZE5R0weIwL49JIui3LOoGWzepMe5Pu3Pl
GudIUNpD/sp2PiwNgNqI1VBbkNl0os2iCMicfrk4V4STlsWSkRLTUfAaRR8X7WJV
xFmF/bR6c5K2ldmeIiLxlZwnx4bq6wIE+cgkXojw7mGjLv3hq24uFyeWOynm3qEX
uxMjkeeMFfy9lgrhpCWIJg9TB1gwWxABHuCvYEjfVBRjp8dszT/bWB9HX8803nZ/
r5MrqKk3X6f0EV1U795use4DTvT7wHdJYYIdo3JQpiR0DYb3EN8Xowdp12ikpMFd
R+pgW4vxliGSm05ii8jg78aUzymq56F3rXUMZJe+QFODP8jmF6T+1F+rskWyVF/K
Ix0+PyX5E21K37Ul0Ix7Wlf9NmH9+ig04KoVB5F9hzws9fXSlFWJbhzRlR77bdpZ
tN/sHglLTOElFATWf4hfF+YKtjWY56Y3oHViw1A9z3zSQwKhegR0LYeEIxGqn7PR
8aHS/ygfCJp+BTLu5cQyRy/9KnQizprQxcTMWboAyDWAPACdHpB+JPzUXW2BW4zB
2dI1ho96NcpEfHYEzWTrYCz0MEMlSZ+CcTGTmr0c+eLFRyMy3Ot+/N35WmaJl9KZ
3+V81Js1ZEmmOp6XstaLcJbaMY8sCHqrgwdgGbM47VYIUk1cedHM5YlXY7iETAQQ
jzfZdd1hIkSgEDrGku5LTtLe+fhbVZONRPuRXevp+PeOXr4DOaQxyPGGv6L64iXo
Y6DP7d0BrI3Mntqa6Pma2c5VofcmOjeH7wDI9FgnMD80itD5U0Zsne1f+qQMJDD8
0er6BCDtInqHnAuvPihxQqODgD3NPLiQWizQwnlyAqb/R4x53KDvCE0/wIWtnYPZ
PATFQ2YZwcNFAUiaYDe6OSWl0OmUdrfQ/XnLvKdD5PKwR3/chmGs08bS8nW6mVeH
rI9LXSjMRDnfdIHoTOOAp14OvnrCA/Zilozr6Dvhj9miu5VOi8NcLJbD7hoabX4e
VIsdgv0AbhY5MWE7koBjTNjO/czD/ObyBPU0XETic1a5RLGODLGwdabdqmjXpBc8
VCRRyWQq0JsUYWvwGwABqenaeVsBBoJvKuonJwVsjpT8Qlw/9u0SmzJSr+xCOOy9
3Z506MnZe1OCXaQ1S03JcPqlHYUuFgCUA6qzznnHcj3QdCj9Nbi+XLHnPZ4ZhVcG
IlUG6K3p7n2UaIdeSh5p6eWxKtnDBySnrLkYemo2mH0qD6nSL2EtWQWafOtFD2AG
I3IASZOb4WMRg3Oo2sjS0OYa2p8yV8BFlqpbyW7DKjghUydtgP7c7hht3FsNeS9c
I6kka4vk6eKmJkdMn33bc/lqRyEBZZBUpMLSwEBGOh9+WSoXHhIeuy767OaQtkUA
c12T56sMURtvcyrJdvNVWFKxJXbRAPdEtzfwZRAxbigwNdtcAKlreJ+p3fCrZjB3
dgLeYk3gBKRQzd4lF0YIVeeZpGwI3ynoH8J3PyvhHFKUPg7kS0f2Teeux+IJ4c7m
c59Zevo/KSHY3Hn3LlNHpPS1szm1gqCU/BjA3g3gKZJJ/gK43j+JDH8u44nMEV9Z
XjkdvCj3aB80UuHsIDu7c0cdC688r61H0RlsZ0+f1y/Npadq5o9wsrXcE7QML6Mv
45znzwj+fOtSuyJpF1aZ9/WRUMpX1g3j5vHEWXsTGd+hS9t8U0XTZZZ9Z9m6B3sg
u1JLjcdYQUAwIj7Ih1TrK07nRzrvRsWn+V3fvQoF8hew0r0F7ioOW8apU8YUlJDu
HVPoFsCWVzswyBlsdWQ3T6awsEPIBkOGs9yUg+lzVUL1pThe6FlBQcme8LhBkkup
12eqO6RNL0r3mvX4KY0XEn0S1ObdYtCycQUG6Bix3Q1RmToS21Eu1CatZfPFwe5H
e5JlX279Oa8OpER4CzxAdPLjEnFjWlxKJ75e/R5prJzdutpvIgacBTN1EbUkIdTZ
m3dP6uEyC3tI+A+50UKgI3sDDEg+sqiYaMIPJE1ZhrhasZo5VSqJrEAQwbnNQD89
xaE3RcMAEyWVY8m8KK7gKiJa9DKJjnnrtpnDIkurg40v3x5EA7i/o0Z4xSL0xMk5
LTTljttfjA4TXcXXjoHoOqXqxu5H37a594MHOTdNozuZZZB1F3BPJ/GslNHvWjSV
p6tayQpgoMf9pWelvKuX6j+t88wEaYtAkZ05fr6zIa1kHkwtYnsxYxEzpXCk8YiZ
cnpVZvS8BajyBeJP1a01Y3CIdQNdRTM316VepC7iOJ4oSM9N8NfQSZ6dqa8EzuNM
RwfvychwWebDbOXjgtaVnEdQtCDBW4/c7SP87jEyEexnUwdyBNFNOshTGa1zKwzp
XMYtctmdnh4neQGbxA1yLjG1sB31WmCzVNGOoycP3zf035h2PT5BKMYFVPDi0L+v
70xUr7QW9q65OMR+IjgawNfBpM+DI3rK1sJXTJ+WUUV27DaJgyARyQFStoecWUZI
VpFJjiV9DRnFY5B/l3z3KAOK+tuG+AyyBiO3H5/gJOxc57VCBPbmlTFRxP/joPOX
Q9KhB0KfuXmu+KPUH8mXYAHIod/gVlZ1IJZAvLNdzLWmmNHNWEbw2DvMdTQ9KqxN
Iiq9CEhC6oHcQsrV6FdM18dPATNTA2Hjvhm3TTpd1q7sBcEV9Uu2jcsgFt0cme9J
Fk70BkWnKUKci0a6Zmp3Uy+HGdDSrYAQ2WmbK301sv7dIiW972CErXh2Kz/mUvpr
gl8qrjs2VH3EQTwboo1umoaEeI5ZQzYQblm5WA9ppHU5gKIrpEl5xI8F8WdpKMo/
ybnJ38TGl8ip1CkW/Up9RBE3vb6rGjsuQK0o6z2GH0qriWWJ2PpelyDZ0nFDmL4P
wPFQVIhEj83EDNSPnLfP8gm5htCc7Nauehth0ZY1HXdGgFRdvj948HN0oGhtEM+N
iAmz08sq6WgbjaxP7CDp1UMb1UNwM+wKhPIUdbNj4Mu7rGPATc85dkFNhN5Rhf7i
vPaMHjcNL21EpurBZ8PQyd3lG5P1Ds/qxFUyrr3/Gu6YRRWiztJJz38ByuNQWzug
zfX0TsHm0ZGLqujPtBKJpQ/QsVsTzEM8bs/So09JHbq6MY1n8enqYLp8FiTCtO6l
XueBzYEP2Jfr2ocbCUAMNGoB9QRDP9C1CGO9y0lGu8wKdIPEipb8UUfnQ75eIyTw
C9Vceiwy7vWjfKFpoKcjNFg4nK2wmhRTowpwCnOkuEHPVrbZbB0mdqqZWThtsWh6
rXm1MdiSX0L8o09wMn+63OSvs00DBlTFEB5/IlZYX9V0hRBXb8zMxSe9GeM55dvR
k1uYOcum9I9RBexH/nxsr7QC94vcfeJlzPfrIhi22AJsTp4GMy8L+eY5bCr8B78H
ju0qKixbMt50Qz2xtNG24rxtjcnaarjsHhhkT1NbDnOiLKlQR8Z7d37T9/icjtW4
o31R7GH/DJ7Wmk+1Slic5GSKKZ5Zy0o3N/+mRmkQE/WAlhW4s2tJMNdUQQrZ1ca9
rdBBHLuZOqB8wV8WPvoCVMfFsYWlC2f5BshWPmdiHFoxnDQgOMrCBRhWhv9D/fzl
2eeZzLVtg7Xt9TyUFUMjUUJVYoecjh2VsR1VucHW6w18FFBQJh9EaXU9GXi5u4vi
b7tmZJ4sBXo2gRt+kgdpP/BfX3szVP7A4uw3QCySDDe+HFAC0geJvVio0jHCenPN
Hec4EtwPa2TvvC5mBx9Pqas5bkUoaISI6Y5JQw8f8jXeqEM+VClYW4Umr0z8JpVL
wz4YoSN2ISaBDy8GdIQ7488kVBBZPDh+NWeW95mEYolaHiON6fVsy2O3/Le2fQHV
2lo27vaX+tQwZ75JeKZYAk37XJ5W8EHv9LR3yoRCgINewb+U7c1ta3G8/YdNfV/Y
7JZdog7oMMM+qaCy92S+amFo1+FWt2cCx6pvTNlUXsEXNSiG+Kg+fLENxLrd3Bmx
tFbUEZQ9XO4RYbz/pkxxort8xYWvpScW964MPts/Qg45YFh76bWaLoGPbhdNpaJv
ZU89IDH8VDNAAAG5ppLdMP5ueXxRfvRxVXpoeS9HDACg3xvlm4FP+JA+6/b2WH1s
mjEG1uWYxxQuEafAIb4pLqLxMs4xOwqRU5FPJ7Cw3Argzj4WEhAx5AcRE7ZlcsZo
pt2k2/ob3tS5q6gxqgA8fwwWmJpiYHNdzNqPflenPbkbEykT6hr7MGCpPv70JLZW
IyEXEfZCN68gf06RGj4H3hXU11AusVJVy68wXG1FB1CjWNld7bIyCCz65OxjkJPk
Utfe7ykY0IMIMvjN3KOhRSbJ2uoIDFOGUCxTNHl8tlJnslbob18yESotb7U5jW7s
L1z9qTw2hbwUgBcYdsNzBO4KA36H715X9hIe14aBTYmxXvvh405vW4wqzgiNN5H2
487S9CMt/0Z+GX+/HN6WdatO+wDhqDluxMdIoqEPVvdbPkKl9cKtHmNgHT0tHEyf
WuXL4voGoEYzsB0KRg+bNh/DmE23fgdwsKzRnZI+FwGfSJwx/LngMFf/pbGIClzh
LLeZeSrcj3lsgp42Lap8E+Xy/k9CYIwtgEvrMAMWTs/01ziyMnx36trMlh4gqybQ
PKXIzQ/lxZCDAXMwS202tnfIihj9igNzLXLnpllC3FMj4wj+dP85/0LPyuZG4o2x
j01sqoOf7FTuGpU/9aNjEoh3aaku7YD7ff19NgvpJfmHynjP6qHDFp74sijMYPCS
TKp3RyKJ/K9SjB/51IfWfE6eMKzhPYztWbBm1Y4LxiJuPKGZUUVGCRB7B1/N4eR0
qnvjzpJ1oUy73ye/NbohUm1+LXG3IHIci+QKUYFAXuluNdBxYIBYn+/OtEJ4KlAK
kblksp6dmqeaXci670GvknStFvMPS/sbQ9aD6hMC/ToHmVHEVvWY9tgPV2LmagGY
9RJvbCOnK4XPbhKgTzwMnAXr6nLCRZw+4IHc/KKgg8b03pK4ZHNGe7H3Xh+QEz4g
/42SKhr5u6/kSN2dHJbjyRT/XuV9uoJVyM6m0sbaAcDaFNysU3BwZ9AoR+a0zpaH
Zep98VfCEqsQEdIhS11WEyOeGTVyNxFYxH9Zyp+AxZcBC4R6bRfmZKOo1FJ3iz3S
paQEzRNzc//LF2tyu4MeW14VWV5z2MGTaPcK03Jb95jun8NqzQnQjbhq2wlM4jUA
YgTGmdiWNsf/efpRmtGH9lpI/jdN0NYwMW1HvD/NoBNtLRSqu/ybxD6YoZFhyfcZ
U7ZAk//6ZhqcNPbZRbxCWa7Ys5QSKAJq0e0Ri+zxWNKvsRMpCwxNBHCE8+EyLPl2
rvjW08A0feL1j2nLV4UHhtL9xDemaFJuzlUK8Yed3ziiIXgfjM9Qj5cb4Ehk8xTc
7vGF9NnWzLulnq7dnsrpEZK1K7SFSa7jU5RTZoR7Q2/ew+2JzVcReZ0Us7A1hXFe
RifTWffsG9NxbqoiLpbvI3ZczrRHYLsCOyapYIYaW1RtUTzQJ96tKE1yEOEBUjUR
n6QMTesyhi1Fdcl6Pehj+lxpnMVQqQHDVQfs9hLMbtX55DTZ8iRCP+zwntrKb8V3
3GqsY5o6q/pI90lXNM5twhHrp4HbdSHcSxO8tgZwOzbXQ+XtbbMXgM01FZDweGbJ
Dv/aIDD4WXkT7cHbXxWzFctxxCKczaEUyv5rqdCbG7GbyJNq7jzXeznB2akAEuZS
qo+rnQ3kfj9bE3Nk52sc6sF7uj87VjBqnkKWfxVyjYckH9poFgIBWoNPe5IkkyON
A2q8HuRQabBjMidORaeWcRqZIxoe27YRmY1g6V7h2VCn2f94IbM7S+WNMR6V9Iyh
zYi+dpxIIwbc9eY6UwB0vlpbf2/OEami12870PHGNPYytu1WX+EApZ5qMUQnHlCU
n7J9inAiNbMT0Fx8V8lljv4LaL4hGF37nQoko5TuZUAqCAs2mSBWRC3vnj8yYFxP
LRrZIOubNM1pj1OqQIHss8wSULiFEEWeGRPxTh7BCrTBDdD0NllamvIVvkWCGJJp
dqwhqC0ciKmHsaiBAVseDEFgjYeDVNcuUiGjMcsN+gZxqb0VJHfok6Yk7ZnkR6Oi
EXec237ZLPbd787nFCMIyKU+p7q0Z4vh+3fmUu2Kie3LkYTW8zlvD6yTJZ6VeRQl
7aucv4ZzWkHG0c048ln1iEDsAMwz+nnXTP0nWLhV4TMfJTlC06QqEhtpqXOtih46
5LekJpJnq4rX8CmwFt0EMXM2I9Z3UU4MuFsqlWz2DubB6OrnR9+fS/REWf2BjLOc
tZTAORhMDycJNy3DdVMaE+V0oFrfaevP6BSQc3l4yYaQigZLt2t/ONrY95oKiGJb
iaWhfo6Dr++vVHj85naDFJGsfF2XJbx2gCqmcFkJJ4Ekkv88LLh+FELCHbKV4byd
fBm+ihYiIP25kreH6GUpTjRW1Qso2IyjoVnzALJmERhJxV9RMI3ai5S+4EgOer4D
qts+eh/M+YNX2+Nq8f+l60rTQph2YmQILh1y6Fn9AOHVxYnrX8EtCnvEMF9ZfEBS
uPsyAaaGCNTts6xHfYmGFp7adBuertZDvysMOieFfFMObueaKT+8RqGaETtquCLz
DOSqHthLA+SuCu8OreV2Zn0m6d9oxPG5KGdBNLv9RDx10mn/7N2g8lsVeJGpJxJO
yvxt5A8B6Jt49iURw/c5+zME/W+ZS2K4bofj5ZKbohSDAPVj48ZcMNY9YIS+b+rD
e2kIHTBRFH0fuDF2BXmLVtXeKn29Hha1Dwzq2k9rKx+xroJ40dePGvd67XmOl49g
C5oZ8Ue7F/42DDIrEUkROvEOXhSvTTpTz5FtTdNxP2zJcEqrPPkPSY66cPb+uQan
nnYavxe1IXT5XkgCKJiyVOH9BEYlpbO25Y8A+5AhH9mMKU8LtW8i9ZG+L/KOLDPr
SuZYAHabyusWMMOvark0InkSgI1BSEzG44k5+N614XFov+2AfVTC5PZHJo5PRtP8
KUkO/YoZLrvNK4JIlIblfsmqxJNRGXZmsAeZYBXH9aJy13HfvyAM6n35K6hO50hF
5hDovGG0RlnYW0hai7a+XmpOlscppEdqfhxfRF5VADFqQxTT9MhwCgDJdsFW+Y7D
2zAH4f1UqY8i1jNy8ASD23pwHScSumLwYEDkdkiBdczOi5FQGoydU3dfXwzARxOr
jTG/1k0WgsSds3zdcyvoLw2lCYrzK7/0mJOdmA1JSm1hEHD69RkEi+xX+4fYp/fL
37RdJYnSOxgrf34LwrUb56TzJAr+3+S4xOifNubTLK2qXhTg9pIg/EySbBPWWuyZ
nlS9Ki9dNxh60DvL7S7/mW03LA3kpl9VcfSSWoDx+bjYHlnIald0f573Z46w0ERW
HeTNR17nScDSxsgEA6HMFY9nrFgs6igyTEHh7ZQRit6RSrLYtpipgAeGDVQ2s/ah
HNqGunWIkBZTrWK8PgFi1mjzhWzGXo0BS3fmgSUbX2YmzTCjW1A9Ppxyu3JAyGD6
5IwfF5C0F63SESylh16iqfauZIjH2o9LPHChABZNs4YrvYsO/n9drzU1W7eRyxeX
/gc+PhwKGI8mpJ5PBYLp1Sl7yFVqvbc18EewCtse3bQggkGuNpRVDlBnmWMnSPx3
Lr5j3lNJw7/sAXDGGNGmd2qcC/p01jVOnWtUXlkT8KiKu9HOlyThUO8aKZ8Ddd2j
S9wHkxU6UD1P34qVo+p4mgtQZYoaIlf0nwG+JjDRu0o49aEZL29s9zIsDBQH7b3J
DVxykzwv5UfabcXSg5ozBgm+OniIFbebmxNY7RDPxznn4x15ritgu35aCN91xkEt
mftVi/Cf4JXL0OtrmjbSKxvG8fKFYYE/ZJouxZ/MnsamsmEdDNoGG59dXO3MKHK4
guhr7eXGi6/8l5kArXgaisHAZRrcNotqMxWfv8hhqcUhXlBldeW2XTWRaqGzMtZg
cTpnj/DvVcnhC96Z83IFB7ZqYxy9NiGj6X4ztsCkRpCKp2NSEx5QDL6ratqj7WBU
68uffixYvuOPcPdMmc0ntYFZBBe1W7B9oxvh4X36edhpQ49lp3yNdKtDKcalR4lH
kMgtvPGbGnfuiip47sKKJMCPgE61KTM+tiryGHUAyERtjUUle6p/YIfEn6udMEaP
l8nnqlD9W0+TN90sil5byLa3hCiD3YA8qB3IveJ91+3VL4fASQbv/0yWaspUwU8s
938Sy8g0/05dtKW7BSbFP2676/3sV2cAnzxkDt1lzlYWoXv6ZriHIcYLmK9syswL
ufZx9PreABFBJIWkzFBmx+K7chLRu9RvLxOhXFw3YCE2/5nKEWZLq2nmV+r7bGgv
3KgJ2sPXoxjfn96A1Kt3yw6/3FSAnKCyVN5Rz6gcwfss+oJjFbgLxEgWNQ2swXIf
GhSpRjKtC+wSv4W2PFc16hNYYB308sGoKgvOm3jmDuICpXHlm93CfDf2V6ggjRE9
jjsXKrIVpVARWf15GmpJONb8/h5bz1G7M9L/avcN89i+oReMNqsFDwPpIuPhoppq
upcZyp1JJEkJmlPRSCNG71+biWVIv0CqNaf/sD5KTewOFAUiBa4AlRMDljfnimXa
xYDA/fgdHvK5RJysS48SmM1CV1Ubj0/VYng44jL6ne00Tbq7LSqCJMWABcU3/cEm
cx/WYsH+4uOp0CQ45Ye3DdtKjSKESpjAHjEnECQAGZAR/eLpf6vpx7drjEkemfAS
90qMYinU+K1KztNag9/mjmByflo6h+ctFb8XgzyjondsNoNf9Ndj5OodY98QRHyz
DKdYSk2W8lv3VJdc7R5KNpZ8rWvQcACQ1jp6gruJF7U7z5kn1o1m0GboTY1ZkQno
kzRae4ehyJxU15BAdo4UnRph2OFrkQVU+1t0JcnVKFV8liV3DirFpuQ4i5VvwwMv
gFCAgViuZo9vW6eLp5nqdNV1cY+Bn3ze8fGfS2mUc/tYzEotoCP0ll1+pHCIaxAt
icJPQXbxvFtb5a7hTzh+EI4csNvdp2EaZJjAXCyvXIGZZ5OhQ9/gwEj/OosDyTqi
n3HW4LCNbDMdJCKyGl9h4SRQbqJwYcJGJ7o3Gqx83mPL0K/BKCXVuCFhLO8afjav
/HHkQ8Gr/GllwGe8yUkXFCR4dbDJXbKaAl5Rdu07licaX5JI9kZ792pP2QHHpF73
xi2q6BPDiwzVPrRmNTsOG1BNfTyrJlLRA13kmViT5Ysb94272Ob9UlDYG79B1rsU
yc4rGkd9rtKOe71kwEn8p4RgVYDHBGijdk4qMkK7Q8VeS0liDFc/24eDVqSZjWhE
+EzI5JBH+WcduQCQtc/pylkemCJvLcaoNa0U2SyBh6ECPfd92DMP6l9PRdGTtUtv
BKRzPEjCNc2FEaaHBzS7J9EUEFq7OObZvZLJDlJSf1hs4uR7h3thhY4VwOY/mkXo
EcQ1gfHcxNgu978BOT+IKkqhTvdDc44EM4h1odMTrOaxXRDHaLpJpTXqJ68lOc9A
jRvczuCh1S7X/KMePH0xAtVWc1tc5rMQ3uLEAQgI0TlsW09pWw3S6EIvjAIlJ07L
E0qiOlxjBcysI8HDBGgURYHiK0Ec3uHPq/3ppM6bDuPvfDB6LJ6S/nYrCoHMGLpZ
bXqUQwLGDIpQI59vjQQgS8i4hLQq4bpjmnGMlF5vdU9Pk5Lfze1FjDa8LkWU3LRJ
oWoZ7msF3E7XsFB9EuW6pt2CdGmeuQL/xcA8JLWEai9yWLSBX+2WTaORIQQpP2Yp
LZDHE5ovoU78PEEBXmhIeTfQndqCi42eB+j/nlnfepvPdKgO9bdn7ihJRF91EX8C
2WtERWIRchKrMa3gauAMPE2ya3Yr1o1PEtuKEKMfAAwqFWUILm/QAfBG/UnqMtVv
4I/aURPRmkEiLhzwozgUYOP5NUVBaWjeVOcOnr/jewuIwS5CqNYK1Wcw7f0cfa1F
euf1Z78yWx90X+eN1eLBEIsUWDeyjb+1qDEnI+zeXaR36F63uG2BOt2ddPlb6P+6
tVg7UQpHMZAOzLowLqfWRuooPmNNx119FGFIzqw9yBfcIO0kNueYxnpB8fuxhnnc
5c1xWONv+H1D1Apn1PbZsLmbUWOq3lvqWJfAQT3GU/V9pn7mcx4VLb6Nd5wGEqME
r8HbVADsPlTusNY4BnyscQFuy/5zEAfhk9Q6JXN0j5ioPrPrxVVAqScmA/tgUD9/
zS3u106tCBHIv7piZzMC9HCwTGuvzmy+ypuILB4qiao3+2KdJyeYZu82d8wBCzCb
9UWSrdPtrZ3DhmrhxIXR+YvTtwWyBNSp1ccwqwwcBO7KZEzE9UfrKVZREXZR0mhn
GgvlfcwRMIZS8WcapFafnY1segGcBUjPKRadKkN56Wbw1LlQy/TUlTf+mo36evQp
tmNIfvJiboAOLpMpl4YhWR/hOm7RSdA2dg2qNN9O/RUH1McOIoADiQ8P++kXM1me
IvGqucQRoHO2WwThOEtSamkM14VuDsGXfbTrkn6KCeBRy03RmnlnJ9dXDT6fnZRT
DhJvRg382Kl2rWKmBtoOPnH/32KxJpU2VG/WHITN2+g86OXKYfAsZLHhj7EUXU1u
r87muhVsI6cS7M/Em+WJBShGUwAikgCIRTphehUI0/2iej3qEK3XrAoyDE8h3+8v
5zH9+WjfSwtFxTzUypFSii0sRodpC+scqRIEbfkuYtqB0QXg/Zb+Vctr4otMnIvU
13auGD28NjSAvc4VwoB19sPUxo310NeVxxC3NeEhBVBurwySMbXlwLd8iQmfDdZU
fDCks7MqvFG+HjYiZG9Pw9xCkuMViLufJWG8t1KC1EsuNSYUct5jMEAKuKBSHx6M
FeNdLf0dvKDIIshtAFzpD2MPXYglcpG54fIY4fPXXgE4xpfnjyC+hnRGTkQhz0cJ
iES63Mq9DVj6V86yj9xIAbTO9+jt93US5AJZfWOlWlsLQd8bSvGQ5Cn4CTA6yExj
CqB9cwzB2HkS/JJKn/uoynY+jD9Rg+vjlFb4HZF2aoTiyFozES1uLEyGyVbKcorn
Rah63IE0p5BJjCCBqJCUAFHAk/Q9EFPP4y3upB/YfEiwDUKoIJgbOw0S7bB9VetM
a+bmqWWZKgBTI3du05fWQD1Zt2jgvhmeFCk4APz8wxTBB/8GIcTu3Eg+EZ4Wk/St
j//PFV/EjK4/oj4Z+GqWX1CetPqxw6q53qdA8fVSX2zEo62zTsfz8jP47JrxGs9e
8wJS3j7AfcVuxxu+rKd9v1ihzm+x3TLlEG8kHRUSODF/kO7eqmoYU6C6BPv9t87M
pRX6KlucFKmg2ZX8+qheR6ZFHEzpOpYOIY2Kf+Skr2zgtfZ6DOuCAKt2xcR7M1d9
xE5U0DsA9n8+hTBzvB4F6tyt34xu0EWkuItYdZ1Ocol9xlsGrciFdTMge4az6X2x
y5nLv7ZCWntoaNtF5lJ/LC2/UQih0gcmHw9838PTMpMdzREwQICLYKpham8TKgZX
PE4+IQTn4/5ic4At+UaFg8Hwchz1HGV2nfO0dzMYrMr43xxyFcDUwUgRZOBMg2mb
+Ex3tpDWMTIZLTnrbr0EKnclkbwN2Y3tiiQL5ljjolxkMaAodC/etWWf8DcmnTjP
Q46U9R4YXtLMbrXC3sqYfGVLN+P3qxzXQy+Pd9V+Lb6TaS+YEsUY6kR7BfQ3cqSs
U6AuPB9cF6DVZG+LhFYRK7uHnf3f8AwzXLv378SzzUzcvGOJiyK9Z89eoArYzNJo
KF7VaE2BL8EeB7SeeeHSger+GQk4jNoiIEtgztNM0yRbWvJGBSz2pOpmAcGIeCsI
Ua89f9rjjF/Q5TAth/58T4VIVFl2+vYYRUrmbdx1BMmVHnz7IvaSwYXWfKQ49BWm
I6PMdqZ0IbFGtbDURNbdWcXKyYr7yvqwCmvQRKz8QvC2e3P/FHNpSnUxDOBghbUD
RflqIqwXqIU8FPs9YfSxzoKXHAPyfFzhd9VryhJxcWXPsbqUXVxafsd/sc8ERGo7
si6iEx02/BdLlT65nZyXnCah1FWdHx+Wksoq48WmVof/hF5lWGZnwnI0p/P4PqvV
cYWt8mxo0a4jjSD0A58uI4/l9/id8xhRyG1pdyE04gxHUA3vL3TSopV7+XnQChWs
ucKb5ig24tc8Qe/3m8JJM49C6zDH2jHMhtFAFAi+qE7dCthw6xA9O4uOyFQFzNUr
mj/+nhPvSRdPHco3UwqGbBc3TuKSr8Uzw3eFxVCvjzHl9VXv0cIkb4x2IiJ13SfF
YNaryXszSwG98c1QB/V+UQaGi7CW7BoY8x6jXdLy7YINI/zwKEYyq+2x4pxkalFl
gH/n3aD6JcYAdEIZIw2d2d9zQS55+e3VsYa0aG5BvZY0VbMqlXomwJRJTU/Xnyyi
zD+JCzM6wlFcQbDp6Y8fK8NnPGDbN/AoAboAnyB8Km2IQtuqfN/ECxtpZSZ9SY5q
rcwqVOILp8s2wQv6wfwj4B/1oD98BE5moPuXxZvYbTYwNTFQpiPvQMIPIyUw6klc
xLD9wUMsbwAY8ki48neYg+MEQQaVa0gfAP2wO17zZ38OV55PJqTRzlQ1JKc+IXsy
q/gQ46Lc7OA1uW8JGuIAIp/BehZAelyY4RmVeUdpkDRSE9Q1GCv/Nl0mncXWGXoy
PY2s1sPuvYAAcUUV/TxM/haanumQjNIsXWrsTJmpmItM02xs/yypFrK6dzO2hbxl
5jdc0J1kEKi2nRXpqzC3GyHO6TADppDgAF/kRdf9lgh3vlyYDv5RMKG6rJ2uFmS4
pViyd8ffINoi9Cy07gPUJ+SFkF4/il/rgrGulz2sFK4Qf4ZzGFdhLX8wVMfqqjt6
vMe+2jIZLauTXkBq5BxwAUHO6CUGThN0o+BsnED6Hbs5d5I17lZcrKp4CDiSrnr+
DMK9s1FyaBd1i5IGW1E+Xr+9j8uAGswy9YWaOfrZs289hpeBpl/2VpHpvyw2BeHl
Z43Ua79TKYpFr+zPDSv3PM/6/D7EBEMCqdO0QoogN7JDdbQ1xuLrIZzWlET/GIZ+
TBcar30KEbRu/IhUiVXhfFHSoP3f2Sx4ptH3w/y1l4K1ndLvf5hc1C5u9jx8O6WQ
64LTDTz+7tERwYwpsbeOdu3qpDXMcF/kRbXNkcD8VpjYPGa/MdFugLcRKY71ysh7
NSerbMzPXPKNDxpn/q6drdOeuYrfY5Xp7pFAdUFOXC7cde1W9rFnb63Jj0x5xksY
pPRWGQctU+jRC3MBU99fkhtBdz6d6/ysy8rvG4Y+621CWbWNKyY4hWx/zlEB+j8R
oPPnOp0VL+RynmixL7i7tXgd1YbA8UDk/sG1lNHQSPE11Cl5WDFNeXVWbd5E/Y/1
qLehT1Qetl3DAyB6482aRWZUBSaehhWhCv54vV2QlYYA+1gImv6QHcupq8rpxl5W
/1OPyDC1h48XawYSh1eQKQ7dFg9xVNS5U78DUNB9B8k7RdEgxBFywUBDD32s15TJ
6d6F86Ifz4M3FXcFEplEJWh3KSml6YVkitN6fzZKMdZsx3HVDYxdLGlitEnjiJxf
aPgxFJ3NnLAkBmHA3YBGD5eWySNPsCWVAMLXYlzNfdjzhju6HJq1EiUkVf24/Us3
VVUf2he6rjFVzWoxpZ2UkaPMqsiTDqv9bPRxJ5ihxA5VAICSBZMsIuzGnzWqwzwR
lCP9jB1NeMPnOJZK4uqwuTOEd+Gc2rpXveh51S1j6giupsJOMJlh3lkAvJFar1qi
tyd0fg7l2fj3HPY5MYDYku6uDd6JPXuGTe7YDeCT23AX4HeqDCeFJ/sJjTNMYWJ/
U8BQXTCccv/mnGAzKlfCOeKxYh5cZfZL0780esnvEDGrii9Nb45GupduZgLcds+F
p1ixPEaqzZWA2ukJ5v4PPs7MFE74uOe/obGuU4rb2+0xcr1Wj7qVhTeGkvrwL1u4
aBvEG/H3UYGKbdQlmIwlMBXaXVr0S8uhq+zVebu8Gs09PdP41xmzDb87L9Xjh8eP
VCDfMS3nocCNe9fgwsL6y0JjPIwmCkk/JbCHhBFJyxyEZdZ9qjDxgaT03qXRSiTM
dDpN2mZkWBKsWFgbDwFHe2UjkOKR90u/BFxjQXQ6h1XIpNVVSXUXVDO1QCzNbiNd
i7nhI4/V87KVfuC9534+0VkjiwymPQCsF5snuBw3iPQzz29BVPQdOftjgpU6Ro/s
vYqmmzMgiJ2B+SdsS4bETmCitc6CvTjnR84jHx/rRVuhYe/yVnKq3S+6fB6ufJ6b
9uX/ok4S/YudXoFHmkBwc0WIjQcwwbt2d/T+RSSwI9cOtg0EhW8n3vhpGXZEQZRa
9nUFr1yyFFjZF1/tJS22w2RATTvKK23/TjRu9v0WMA9Z3BFfdkvt7sidD19zSLNF
2L2B5lM6+cby6NRHLC+XwlnnIRKVKGgpsQYDy0p0AGgBy0YkhfVCpWMEOcj4P+cI
ZUovFR8zRnirx3WDqHKO8viJbSjcHAT8cg8McdhOaZen8U4mHVFB8EIdue99CMNF
+MeA2dnxgoDhzmxiN/hjcOwXXcKe76Zf0CZfGjMPxSJ7wyQaxWjuMwSnVaweQUw7
+NeViozwwSP8WyvkzfK5QIKSTh8FuIYmVzplhBzwR96stIZOle/w4T7qqMV1FcfP
AidxW23sPMCRQR2fd0/Q6YLkgnOrrdHN3UODD1f4YXgRG+94nrFUVDv2Afjuh39g
lHCF6dbJcVjAmwDeyaf64ouvGFN+g7hKQLjHU+o/21AHSCH+WgXLXfFRjxxLHzf5
zArUMJJmrCW2wcwrJTrG9F6NrArwG6J3WcEyM7pEnujvTxrIIfhaiDcyItbVCBHj
PvFpbB2xhycHGMnTg1umrsdTm4iBNYGiFO+L/7P5s+Xy8pYZ5L2691VEC7j0+Jxa
pC4fdlzlILrgLyVdXVeiDphzHPvSmtBV95x9obtzPuSwAu0JE4p9eYOPcXLsn6b4
lzI96uPKLCTrkPVj7xA6K9RvN62H9PSaUfiqWDr46L+kyFTRncBPTOTUylOHker3
Cz6/j635mSicMX3m4bFcnJ0Yf/pS24zVp8YAaNOze6LaIGAssn0QXpdWvRhJjlBu
gUPWb3wF0RbTFCIJ9V0AEpku21oSXLdx1VQA10r8eju9STwOJtJvVv0SoF/e9inR
QWCKxuCSdLR/EXUXaLtY5xVo2UHDTkcWTSqptBy1hv2YXmDZS91IC8LzRPdHqHMc
Ro+17B7uc09OWSZlYLi47dQXNVWwBMkNDHmStNS7s2i62E30bhrCf2bI9Z5f1bm9
JZ1rj+ISlINu2t9CtVrs4Ec1EPcAoFU2ilezGirFMkVE1atRODcJ/kfuHJdtM0Wa
MEohToC5/NmyOX+HwENvGYwdciX1fQmBYd2o4uasgG+LAJbOmkV6Ta1y3W/einy3
Rd33xa34E8aTSjqkg0lXnlNmEPKebdNuLW/Se81JOg6W8/W+z6mu4l8cWFqHfrNu
Ne2OjYTWohaBS+HLgoNHqqOQM4LH3L2CZdQ7FHzvk46qMf91d9k4oeQJgu+TGHpN
SI9x4i979MjFQFcUNJZu1+mVPe5ODJ1IXHsMwI/KGZ9C/Agg+LYEdgYo+LgxckJL
PGEVK9lCm5nrQ93i65nt6Zb5TGm2VEwfSzq7giBVCG9268jwsz8Bq9bkKggNUCso
Y+RkEeegktSbKyaKeW76svQ3GaXpgcWxqK3mhkKlVnv8VJZvPumcgWdGUVC9yHWs
M5LehbIz9e5d9QV36JojEJzX4kTJe8lC+dGBBIUZ5yGk3dqYjwGLBWlBJ2Yk+iaz
h/SJmhtII9YhB3os9d/JTk/3WwSAGSAN2pscJXXQAUi8rLtgwyxDSdqHeg8muslM
BurHhfKGDOGrHv0Tm0apcwHYUKbKz3D7wE5+zvnretqIlXaGE8zryuN6anF69Pkq
sVn7uVu5w8mVU2Cm/c7GOX6a8TvfIG4+U5iQHfAUBOYjc3GEGskkQhDY5YEjJ6tt
ibwWOhsEkMn8+7sMTfMYPsaGsCeMuTPPsK+ohOyXpAGio03qn0sPAAg2PnNUA3gT
KHmODOi3Xg9CQdHcX+NnDJHiFqCkbY+9Vd2eTGj5fo9JDTZwY1U6ffLp29QgrvSp
dPmqhJN+I9ESgZjboYrNeL2LYeKDrTQS4oGiq27ICRFQYH93+Cu6gsxgIgrHkOqS
O6AGRHzQK7z/urXX4nGH6X6ViMPCVvyXGtsAlsgahCiuKlBk/t61LYtXBNdS0yIc
4mS1KdpdxuP6QvVDEQKMv46uWNa/d/tK8/X6GivydQOV4HvY21OGu0r5W/xSwww3
tmsVBAp6+SMgRTEk0DKHQto9Er/Z9QLBDXIBjZjLkO4vEXBHlXNOB6HeZF/rqcdK
puMPmIGuuXmpTsTNxpc7zzozxwFv/jP1B/il6WyVHSSTo1ZChbfhS2EId9ZTsHez
wueC7J7WaCloFM+WxNoDpzOlJZ/xu/0IYvCdgdEeJ2bODhk6z/PCnwgsWR2C9ozu
oiDb0V1CUWaxLe6CJdOKUXSUPpJ+FDqxuJEt6JjbFvrjbNj+o0uYLa6sDr6Mfrs2
xT0088B4KUcVVU/NjNkZMmdwpY6ZbzOdR108Bh1D6us1hpqSbZ57AqyndlR8IX74
QWKUrUcUD1WI1etTqu3ZHU9UhIGgESKzZLqnQeRRH4fgW5VDdS4FZnglYRjr4sR0
2FLGqAdFzw0TEcHQaO31Wk0yiky+7Jj00QD90dO2PKgTHKiXJTaSxcDbH9OHS7P1
F+1+CjXf7eNRCyzXruIIsOz9EEgXArPTdO+56QUvVFOK2P6npT5Bw1M3UHoUfHGD
PPasIylsqQKdvM87hGEOerKnhL0atHYZnQsuxuQy63gRqJM4R544yclgzwm34OTo
jnTDO3//CKeiaCy7540/Vs7pittoFuLqE6+GUWaTljcKiD4U/SPvcifEtxVthNig
JPWmQOcoiMEDgBW3jvd7YZMrL3Ckn2j8vQsYDUM1RU//QopoWJ9NV7zJw3Ju8iFF
JYZLXoUumq67Dn4Lh6DAxiwvmT9516Ds9CY2v7u24ufqROIs+ba+w+dqTAWMerNd
U1bGy/gKM6fOTDdmDr7qzPUKX4LdITRx7GwLCz0gG1lY9xJ0bkDVZoPA8HguZu9G
qEH2yVoSsvwGAJ7vJjbx1RLwx9XiHzLO+N14Tjd+CcpSZ3XYlSaYXpl1Ei1+6lXr
f7gdD9Jd2idJj211Z8DmvLQe82w+QeCifXT9nhoamBUhe4a0yWzS7iJZnPhfDxUJ
BK1ctHqWuMe3fnOC0KhzK/xK3op7dCnO2Xt83X7xsCYKwv9UprpdXCWxxG1VzYJP
xrqAVoL568+UiFPE9slmd65LJ86P9jhJAmHkNs6qjuPjpv/8JAGHEDQipD8IykVe
Xt4VVC9ZZd0UDIilxhXkutKCKgE/S5LQMnfBU1Z2VAkdALzAdxhf+dYxy6yahgaZ
k48GHcj0Vsal43YajycHJif/BmFrUYIIzj4TOEsvNXzJpxapwGL1JRGMoyL+19ii
0b7qQFfep2Wuho8LW9JzUAjO5oS4pQ2k61bD1+Hf/D/kj3+uvT85BQfcmkSGIu9g
zZY9T2lH1tlj6Pq2nnvX7fRC0PVOvpeSN/WnrOrf3qZz5WNTaDM+qlXzpZCPahyo
cvunwp/MMJdta6TiMu1Bp1rgxcDXqdnMD5JRcPYk6x5FTQ8nUOlmBeOgosaOah91
jnTMLRtmdLe25Sh/TE5nN9cBEXL6exlGIoEvC4GSSOPRuGC98hTI8HDgLoKQE0Uy
01S+8NrwmUMKV1LpU/DVwr53Ix4600xVs/DyprkIoZPWjoy7Q1K0AxuUi+aIw73Q
51riMXi0NLEYf4WnDRhvW8LVmmO4vfTL0apYpaYLTzKEQgcUJCr8gPvUO3gaIW6E
8C6vpb0ejKxzatC0Y1xwtR9qaCD1FKzxoROEVW+v/haPG8PKxAlzovU6DFQ3tERl
ygp8Esy6kh92zyug9DyP6AiPwM3MEJM+rm9VASS7n1y3fclekhv82F4sqmxbKDcV
brmsWR7Xgs9MIwA5dXUIKuCKOFrvCUoRVOpbLv2Ne5DmVJhcrP3x0fzqqzUjiIP6
m9H1P8dSIXXglbdaYxMG1YHSosB02BFY4Ipd9jMpF4Wj0exUBJK8Ckg7ysv+qu82
wwJyII+2hyRN1upzkj0IRa81Gczv7PImxwmbHllYDGuzsRW+mqHn8DsEdYcqaud0
11AwwvgD+j7qdjKk+YRRP1MPrmdWlaZX8ZM5EptTQkRcGPL2yJ3BIRPQbXplkJjZ
S+5OzHQnvtdUPIpBFYbk4nnsi8OUkotjokrw8Kl0y0TlPZqNjuBXaWa2p298r1RG
PCEq6WfcPFso9DGIiF6xeONVRKlBqY/IMyOu8OXworEioHTavSnBbi52Up4eM2MC
3oJH48uPdaUc8yMa0ZWsnp94JgWYdsBvxXWWUJxFW1tlHXNy1RqwasTmpOEQFGnN
Wfn9at7VFTwc/1DgyF8JQ/LA+d78SxVLH0HNkEaIHmVmEAPqpS0LD+jggN0V7cco
sJaB55r9uhtUDBSoesZh/udWCDvsca/FCG+PzwSngj6KNmVOnp9m1JY+ORTq7Lj/
IXWuHp5P4JP1pPbjq335GPMg9Zb796xzmwZNS3COxP2gyKkP2IwyntJJbGExLXbM
MMuCwOda+LvtIUUDMdeJCvj85t8M+FsZQ4MqQdW4New6Kks1JX3ZZvo375MR5585
days193UfPib2zclVWAMOKai8Ir5YmW9djG35+sPSh7Z57UzBLhAeoJ4xg0LDcMZ
oKiDv+tM2oSchdd2KQVd1P5Pqp0mZFLsXyPRF4J0Ot5/tvxyIIYaHS6RyM8lmgxf
lAfrDSzFJZko3BrGlV6dr04AEvm+zmkVj4Xp7GrkBIVjK2kDUKEI2htelKArD3cj
ph98+3HLghip/Fd6skWcrSgl9mff4ZFizFkECxfLXh9ua3aEq4aeSrWZHKb2C5Jl
8zLIIRpzvS6lIl2zkPe2bnWeeSyvANP5vOcxxBwdkjF0NqIk8N3dk/8MJniRTSzl
DmgUZlJN9k6wjC5mUI6VIhwKKruiHdRqSOHUZFfDnmuEkE/hxsNp5CStO9/miY6j
zb1DulJZ3u0Q69n6vODObwobao8N8UX+PDUwBEx3AGAnrMbMdiYvikWqFD9MZfBh
jVhM33S/5PRZ4YC8JjJoyHGaKoHcHNBFMxEWfcRmZ9fTK5wMFebxnSsxVmJT+8+r
TSrAmSJH68Q36JO2htxr6vt5sDjTYQEPu8pbEnh71sPwElErkUJlG+/gSWygCFg7
p8Yi3mrcZbeHNSYujRwVWwpv9+7D5t/5RGEHQqW4m2oxC2RyxE3DZ/TqB2en3ITr
3x+Rk4fw0xUroCUz4pdQMQXLFTyksodn1Jo0a5AqAAZictO8e7vfg0TfBPAFjodD
5W0XtZmrLdyarzm9XKYz5kSK+2zEM/SApZtMCkAypkms4r31Ta1erC+JmONXFlqe
h0RTAIhRegXxHMSmCDR24e9+PYD4s3omrjZncBDQ9EwvHit69hhiSgcwGlutwPom
FkgI6VtX8KndsQ5KoG0cbSI/sMHfqQh8TDWXHClgZ8aDe2+gXe2DMK0eqjMDgP1i
/sUT6qGOQKyurROg6ijjB6rkt2r6ZE1/YewgXxZWocuIfX4MpMoS/RI4SIXM9B9U
MTO/rpKl98va3rf4VjsgYky+wIYd/CI8ewiyI3USUrZyCLccRFhLpgTDadV3PMbN
Fk89CZH31d/ha6VHA6oLt930fbS97LlebUjjW4PYnX/S6xUZH7mUO3ocZ/KyGSkk
I1awTnNZQZpG7dJqVrkW7paXLNQZzvh+fEdeS8hzCCvIOimg9jGBTPZaX4AQUmcC
o5pGVrdyu2St+xfu08R4i02MpmPp4VMpSWnucSpCYronXBB+rn9jKivvT9WjN1S8
HD3cu0CgVB3MDPic0GRryM/swuFCh/AAIqJLuFRpwtw9b8I+LmQx5+xhJY0z4Fmc
xWe38SzWPGqIFg7MBS0rzvnLW+5/OhzUzwmtZMvh/Z9IM0Af0sRAt2uzE4gli3wM
rh6gbz3pGEfUKPt4WlgGd7lnYDwlqfiMcKiJVRw3tm2PDj60NOBXDcvbojmchnYR
jTxsAJj1pRAEfh1u1sN5HyOiKdhZRzBcUmyPfpjdOdalXPi5aNxIHMxo+ijFgT9S
vEkbfQNDrGe29KYn5JvP3r8gQcFGc5+w9JLZF4dLwflQiNHtvzjsDcjBkyGRguoA
hWjQRiQ4qyZ17lo+30Bbo16/9JyuyJ3TtbwYLRNDSyb+HUBAME+GKh4ARMoWYbl1
D5dSZR6PoC/p3KoPHuZHqjxWsN0UyRg6ai19ZZsfxT7Ajx/p12aAkDJBBWDCSySJ
ISz1rcz7wdwM4xDn3XxspQpy9WLqkMQmBuY2BL0z3rn0XrR3+GLBxeIydh3/MDL9
YcRHUnduJcPh+NTHDENzdbeR5dMVT2N5WqcRi7xotO5xJ71jeYnzsSfD+wADPJMu
E9bQmPJUzqTJLfwLSrTD3bIvTbZN8kbvZSF4KHKDUewxwl0abztFi3ItL/DU1Mer
sy+ei9WyhYgkmSIbvA1eHZ/5g9so/sp2IyPrbCRpemonArmDxwePeOMvWG95eYKu
hD4pzWIcA5E727od1fuf8acSXmBNfcL0mjrc8j9Er0zIewuarsiLlpGSVlSDRaqH
Mbwdaum6pWk94YbpbuNitxlJ5rgR/tJePprTdHF69RYO7BpYJoubpzo1Wb24mNmW
qBjyng6lBo+cih3RKqI0JKNurx3fnbZxQpMDk7KXm/7JU9JYOZnRzi5CkqAfi6Yq
DQFVRPJsTVnf6OSdTiODXTCtdEHnf5XmlKVRZI1IZ/+f/dnp42W0Az1f+F71LE9Y
t/0x88ZIfaQfFN0tkZN2Fjmn4z8KWEWrPuA/X9qf9Fjavp2p859rywCz3z+sY9o6
B3cEl/ydvAZN4ZEUAp8Bur7slBEIErd+20rH3mnbrNBXxT6JIL13cmtnhc//ljoy
vEeWdoPzKg9oERKMGC5QHQl1YGSMEYk14UY+H7L04BT1pHeqGT1PBKYVHPR4iEEb
D/lj3e8SgCBO4DYdShMMb5adM9Jq+iHocgBP0XY6/A+ycr3GEVDBosXTvcii7AB3
NEVaS+7g/DNLanu05qj9sCmxhwrQX0U96Vjc213ib7oRRf0fHC2m3OtQvYVbD50r
UUnpUU3jN8mBLqAok/02DuvtKKuAjUSXPIDtJsTyw0l2qOtA4WJo9SlnBS7ez5LU
DyTtjYPvwKuUwMTony7Hj/MMqTQbYtEM5lNMNEoQMv7UoLU7EvEM/pnAFA9zUpEn
pQOUAgoI5qUiQSgA6ord5wkRcjUfDM5WlOqgtyP7CXZFL6dUWSy9Jn+XEsmvrZ7k
+pZX/d2rW5gd8ucCRyXoz4QJIKHc82wOPAVMaL6UjAazv1lHpIGerwDi+g+N0Daa
EvnWnb3fzAAYmd62vULtghb0B569Eave+zwBLlTl4g9W700/PKah6D+VL00VxIDb
uhSPwVt+BDRk3P5WkZDUkxgYyi+jn+kBr2iPMStdyTBhsTF8wYn5bstZAQFK7Akh
xaLTkRq35+ZCfsphzkgQohgrZwyulMPuzVNmToQcwvnB4KUsxcTFNxgW8A7oBkbC
AQAPOVWf0p7kvg5v9hpF7WZMYnWgmC+j3/O2AoNVvnGVcwTn/eat71SoEeSuveBK
7d+IlQf0PTleK3O4LnoP185Ks6/7GS6AXM1suEufINiCdts8L8J3mijaKR1xwE9l
0qCiJl/AS5n7HRPzid6wVDBKfH8Z7aWEqQnaRksalKsgON9Wctet/e7tT5KW8XIg
MSEa9x+l+Hnlq02EbQLkJUzyasfWE2+Oj8Ue7RserJc3eJdfBG6kJaXe1EpnYZj8
L/g6IVy1D3g2JKNcyF/kN89IRucMDvtT2xZBMvHwHDy84prS0/FM/Z97TUYe9fz9
fBVepYftnvlO5EbekK0Lh1HTOQjjg6PFh63ph/GGmgR3AJI4pCWz0yp4Em5LWsSu
ABt5uh/YhjgnobLrzjeA4Dous8XS3Avv1h9WkKOtvwsSy3EFWRfL22LOsaNGUfFg
mUmWIiILxrmtMEEp0yUixwiS5TrT9FfG8ghx+uLInsQxljlhVHXAswEEQeaa+9eT
8Iolb7Invl5px7SJAzcPxcHuVyevADrkVhEJksdJnb9CFYm2Uy6eaurwb/LTgv6l
rtXWNcF7eeTQhMImQFZpumZP9t1dhVc0YX7EEtj8h3hjQg1nvn5/thQKJqGUIVGY
2+YVAbCL52/ccPdvfXU3RL64GNfnKvX4DDQY2FOdTvrwnPbQzk7GotnaDab4MRlF
E/AXAWmDukANSODIR8S1G8CyjsPrVUZ4RCK9pH9wXkBIwEjnVwFi8ieja96vl59V
wDKqIH5i+skkb3q7o/tADq1Km5glg3WCJv9VqCd08sgn+a5jbf3L3+nZC21SbzYu
h3CHZYR0CjCC2r1xCVph4WIK+Zd1dHs07zoRJ6KLC1EtPxBG7OgXmNGE18pxQCvj
PqqTGl0t0E+2ffJF+fgz52yoE5VXVVGKrcvh0Lp4YzXNJhXTHHLldtnM111+oHMT
4OPBhDazANHI339QOiVxaG5sWFnjhNa+ACr8APxQstUIPkoprqyqwg2tDLnQxIPY
geEuv0D0UxEJi9SupylZsguORvLIAWcofkIe4bg8XvIxWr+rqladBbQIBiBnL+eR
0m1DgvvMbB82VDUXLQM9xlkX7gFHMJL17/CNfKSwMOsaobIjM9mdGQ61CDO6EfOH
xOt/ox97/iwdTsT0MRF9npNLLK0tLipFLXeaRfj9JilVbSmA6yD6nqLu8yXiS+zd
94KOdGGWrDvBKFHU0LYWDMSaPaEVd7OeIv8MAw70hqcVIoW5gobtgF9IGf+chRYU
L//jUnGMJZWnGrVmDW/Mrd5wsQfa/ksTvmlD9Wxq+ZvU27UJ4qqK4Jw5tTrF7RMR
0dwN1sgEwzfhylsal9y0cTLfG9lRaxau/hYaSvE9AKXJOG8p6kBb5n5Q7EoZYlEA
G78zp+w2B8ToqbWKm/odRvEGRpDGJCfX5nsw8Mt31upEW3xpN6FA2aNTItcX8U+a
63A/yTjziWmYohONTwt1jcnheG94Ex5FUGt2RmhlCB9X2iJ80yEeOeHgY8QfAkGb
dYnPxh6H9D6AELMOd2i6FJuI/kbiginvGKD5bdZW/ZbFLh+7tw4ds0HJkeBu+Pwf
U/Jsk6px6sEPjrnWYQ/GKKQMnUrcyKbir+ZM8/Fys4Om9C9zmNb3fDcxsD4G6W+A
xiMxQZT1GXdoVQliPkokv6f0icbriO32poOS0LbLAKX0XhE1TGyQ0jZRMATB/6sM
ZBlA7mT8don+nioo9e+W5CNIK98nA3MNqBI+ON+HDT647cUJTPzDm4mT5s6Jisut
ydIcBuO1cfO8fomhr/7sL2wimGdNRmU7+s8Q2whbioB12/h6oTqIjYnvwJx49NEL
DCVz4GLpJ4DFwFKSnFxU4fFsk6An37NB//1RLZkkt6GmiZRttX+4pCD2OYimPmnn
MzIrX1OMf5yZcfoNsLeEeQRmKlCe7pRMRb4VSJ55RJF0F1bkCNGnPXZjjrgo7thp
u5KC9v7QVVZJfTF8EGXZM60NHvVOvviHHAraPBmJI+JRZ8QIt/hng+0b1BzoIepJ
BDRz27IGfRfa+zvwOMhAUs4ldVlDGfINmhWx8BMZqee44pdGbE88mykySKl69wnb
bMJHLwvbFw+ySkbzTE9duK2lJETW5wkn74y/AW1BI2GXW6ut+QsQ30b5jdjS0Q2B
sbHUZsmjqFjAoQhYwnO1y0OiUD6nTYsEwiPIy0LHRJgGqVpLidtlspdOkalmewJP
RnJcw2xyqvjdQC/5wiPNgib0scYYQbk6PX7maSTUDeb7AJYvo8oU54VSRoEB4iZ+
4uMUqnybw7ruiYO0LRg2PCEjPi6btm6nbqKsJsgZyIoiZGgb6+zkvV7ogryqSs7b
AhhpLN2vQc0eJ3+5crSk29f6aWZFbvN/HUAjmJKMGO8wvHqeN+rQ5PnKC0DqYbC7
fSSdY5PXcQiaj59VnRbuQF6ey0LwxF4CvW9iCQZp1RoKvg2ZRxKmv03OX/NS0yVz
lqnPhDzcL3/gtL4tqy+c7eZCX3nEle3j/0cUt+r8A25awYA4JxfqI3DLq+XJMZsu
23t/gNYoxh7q4OT0SNIXgfAzktQF93s38W29R2b6wz5HjMY01XSrctoKdrpOGkpX
0DN50V4RnNm4a9tNJ+UVCtStJNg+FQy919q68I2kxXnEuR6fhi6w9K9nRgUPNa7O
mAmoSRMQOCKAP/nua7gKy6d7B3Jq5tEvBsyVJov0ArWidJKaXghzkXX/l/lYlVfd
U7kOpUlxzc3271x8aCx9gebAXinJRTcoSABmxvW7IDFpCD34zyscCqkzlXutWH89
GkpsWs7JtI4iVglnnbbQJ183MKTig/Ll132YKHvSFTuxD0MdiD3lDkSGbDavIX+2
mGTDBLD8avfpqrZ+die3LHXmyYWz2deeMQI8oWN/BCN8O24erN7xRc7/TvacNR1/
PDFVi3dvVkcrXHShPx7+AOywCCprAjkaAyVgjBG8Bj7RS1I6Unb3gZ/QtAbQYVps
OZKus9Szp4PPmJ7sccc7nrBVnHqftvf5oZ+hHfHHTuOxaFD74nbgnq2mnc66h5s+
wu/xoOCg6Vh6PgvKnVEXmtJK0J3U2COltfQplfpgUEUsYNDJ2rhi26pe9oXhg++w
73EpBoGgPKxRHaJYo5wxLx1s8nneJQh7HyqRxGREPTL6enVcZ36jjS0dpN88jhj6
DhFJ/S4uhBml3dlb/Xa0GdMoyBt1h9RD12RTgoQ+WAMbX0FL63XuSS4VfasuhZRv
tnaLTR/9PsEVnbps2Ne9uhNGMnCGicxn2rHOsBVvq7ZQbxc14YmFUPRLwENSg6Wn
9SroRtN2kPdcoPHw6OHgK4RsfZFixt2Zxfrp/jCL0WaPPcyKBMotnrl26kIr0DpK
WPFfsPKthGGAk4tK40Ho90TgMVKuK2Vff8SL8m4bjTDXpLJnOO0fpc+Bac/cbc2Y
oeUwCXy9uD/muVp9DmtFLGB0ifkay4riY5qyLodyEA4NsL2oRQhW/tdKwNI25pka
ZOHRTUMZtQ+KT37EgTgy7ffWM8uye1niydiClNvzPgolnlQVRsDEI3DVqZ4igqQC
A4Kp6JMdiaDHpT5XLBP1L21dn3sbz67g9TmydCRgNwRggWhpanTjbe/qBSI8/saL
eE/GniPYj9djkbIZniqftj1InCG9ywZ7QbCwzpEwcDClZMicAYW2sENs7RB4/Ak/
ff75cuPGYhDGPCpGG1VyPJcdvoR3UI4VfFMZjOFsJ+ajNAULt4QZxUcZG4CO7ZfV
fhgXzi6CHze+AW997BVnCJZoJVwyBO2TUTL2cN62GO/Uo1nC46zFutwgSJ7Bv51Q
b0tqUxK+TfvrDRwH8VKXSsPN0JAMbZCCPEdskkM/5ZfV2/dPCmNS/IGIcM6O71UW
vi9iN+cYm8MOwwlgkBD3t4pIdoL+C3EiLprGpPET54+SvfHo+Wj7UoOLafZ5vv+M
zK9VJBe6EvFWeW2GoHorSjpO5wLq1/DXKsJ59tOSdDEz6NsSm8/nQC3+VPxihbse
Yfn6YQ0bEKq4csvZ5P3eEPihK267vMJmlPLUx0OcTCKKitBoy0CHT7HxnfRoCHRV
xjFb4ddLr/gwEAnF+Hd5h9NPy2evvoaAzzA2yNQhV0mHJVy637p531zQpxAn9DMJ
MGUIZQKd7CTFnoFr6ED00C7YupnE7hN65AlEQNZl92ghjf1ehPUsvrQDxPGeNAg6
ND99IrbUp1Kyfx/LWCREIZqlIW0iMeFPfTZytNRIEkO95TF7wYARK+lqTtCEKg1Y
jYJFcUQl2rf+Ge73RlUwbFPia5Jusd1mFt5rsUiByE/CAwC95Z1R+ZnX5QaTOXQx
rW9T48aqAO7bEjjMz0+G1Thklfi2pq7hoBtR2oEe0ZGbODG2Aqbo1QMqF+jXbFk8
ATHtTmZOgOaGwAkzhNsezayJNplzrTzBglP+GDWy8Inv3LRKKmC6mZz9EjNwdgGp
Cg/AZi63NiVv/c25pUIbXw1blw63Nu7mH5q+8LLfxvgZbLE1BsSgbZ8KOaKR/yLj
GzD7UxSXleATScY/0nyUxcHI5x6xBxgpPmiXp36XyGOujtn29j87Hc8ONGbbJrNx
b2hKCoYjcLuCixkH255lrLfKvY43sjf0H75oE02SJ9Kx9WIzuyFKLwKqqrOUTeR1
WeRXE6/+rdEuGjiJn3cG68UqklW0sOodAgDfd2Ne11ePDTgBBGysTPkyo9EkE9kX
hUhp0VtEOGbaBy+7rBz+ujL16l+ULouqd5GlnfHnFTczCrGX5EIZbQdJwB5KOZv1
VA8oYUUJVHL7q+5iyQKtuIevTr4qwkOxS98nMd5fhqzNENhbnbnBWNXRIyNwJsCP
AvpkurVVgvJgoqpgyhRXl/tR0GbcUcNJyUT+V/BFTgqBwbrqGX4VwgD6quWnxThv
cWOrcwc57bArnzI+moNWzVKfIqx0DUWl2Q0Kqm+oryH5WsNuLtCe4kqlEDsz43qX
UAKPkfRLT39FNwpBypHRJCRxATwQemZiDiYRN8TL6YQuwgV6qQ11YvG04ccSm1Db
mAs5rdgTYEaj3gBXxzk4tIZQ30VcgZ3/nYwiQOoD8fcbTH3nR0cp75tbp9mBm2n7
O8TGUCqk2Xb3W1/+b9JtdFB9DE8vnlrXgYrK1dgmdF2i5zeWIEQJnVbel+pMNmB/
lrzrGyvitYUDsfFkogcYW5BYFTGCnc4WRxG6Ac479A2ejfki/ZEdAa0zGjPrpIJo
WvKX5URdm57eTXlixeeSIhih4fHCAlcDl5Acduz5+6aavRq4ZQTEtr4990hsvItI
asfbBUj3TGDYZbtr5xMax1pqbmSrA1OEqNDU22xUnyu6sXMq0mB6yruBpseXwOmy
TQSW/poqPlXOS4h8hn+RYeBT/3N6Gn4n+xc9sbVLhhuNPoEtaB9y7PwGPnBsmdsB
wkjOKcyHRIKhZNQ2hZwaYWswMUDPfrxC5jApqXgAg++OEeV/QjX+9rfZL8k5R4Dh
VhQJu2m+ll5UcTCOzGlYmBEDSBFzP1ZiCFiEp1IT5M5n0CqA/wxQjABlruGO1XY1
H2oGQdFOPH1ozpolB9kQiT1iNhYQwTtKpf/ufijRJTZK1sFIDPq7y4yixvpXn7pV
WNgEDKHytVCL+6QzB/Ti+REbAqwOJnbUp0kjiREd0Xq966lhVbQBR3PFcUUY6eAz
d9iYZPnHdZFVDZvQLeRF0j6NL0dU17dVnd+qrzhMNhCoCSlV3M7WszYtxuOxD1Gm
s2Dj6AOCK3pLgQbCTfk0yvSJoWBBK4JfclxbgbWjkp+uBaSls6hT1V1J5Xac2XAB
4k6CsdH/j63gcOTqn/59JyQ4/hn9QQN3nS7QrU4JXfF2tLqTeG15ywYEOHaDEVcO
CnrxSospRpYqiopLt9EXY1Q004j42FHwlxEirqNOqhQgKBBdTX1dI1SzX9JmIvoh
dgz+7+6XAD3WoxvLm4aUjTJfVt73Fo4turHvJxIkl7rEMbfuzTFZ8QT+WUnkW2Yc
lswpbejlXNSNJGqaamg/xLm/mrmtay3h37SrXP2NEOzyUK4f2Vnq94B3Q7YFU0lG
rY4AUrJNWQsdKry+L6t3e567PzvZ4NohKWq71aBrn0t3QXsqcbByUshtiQjojNKY
/EAauR28AoHftrM68fzXluDWqoJmD2pI/bh4l2A7BN4BYz5TEfjYoN+vmh3mpnJo
lQdoaOej6kmHkUriymN4AKnB/hvmGIq51FR7iTbM05huu0hyu/U+1rao0UOAi5Do
A7a6vW1ecOT1XJA0YVOFIoI/SWzRND/HNemAyDrq3bWUmFBzCLG4jPA+Kj8FEQq3
m81wkZh+ivbJOJ70ktHJ/r1DBiF2drAVG6Naq8KiTw2V/pn/lSh1Q8/5yvAeXTyK
vQb64Ex8DA/yXUxKmlOPL83zobqNcDCaLNox379YWW7bVSlELvrjRaeyH8ebNaNK
UaoZuE5kN7hKTT1q9rIacWHAl1LJLyUTzi14gSdjMZ3bQZdX93bY2mVlkVbhIzTE
8zfXD/RcgPfI7UzWW6cKx85eoIJbVyOsyAcB6ev8Y4+k71CqzDvB6zNHnsxX8ziR
9HOjDrPLO6Erm3LkYVb4zNMXgN83AK1wRMa4FgAYRzyRUbuImKCT+teLNm6BIWcy
SNcQt4MA/N94NyWU7Dupv3N7k9/WcDdF+rvW3kYSFwqt5/IzwKuzyrYwz3IOrGKZ
AudyACS1/tXW7aktZJIol2AWm0cISiwpmowsCZF9FmisCzjN+SZr33K3Rf23FYmI
Pu5SjIBpiEMulHJgX3Hqrr1yppK6WPkNtZsKDj1avzNQl5RywtVorU77td9jbK1q
+EaMDtyqKvtt2XkHQ4+B5uzIngMEQU5lPg/yvyJ51oSo1xEHVEKeLTPNR0CfaRXx
KKBwKG26PvPh5J5Q8R473xT6jT5QnDVN8EUoOramoZUBEpP9qA+UgB0LqSqg0pti
TCda7F1TGb5Eo6UnuEBLN8ic9uCjhlRA+hO9J69pVMBw2mmLnW6ln0eZO1YJC0e/
/yeelmanZAIZ4cDAFwiOZRod48ybBxZXmHhuD3KKnpouLPIb9Rtg0Xqipzqb1+Tx
PxU/3DQGKaMiZZhvLDWfJmgaRA0KxE2ajUciltn2fc2Fj3BKv/5YY/PohopFDVzc
1113RORRnxe2Y1MyEgHhQIUHrfC9QQi9ic247r06gwVg6lXP5dQpzz64wFIVzpxl
BWnK4d8cFRtQm9H41lpwePHWLs3tcgPtN+U66PWyXQOnwvc0OsKSlQyG9JM3SbhA
n4Kx+AVC78VSmw8BekIknyMxHgHnmNZUJkNbtfaVl3CqpF4idKV10PORgYAhXlWz
xOqUdYiO1eTM5GUw3zIrBlOPxYmf1bz05wDTA3K45U0v6uQDcIxkIC5OxAgqAf83
YXpTq9By9AkRgQwVxsG86NPgosD5H+klupZfu+eLU/1wZ5grC7skzG5KeR6PDrfm
U5Mefpuc6oLJENg8X4wd9XhUwHKDeGnwebMMYXRI9I23XRws8yU8VwVik7kOUxgt
RBVsqGHIrT9sICwU6x45vsLtucumTIuEeb2Ck8hE+k2iuracYLTQqlX8WWtJEAhr
Y08o7iHyuS1EI5NPjy6SRQxMD4KmnzSO6bsRTkzKwTgnW7CgepBjfKOHp5LRg0tU
f28khLlSGWnlsu5qfL25tl4MMIgrBvuzZHLRq0PsldNIEyr/V4YchPsrljDb1G2u
0jlaMc5osx+5iaYz6fdEl0RP/EnXh2+hZ2IHArL82IXOFpmmru4an5Vz+u+s+PxG
UL4WFIGuGXpaeDkkzrMQEue2+AxxVAL4Dis5I3C38A2P0TdHvLahD1imp/38PwUx
/A2dNtmDRd3rQfwpfkl7lnm3It1RPDnac0aB6SHnk9ICdPyhskHKLw4ljcVmSfci
1YNubpT7zl1IOmkxW33nUUEAFmvMCmUFAwJCbo6fkgH2Et0oHKuauefzbUOpUgey
3mwY1hE0B5iYHd01PTEjV0SDD1shtozPA8QDgYgTZU7rLO0/vlrBlvvJC8v1CZ/B
eVXDZvCv8qSFdvtgej+XJAEp1SiKe+pjimABWnDGsPzBhCH0rWIshGmT2zz1VERY
1tN7Q+16LLsYZ6U2dUWpPu/W/Cro9VNYEHHZoKy1cBwLZc59wDVVcSBCCdU5vYP8
nmAeqEffSIlGAFAOwHwcb0jkMJVUYUXKipJDD5rM8G2j2O6/Uu62Q2e6M6Z/BU4c
SoLjo+Yee6m6iqXuLCUbhvej64Tz8XJePT2C1tOjm7NVguvUV3TB5r6qNTMOQ1We
XeucM6UJV9FP638KceXR3IlOJ/DqI9Ra8G1M+YOYkCFBwgNfBBfUp/FhWujHoQWa
U5NqfepGXBBDagcHqC1hJCvY/Nyl76cTUDoWFsSegOfmlhFKG/+EfCXa6pxxCOxj
hcOPp5a+aIAKI2XvcYwE8/V5F8FnM5wE7n7IVbz6U4ubGUAeExJ46zCIMf6ihL3A
Zn0O499B2E2gsyHGkz2X9p4teXAdVXnTL8zB4Ko7KAu9k4qmnL/GZaGiC5y6q1Im
AGZ9TsUMs9QWwdYKqzWOHN5Otx37QDlDBOvTH858zw3ijYnNnYpYdkd7Pm2S/s+e
ZiMfbnnPT4QY9vSrdT5dgNLysC7CVVkmzCxQW74Gev6ca+TyZOKtXbEERGP1oW1m
L9A13uIH62jq5Z5y4PIvfSbEBS9a6SjHcs/asUy7dqDdqwogxhg9ScNH0Qm3L+Qh
U8Emp/MHJNr5yze4GkUFbWIfbqP7jg3jawfYGxH0C8laACg/3kL048g3zxZdIzfB
xT6XY4lv4faW1b7Eo1Q5/rrhywLiwhUJf9bOYi1uqRJCzLoRx1ivAXOhilxnqn4C
kNaSPfHaQb9gs/syAOsqowB05GoQCFmp0kGpHQPF6hNsjVM6SYHJ/1WcaVoPk5ys
B7njsbhhGFBBcVjRpK4rkYlEKplKdPelA2IN/ZcB/bVqMfxgMQpXJLJ6nPf497QO
gtJcxd0aW2hxEreIb3gdNqK1R9sqPoDq8BptVtKTGis/YohBXbcPeO808J9ZbGXy
4dD7gPH2Z5k0Y1/nzkG/f7xvYmZl8eNCE45fMm6kJ6lrczj2I5rDXu8NrrPoaaEw
jpfbVyauqdm/28Q7eBmU0tWBpmve9ShoOBFw/+IUTjM8UfGKkn4B1TMC8gEbllLQ
X3RPQjtYKBSYT1NuOtenHVgP8G12KmmXc/HFqBUMuo/B8sfzR9o7NWD/SRlbqf+I
6b8yqeCrL5mjM48XdR3Uh9yuHM5YLx+RkjsKUJtjAtfE4OJg2uTCc2w+49g36+d7
cz8T1Fkv4vJAfjxVCz/kYBP4QVfIf/qhE5vUl/01O3qhFsnfrpKhMVXzKXaX1vSS
hjbOvGto73IEgT/wdh8GHoRpH/LjGxVd5vL2ORZfhduYY4h/ERqKnvr410HqbAPG
NmjVPj+2mVND8t6mxnh3LfpvBGtnBv+gCrRkii4GSZkyE8te76PH2a64T3g8a6wx
LxBtp0CpzR28nRb2Zmh6cPHkfbiu7cfnQ4Am9l6/y5qRkQMrDp5O5pqKMOHST8tW
77IWHv5L6FmmtU7hU08srccC9N50hV95haYqZy1ESpBDGSZ9QNZ19aubWbmfos8I
2wJa7LZn6HahYZynzfram987b1JvJHM+xy+b/WMiC+y2A+QGj6QuUhhbyYmPZoZS
fYtEN1zlYYl6KK/zPNlLaoJ+1OHP3DxjsViY8+1FH9oD914XtBLUaBT4mLPzDMu4
0n9JxjrTK1A3DF7WW86kibhz8gkOJ4SHoduqR8LrtckTy2t7tEMTcvEwx7MlMqXK
ZucPq3yCDMeggq6jPAHVCF2LgrSQq1ASqWFfNZ+5peXJlSlEot0fT+h+oLQusmGH
aXEo/DdIcQ/psl2UiqjDT+4hf8bYsbXWrA2tAbfE/chylEVS1cS4S7QIWHplPC8H
VprlxdHEZN4h9/XTB4QvI99AOOnNoUy4+KLD0X42R5UNjGlxtzsCMn/ZY+ypgoKp
UDizCRY/o1oRYArEMUBt0X8+UbfSBHFfvzo8at9KwgWZ2Tc7TiwJ5OFHyZgCWNMD
GkP/Rxj5qkfRRjS8T98yYJykLUlt2hMrc75gRmvNNYBWf0YJbCOKpW1STQi+Ywad
obs1zDvAJaqoFsh0qnxfoePnWQE5+vP0nzMl/LswAd+xkmgWlMEHIr0HArsf3VFe
HZy/mT/k/qyrJcoBNmtHgXkKHLMG8tWwBE9HV0c8yu3ixuXa9muVrgdhDC/ywRmI
7LM48vT+snNd6aryiuvcYq5CsMrnl+0S0kNL9NTGao1ZsqIlylV/LHOiB/UpdEGH
y8uLRqw2laQvlzCqJxYhQKrVRJSNeWOaq08Mb/q8IPy8G5DEO3fNcV4S77blYGqW
xL6zMMiykOKmkLX+rQdCqg+/tZ5+PIqWHi/f8phdrvgIL+O2AuPMdkQ4xuX5YSE2
k3QyXceiV6W/Hl34UHKzRvZY/YfRHSqEyANvXEcwf7mjMHAO6mNvKp84yNgek1xp
Vi0K6Ie3XmL6FXezRcBX97uCJb9LKWXO02o9OvI3/FtkL/2xIAePqRcHafjM0ZA4
qObniKWviHYPQO6crdAOlnKZ1LC1D5to6MYJdOiMp5BlQvIM1PO2ELEMQPMnxXb7
rFcx3oHI1jE5kgtHIpxdJBuvEzPQ3Lwg4ceyQ992ToA9yn8Ci3c+SZ/Qjvdf/4nW
b8pX3gLUqlUOiTOxRhSKgM9u8qnO5QqoJugOSWtpmQ7CeHuX5WxjjPsJ82gvYiOB
sFbZpgq3c6Xzi5Ps1F+v2Na01yduaWjBR24QPObbWAXtJ7Ep4/K4S6YY004Di4Q5
2RhOff4akWFWUZqqpeRbDW59y1Prwg8G9RmQ1V2EjTiBFkDeLI7IdJAG4EWzj4CB
YNl8Z/tt2MTglRm/CEC6UJ79dmCeVuEYxHWIy3f6f3pcj3YnmRnwu7MTzbPUS58C
xsbrUcmbMirKtuG01zX9Lc3IftU4f2bcAjx7zNwhpaK8JfUkdGBBmoW6etUJHVAA
b/y3eoEgr5DLqo+YqDaXGLnoFiHFZfoLmg9GOlBUy02lxRB0CQJTi+OxiY6Wg9Z/
8ZotUmcOmymFpEag1hz8QxCCisgV/sc2prmXihdANrOQ30YIJEomXQDNP9aHXOHF
OT1MbquQTmWq/ouCvjnXl6/6qvU7i0HMIiCBdCipbU97hggtzJNpKbD+rN5hQcWk
lVbzcAquy7LbL1Qe5/7qF1hVgCt0PTODAenOdB1QvtgT2t0BS7M1ycwJGMauiGCX
Yil6J+EVGN2dZoKTpUTVBdgoyWxfok3VKmdy2HbxxLUAYcRqs7QopBHTX5CQXn65
ZPOir2toNOawt9e5BY1HdkFAzhGJmjycvlbk7PIaHLoTBUmH5Ek1NfdUFyomC1Oe
KIqv2hcCvVGg9m8V2fYH4aHaNDWSbKFkdKKREEZQxMEHsbm3uqy7YmXeaD7Hf7mu
ANXlvyy7AymigoBygj7DSbBquyuks/cLmEk6kilJrjpT2qjAlKZqKPaupY6IC80i
2DHrfLB+f6SMqIQibS9gmhNCvRObG+Cifa20fj6qdwM0UNf3X0USjdjD7NQ8z7uf
c1ME0kxYqZFfY7ojfAgFtr6w+t++vssAQnW0yE5r7cQZLOCxupQ2WTfgsmUOB+2b
ziwNugIO/yLP9422KTm4wQ6IEgx2BYHX8f+753P9+yBaxEzOJ+YwjDaa6hwbzD0z
/qZBsrub5HPgnfAWkqC4rft/7PWj/t0DugmJkqdYVkVMmQ/RwUn8tt3WK4VM0eAv
ttIDVCUjX1dgpNViadlQIszgknnTLcr1JL7prr/V02pjXdGHZvbMopdyenqmWt2M
Jc3LvG3Zxy4k9eFgaeYqjhuWylFzg1VVI1qrEQqhMuVu72yRR5I84efcWjPe/KF7
P3IRs+JgpQAcSg4TXMmCv8il0s5i44xaY9oAN+2ja4mbsdAbHm6gfdCUhis+C/4P
MJn8kI65Dp+wcY8caO4KZBKLz0Dc8Gss7NVXv14+pEXjpVZKUPnVTBYoh7Ab3Vm5
fLQVneMnNQCJGobMMcFKfGuWbeVsHmGOtpYpsEC4gO9VNn9G+69BcSG67sRk9dH7
IFtrdkfRCFLHPrmpvG/9wD0RmnGECWxNn1xJVlNscesVpDJ7wvOene80Lvxb4xSN
MpngicnwkxtrpLK6vTmubTbhbWt9biV7GS74YWp7LWHW0HjHNNNSm6d/Nvj5QWxO
wtMNp4JsbX9qfv9es8KzFJwnm52gU3IvNvxFIlZDhSAM+0/t97sVyGhdtRE4NZpD
ENv7L3EjTMQ56MsENKIs/yCa8e+l3OMMwBVy9GANWFJgWClNZv/QBuk8EhIPeZVh
bJo9FEc6Q5n4rWDWJTJTveSldEMk4XySSDn5egDFHDvKVWoSir23D1ECknTfUxgR
DRV6HLtfr5ew1eaGa2ZOa4Y7IptcV6ZTK4zcV4pG0yU9Y8cRoq3Qxc9DayDE3BCp
upYr3dPvfqyFALhCkiVZmcK+iPXuv5Qu0cGKhmErKF4oZBaum6AsfEcA7OTFLzHY
CjceRWDalQfPoDaDKVsjIKWWS+5pbwP41Ij/O1NVKDfgaJl1lKajneepNfc0pa/f
zqucNZGAWOsNLv0T0bcxyursKc7UQG54xKKzT9IAXtvGDvKw7jCne249m2Xrlpdw
nYWLljY+0tKJ+lzVG5xNxDZC91/+pmBJ1v324UZWadk1ofk4AqHSK8jrehzVy1Jy
alVw6BFrs7IvXEsN/wp3dXN6TtNB1w1uHQvz/9qWBTCmqmrrae5ZXTjX5XK1tArb
qzw4BVhHqwKeCFeMJRyA7NNR8+jJXlb6BKYeCtld8umB1iQHKr4Zcz+p4Xrmh+X+
UdRQRgjtdNtRHvneQE/Lrwl8BlfYV7xTDQGD/GN8Ovc/pgIhHqIqMVsHPQOU31cv
vdgxkaz4JcpY2fGVHjrmVjPJQew5bL9F78/fnmyh1KxIK5m86gs5RCn8GckbTG19
Vfvr2vRurAYUlpwfiKf5q+6EutYw4MTw2pUaBPb24T+kjriIFN2TQlimw7RRweF7
D/Pg/nXKpBSOsdNiOkFCigng79l4p9cwyfY1Q73wBKdf27Ox+fEw9FovaN5bskCu
zwIJqFdCC/Ev66s/LmtVm30S5ERbotl8HWYJPnLedpjr2ZlMkCgXlN/OFpUq4wmy
SvglWKAxtB3TyVBfuVoLjQ/+oafpKbojLVC0o7zWALZaUUkzbeFcIjfgUMMj6sGH
pn+FBoMz+9uRh+qTa2Tp2tnVH9/ClS8/pcOnF40rGoM1lLN4UUKAdc9UOXvIMlrn
cm4ylWbUm5bLZG0rOfA5cZLj7BkqzWxSW7l+zNcUhKiFZRWubbkikdFoe0eJty5Y
L4CHeqQZudmW6eplIavwOWQzv4FF9ruU9ti1p+K8if70uza1i5nad7w4YV0+nQhu
g2+VzLSaDfog5tCTq4c2uOB1II7+VbLwOXrfqvRv3X4zoF/jeDIEvJ0VdLnftqep
FxE/XoavglTb2vAnSF+NwOzDOlR7SZTHMYexYyqSvW8gaa7ZX7+1pDOvX0vnA7r8
21zFQ4AAJvtN3BxyT9Tp6wuVG+dc6IgkIa7gVtfpCfhPNGN6YI8N5/IJVupnlBHH
Pf3DIoHpqDVvUXOpfJg+7oZzElkCsnVvDeryVRJ6/tDS182DDlGB/BZh/HkBGtrd
VnWwxI3qtrw7ldTpVWrtYWqd9Zh9yOlIMgyJfVl02Z5pw84lr1f+CeuktPzCapDu
TciyIEIx0XxK4LwDamPqb/j61GdmxqaSQ/GK9iN7y6//BmZT86fHEvsY8AD1TmyG
TrD6a5mmPW+WnBETy3wEADgY1os9JxQJsv4j6ktTfa9Jh43EnnN+S6D6kP0SqkRT
wS5lKjknCNfweU+Oj2a2CoVQCC8UhhTlnoLZu/Y89c+83Ak8cYUfyQYaHjt1dnjw
EfWGBnIBcDZw8cxm+BKxBeQBeRPoK6hP97sT7isQFgi8PUo5OZx9pByzVMzsCg2j
/Yz/1gfCcqVuDErWHpHLyoguD3sB2DVkqczQIut95d7JzBs3lTyXFhO9X1pzvW5A
dn+dIlD9Pk6LrOXrvH4GM8v8uC2rHo7fpxKS0OltbsuDMxi9/X6visoMrhIm4ZJv
EYTgXY7RwPKh8V9LjqtzKvnElSRKdrxYKoIM2lU8YqUPoUMkPXEyLru8tM1o0NOG
mTIdwUDnVfjj6Pm8nZfboIovba/BMV7YS07mVfSXSIQ1P/3GIShlx6OCPa57xtrz
Z17OI3fMDlW8Ew5FPXcn7ouOy210BFLm+uz1cNC/MFYe5FDJFxwWNNgvrn7w9OTk
HfPYZvbaSxc6JsN83Vi64uaPd2j+R/leuYd8wfZO70oQqddP5jbgb8GyVLcbggMN
9gpi01oDypQXi4mo59tl3OEWrVy7vzKj0f18xyACsoezClpZj2CHpDPzwR1qXyvZ
8PsHWegkN5kpt6etGs8ZWH7YhaGbU2GECIi5emjS8KYceGAgCN76lPTCJct51Vue
A8KIOVnX6Zw4VXd9u0sytWACuD6Ljltkjl3ZJzBexxJsb7pZ8gjAVrEFusKYiAnE
cYShEd556PuSGMHQLtcKYAuiadCwWhDSP4BDMFiEiS7CUiN6cNqkqd2bSRTZF8tq
+TkE+epR9PbdIxro3aaSKxw/jhXXT0tbemheAUN0tJ9U6bIWMPhOCzWGbBBS0JTa
1vxIek8LdVPhgdaK0tVkzdY3DGu6vpOJnl0Oyq4XW84Qj76VJSuKk29LglDgM0La
TPvwLcrggzXFwwIUvwrl29Mx98TYWL9rmzITX4KLP/1wEE9cmXb6r7oPaf4efV+W
VjshCPydhPydd02Nu0Ks2/NQsnv1Ssg0LGHWXfKUWPlUAB7TDZPoluLR+T4I1y2w
9K5oIg0o+xPApfYHE8M1cLFhn17+DvvZ8t5po1ZtbUkxvY9uIzywVgbgkrxAXf7n
ajacNPZBgmolVvHA83dO8vV6B+xjjjlVAkMi4jCJlum40IC0LfXOpSNHCy3SKBE5
fgpV4bXKlw8atppEz6YC1I/Sh+jUE9ho6do48URT6MXWPHnSaviZOWs6XCD+4eRx
SNusdhNzcAhas1Jec9dNZFWM6aU9abLRGnMdsQmln89UwS9qCcM6+Ock7e45SC+0
oCKBZ+H3iJRBEoVRrpMLurqnE+Vsmql3Fb5ehgv10U29bvauQRWF1x29iG2kk+qA
pa4YthVpgSZsNet1FJ/iCD1sSxmxY1UqP2r+RkefjxcubJ40nEuNXo0vkuDnCIlj
sI+JSn8TQCgLRty9r8T90ynR8XYvCNJ9VNDdol4RswZciF06sDud2ejzJS0UdmG8
c45li7WseZoYbrvSo5B1tikm4IwM12eV+GFbrW8f+yimbwG2CO4MZ+a1cKnVS++D
RelJzMK/nK+2ow2Vr4M6FtPR80Tkz6qEhfxFmBvsSftF46v8YooXYpGvSdn+UsjY
V5tqVhoMu9RL9wc/D8XqP4TNFsw/4WWZj7TMcyPLPsKoafWHTyqYM4mx9xYUyg6X
AUnqjMsgecacdZt1hpkAUbxZfKmsRk152INSsB4IMEF8uM8onCzHO6MDlX2RW5fX
ipwn7jeMfa3jUjVRhcQzpEV1xtYCwi+ys/QNepJlxNMEnCPZ1nrdgU6PdN2KNUMs
WOy+tJO7hQl3nuz5Rwwb/t/DOf+eU+wupV1dkuRxx4ZnhsYk2xm9v9Y6qpH1hsd7
3H6K4RwXFGLloiHBOyexV1r07+FWhfyjt+1jHS4f4gcP38nrhHrQm2RofE1oIJ8J
bp9lk4Fe+UQotbJTOTD5MZ8SFjwp+KYWkLo+0FJrhCmpRtl9yLzewHeK906IbnRf
VWBusnVyqHXu/9uy2kTyAa7NkIwygTJAz0izSNMAvWUcw8hNFyZemBFdTjy00CM+
lob+qR/DcTNsEjjmFpeH2s+QoS4CqZIF0jXl6xCS2eFJOTnbdcnAKZr2rvqBrQMC
PI+UGWn1jmdFJDwoAZ8KSOVfnWhGm/EbwVXzMr+zZlxfZfau60B2I29osvWUtvvi
qhXw4LOS5H0t5B0nyIfPCff04IXlWsjewKAriG9StVd1uwS2dmz7pGDUV7Qpgil3
Z3famUQGpz5tby6nzn7UG/hWTi/g+VN3r6Yvfmz0hWEx7xmJwEkS7X5ZiK/fNwvV
uCy5Fe4maocpH+EEgj38BEF4HHPkQ1GqFzDNoJU6OrtmsQ4orMycbU15BMWVacLc
gCfvBnmphUSx42uRhdmaTv1hR6Q33HxrgRJvwTBTh3Gz89Art7xIt1j04J1j3mz5
7Md4T+MrPJsYNwErLcG0rG+jP69mX8zvzB7ZB3WSeZBR0+haKUbxeiz2GEfo+p7K
+L3HqgjXqHxJG7TcPDJi23FnIcHp3sqBWMZwkfiuCYiqyaPZF5GXj9MbZcc1xxOQ
g8tTFSoCLa++vMxsSWafo/sAGUKXsLAQy9ie2MTxEuQm63jAynJW/QrMeQq/VIsk
lhSyy047pxL4XIo/WC27NQyljL40YT5x7Gw/Y5cT8w28zVkr1dqzMSRef4ImBoAw
SHJfxI3yJPSD7miEiQa/drVTFqqC0id7QwIpYqxWTe7l+zGpXqs4mJyXuxw/r7dQ
XQ3YCvY3mJBg0OSTvQlEMFeXvipL460w9XXya7l/++x23ZkXZePeiQZDJBTG232B
g0YhwtNySGGycJoNq9PPQ+Sz/2V6Q2zQ99kjQWW5VgXFh6dh0EFuStz5Bj13X3sm
swTjYbLPWN6iqLWa6rucZ7NfMTVtHXQd2p3Ge+qM+xNYFUpFjVTpDjif3xRZYA9/
W9bOynB7c9gXFdFf62SN5Gn4fn9LjD7rhHlFWukauiaUETgTP1T8CUrQwW43JXTr
jqhDvoC3hjd4DI2r6I/6MSbNQhYHI6jVq8SkkQlD8C9GOnuczOWyl0Y4ksyrJcZW
qCEhFYQrPf3uih2IeTWoZ1ft7IvnEopBtUyIaRLpqNfPOVTH0X4vT1zOg08loTX9
6iWca2Kz+u+xZmats2oVL6fTofy73jiMhdLfoiTgCRd5VEdNF5iIIKEVw0ScKBEW
bW/79XmK8cWCbLQsEOQITOBNrcaWP+Qp/IqK+UUqW8NvWG7eA/tJm9fw8TvSH7MZ
aUr1WNU1zkRAs+O6uKAFbc8VPN0vL9ACvf/hXpZr5JHwQ0qLH5Xs1gzuLyQN6DIG
6PQ1VtM/+eEAZZOo13b9wcAD2dLT31dfHLroQ7zL6+iqpY+jXi/Pt/plxmU1YLWH
SzsZZdoFR+Tc4d2sQCf+kc4HICOB21utikr/WRJZzuo5LGoW/M2Vf7doek8M755A
Ma28zEseN5NSrYsIGSzMvHcnv8KMNfpwBF1bKneS2vvx22uaEZ5dHlMc/bM+VI0U
RPNm6/+2IVzclOqNnN6UiQxrBsdZDy4qnx9477ayz0ZnNtOVQG6O8lv3p7y/ys9n
maClDLgc8tPuAM/cgyShxt6uNuK8MNqgHurwJ7XE9E/xL697x9L0xXjHLofpyRvA
1z5WBHHCk4jaC3PBGSJ1hfip5hqTjhVR6J++YgBe7L5YAd56xB+yVqHJf35Q3q69
4bXlD0kDO/1XsKunFIaRPUNdnSDQFmqmasNuSsfon8qlRgEXIhJphgtPg+O+nGqN
ho2+pL7UpCMDPVu0Am4exzBXpCIXbr0PNTJCLiPSv3/8xUfVzVU363IiAAd+du2v
GHcg08zafsAz3E7ZV5gl+mo3ntLT4Z1d4V2OW0/yllyz5CCmszpfXkudxvGptN5V
oeUJ69BvWCT0al0yOhdagf+D5GjW5DzePeY0wu5mFiEjXe6edxVTDI76iAOxEero
sDn1q7nPBm/jZS8DY4KhfRL22p6ODPXUxxiEexpUltivGSxX80hOwc7fBj32JtYz
Fo/zkbCT3bWV+Vw4z1pCS09BY7ZxNjGh18RJDhxXsCt+zUrBQ79JWKzRAPjugdob
j1RjkUuSMACflazedLRxClMeXsz7mlbRp4AaLjLQRF7uafGWrUfpG4+xM4UFdHPI
GKSpDF6Fe1ZnAXuhGtb5WyGasSvUWdlA/X5ReDRSIcHmNoDqoExS5uvWN8dB81Wf
NJk/KTx9Twhwddjr8hL/xnxwaQMgjtyEUdtCeZ1FaSR3+WQQjEhjBA3+juWBiErG
1F2lyabs7QPZEM+Cvwmkw0ulWQgQZrjHQdG1YsolYqt0fN0M/7LYBLZicgvKPnrW
fpWwfQXu8nrVSHLzJtfS368zvdpumvTI3CTHMuC7Qx82BuqpjaC9M8P/rfFO39bQ
PkljsPwTnDFb3h24IewA61BfQiBClfSzUEHnSUSkccKiYS+dQTh1+7npAbumKv6U
iLNnrSeQooV7YSpcEl/GDhUaWlg1hwlYLo0WimqYge3gWi0ODzwruPkz8zs2gi3H
LQoqrU26prICEpaQlFuQGlIP0SDIUtqivTlkx1g+a9rvlS4bdqXqQOYBNyFo9iqs
I73Eaz1Ag5e5L+mEcMGUq5Hk0tI7piqXK6q2f/pWiMHTuNTlZZpkH0WNV9jYjPtP
HXnbKymoBMZIR3wKLC8O/hvL8R70k8zslZ9tp9BbG1KjDrLYKxYFiWKRqRLfsnLc
EV7h4Xk05C7SU/8ihQA40v+E2ROkTVbGHldoDR7OF8t5a3BuZfoo14PyhDT1l2D8
JN6D+sKkuV/ZsIWAex7ntqcS/E5FfQeDNnhAxMI7lIBSXiBekv47nmK7zm9TWIID
hAat1IPRivT7LXpQz/r42cdmG2cpPcUj+9fMZxOFnVMNmGxbjmRMk/zXf7jqAbpb
PPzyBWLAJX8YjRfiDj6Kj1Vbg0CCpmZupoUKCWr61QkoLJe8gBnf16ekgIFao75j
Z8ss8hclU422EQCosAODyyEsP4Y3SBHFCfpMwpqZu1jWenWobb+K8/V07bNxR6wB
6Oq2hn85Ib0ljKzcLnYgdslsfCbZwwvqAFhi7i0v9oC/rF9G+CwmXJDU1TDRVs2Y
gjoozmNyELZjg92GlHVmVQ7WyIE8G+7D2a5HyqqlLr/fGYbjU3gEcykKM8j91rOv
p/By7u8R5qfXDVJZrAfyzrWshUfWKXB/aofTUCzRwVRADIPiR4iJr6oBnxFcV8Bo
U5236e0cHGeVB09bHvkeMm4OW8MEAdCUhkbGjNF4zaxJf7H4ZROkRQZE3D/AsgNu
yV1PDPAoXL8I3RnRG89p6i0o17qroJK/5l9AP48IiHu6QyP/B1DByXncr71QPM+c
UcSZmIRxLunT48En6D0yQrBxs0j+qcvpZSGPQbPBupMVA3CyWkq2QKVq3HJdNXuH
ZIsB3UMrfQhvKWNRHt77MW/SR4/bBsTw40GflDW+5eMeaRxZADY9ndaKgf0JmKMD
g4jIWVbzD+Zi6ujj91s1+N6MWf/htQcU/oRsVokwSBq1B4w4FKAGYOGfsZ/Rj6Bb
3mgcr6Dv6WqxfzhIexP73+PAn7uHitKdz5rQjaC6mnrX9DaZJNey3dVGeNEURQxu
XBnb8RVxgHk9Wn2epaf2yewDkIv12rD6iIGoWOIlJH0h7DFbVbL55eiflculgsFi
SrNAyeTWL6Do4I++9mN+ba65MH3RscJQAhzG7jiU8ce1tGySW0UVU2tanfar5A3x
Yo301Kde+9tBLANWKrkIzL9eVDqqsVsy/TXVNIoCOJXtGLud/LIAeLK8mUpRHUj8
1k2HMcv03QP+uA7ZGGqJDvFPlG+zPYxB2kcHvrEzRDjCK9tYEURQVqtRVnvl1MDY
Dqvpeg3US9OBTb0c/a8/BYq4V+6pPmLxRg/F1zVzvIKQgn7V0RXTrZdAvrXgA6HQ
tH/xNFgngJwocbc/9OlinQqobMSzobSMpXUTNJQvkwPLx3Eorig4QTvSkTbWi0ev
jY86lRxxFiO6pr0kxYSjT5Fjc9OESipcOvdWwaplcGqqS8bHxc6AVAZxvrLkoan/
pKa9Ie8bwcuHwYw2XfcgjjUsndCgyS2cpvh83zciL0FJMyucHLVxFPgp806RUKEL
yCIS1N1UDXI5HwC9p5boOoC2N79p5id8Fn8WfPYflZ0F8wQrJJk2Fo1y1b2xbPoD
ng/nb64i3UQEE5kGls1t7dOSxIJ2JDf/FJ+b25AjSdDQwbEOH337um3IQOFyCL28
XdVi0Jv5Aoe15vLYjLQShnQrhLapN+E/RDWOE0j4glreK6Nd36BveDhc4whveHNs
EhtCQMxlm3JNylptoDq05GMbADot8pGz7pXfhX5nBPfPR4PWefQEmmXeYVKJItIu
9EDBYxMqcn2B0mXJj8TS6Zs8W38AB7tzgFew3SCW8s9kpWE67ld4hKY5txSOkaCq
Rh9ubEun6yef+6Amq64wWMz9QtbdyeNowcocXRdyMAt+siTnVRIyYkSpgIWEqErP
SMkL7POsEjpA8/RjMqMslsP9ZMfMLfPlnbux8/FctcMw4LrNRqkSY0YE76kjbatV
FqPsDwFmMAKypSNuzObmVAdLAkHNqGUY0ZP8WMQCjWoANM/H1t0f8gvVQ0FrSMI4
jdJldWLUok3eV3ksuEgPR1KkQUNr/P8aoSgrUvMt4XzW7A9sGeNespLMMVMm/zjI
xhMtqhxZADKeCx45pDf3c2b3P+PTJQlbbNO5k5Uxl6j8Hnj2hbZUjOdTR5IhMqIH
Xzka5LDSdLc4bAepbqhq4MHf1ssHq6N0ezEmPWssjVD+VSqiNoy+4RrFdjsNxALM
OQ59W475CSwd+lN01UvSiCXb2tEkZuvVcZLu81QB/xACF2IqVQ3ImTeT/zFLHzIx
e6cddyKZTGAZfVf7HWrSml4CwMYJahSm7VwAc9/ri4kKAnQFgyyT7MXowNRgyg+S
d8pcD5xNyD+HKMQ3e6i8eXZjlWi60OIaBv4hC4O20HphyTpT2Syplamkgahj7Fj9
tgpzvka5dRpCXEZ9q0KjM0AWd/i8NWwzzQWVa4wuaNop7j7zK4YaaFNTYnQq+5U0
wPZjbOPr8Eg68l13rOuBDfUqmMIr3zQ6E0kuECSoaVLayrzYi/OxMJPZyLMBbwVd
7y+eq0fyMb67nXmGXRzUwo20En8Am6lrx5lFM8sRCdrvllRfUgQll4Ph/Uw+06dy
7hfTTvb9c843eHLak6+aU8AwUfxrT7PyQtpC8gxcIRmoGShGv4GDkGGCeUVjXHUf
XOffcewtjoRzxeMAc83BufmVG2skk93nmRVHECJKqhEs+T0S837pS7caVhmLLOxx
M32Bs/ykit95NM1HD2uxGtZCeoJItp7BVpyjXqedHHlZJbM+J+l2I6/Nytqvpon3
QZwt5a8QMSzWvUbmhyLmcCsS6q/Inz+I2yQ8kN66asI+3JaSiYn+K2gD8pVKIx/O
+vqlLOKfF72kunLnh7U2sOtP2YdVSe7hgUvQj9lhZq+yqIp2fC3iYFJxdi/9+zbR
q8A8k3M2cRuBB5uSvG0O0U63O0BvlCC11f4Z2QOWf6k83FgTuxZWUDYFpE1ekCpf
cP5SvFls1qDZh5JbNtuA1ZifGf7+tGF+KRSXWm+ltqeXBGZaSbHlDaAfBAa002Q6
wMvF0QSs5UdR0RvoTrUQh8xOs7TM5iTOMWdhoYt5zadMh2N96sEwMIW03jUMYMSN
b6A0Mk2+0Un3I4wejzCJnxrrOFgY1D1GE3WiWLWkHlvye4hqWeLVtNSkVmb4APlF
1yHQ3eu/3UxArK0ffR9YifMMkalocQQNKrvjJuk7pQrc04fur6+ilWtPuUWZE6L+
ldyGgIPQlghds+z28eAVbwoe57c8p1Z+DJHxOuebpCIACjalU2z5nI2B89vGPylG
msmck32briU/mjcdW+R6YnY5l/mh4nBMDWlSO1uMdii8qd57+9TYu4IQNLV5dUZf
reCdi6I8KwxbSZQRpz9NCtNhTr174uid2kXYlc70ZD3j+JDj7efUGTHEvzsebaMr
VHDFd40NjgWLjn0D0XrexdDAdOXxPzHpoN+ickUMWvehZgvibXOm/yJJ29PP8ab4
u8O6fCaNEFwsgWMOnxoZYL0AhK8YFxUMLE1eUek4aYybSYzJrtKi/IZ49iaQv8/M
h1IFnRH1QffVPeFdHL0IizgynVK8zn7LFAIHRLR3ikUG4rhKbCed1aVxQtpqFIF5
skDyKZCHoajTA6R8Ir7xj1FW45E7yf1lA0s8Hbuk0SxDSsqqUoDTV4BCgYteNE7h
FLKXQyxn/8w5oUcEC3aFTNB4gf+EzX1s3nWw09GVQBOFWdCLaxu9bANwHKM0z8Ea
Ye4/uHqqqz/UB1C/uKMDcl6FKU/7/Z+sOHylPMvxA7N6dj2RwipBRxgRrvpc8vUC
szfCOWcR7yeFL+TSAq2ZnCFkIfin6qS/uIceEsA95YlSyl4QlcORGW8kf5+WomCm
x2oi6l9mCzA0168ApQp3DU+sdKAH5cGk8Uxdzw5tGWCjWjxko2c/KT/uSbRy/eQW
ywWwJIZYnC9t1iH+lRpHNIZTzwRalDUUAXYBHPMzBqE6UjYG3bJC+s7Pdis4vS7X
hS/rnA3vNeNZeaSVrZUltmooMIRgFwI1oPzvlBoQ1lbDJGvzJhglkQxDxIjlQb9D
dj5RT5o4sWNC63tKq2EuaZYqQMXjuIY9B0cuURGuQVFaYEYVuExKLRK6dP+SApvA
M9l1ZcCk5TO0g88cnEe0UQKxHAWu3jDhheWCDwiBd+0cBo7kpA0nuwn0smUgYJh+
CfPdpjAHiby2o9DvLBBOzWQqFB+l+R+KRBXHP+WjFJUjjmMKYLw9QZDDLATD0mjP
C4u2P/0312uiDxXZYcRk+H4WgE6s0dAsOc0FFgqnROz1qWSbxkw2ioPr4EHHaI5E
pYUb9TqcIO+EbhgRbfIVA100ViEz4bi4toomkcaM1noF8J/FAHtNzkPcDZwSbgpC
uHTpIgAMbJH3Ct23GP3RmHlf3qE2lnFSkx8td+ghZGciv7SwcLsuiVK8L3lFPhRZ
Rn/T6YDUb5vTd6zkv+/jPD5mN1ByCdjWV0CkE6ynFQLzAbsOG30zvAuEVVxggbT/
/IIULBzeY/3oJkYt8prugkh/kaucvELni8KGXpLEaUAkB4zFFTGuI33CguuKnxOr
mHVrIDVPdrp6KI3nLay+c/7U6B9VDd3SSBC8g+mrxNxoYdH+RBVGx/yD9XBwdIlW
nmbf1zF0hPgcMvWbGMSVfCeQne1Z7eaPE+V8t4gcCVT86G7xQIOVNJeDyIsnNAj4
WLidNSLzfLwccbSM4Df1+RjOL9Da0TDQbieOxG9NiKpxCXWxB6uzO0d6n1uCqlJk
73w0aJzoKGvnJL57piljYoiJ+o4LwEYG7tEUdQD/r5c88OJiI5QuPMJmoWzvXRBk
QHa9oChCVBmdiW774sjnIpOKfyjrDgd3VeNmxPryi5rZSo70g52kzK8ipeTU0303
hmN5zKDE9yIB1LdrxIU2iwc05BMhEDbF5cPSIdm5jXf0sx5Tp8MESXo+UFdsouWd
uRhADA+r7PnqUxZUHpHMKsthfwqb+x16WW5xTCZZo1Qh6KRvuc99w6Mg1JHtJFkx
l/gSzuq5L1CYsPx8S26BvzPrPU0r01Os2PssAP3KDNQmiCQplJwVBA8Vv1GKpMXQ
yFaASx5nzcXMpVpxx/8d8tcucmbvq6qBCEq/f3ZsI4JUr+9wQvml94ErSwd1ciyc
ef0ivbEM04ZG9hft6hqRqJo8iB3Igfq2pWfMcrye0vU527M4Iw74a26xoOgK0YRi
T9VbmgEENcPJb/6cDTNPvUB4oo4d6oXRAdKi1/Ejvf1GDomn8qv1YwMwkdYKMmHx
pohhI4AQSjgVawpL27i0wHgDxrYMZLQKOoxQoj7JyZ+4p+JTqxyODgFAkNCpeE6a
iGUmFJtQiDmNehXPNRCpP68GuoZotEP5slrer8izj+UmlnodccEcpgv8ec0MyTL8
jwHVx1baj26sYdcEaARIHaeAEbJ2Pf9Gt+PYWkc9XVTkD/su5Fjsm6O07Ey2IbAk
HfqFPyGz/abAf9U32urccl1pw6BZXCkB2pWuDE4MLC4RkwpCYhU9/ex9fPioiRc5
x9eQZFhMK7Rc9ltlGPXn+mlqK4VwSzRPyiSKWo0qljeZvLHMkVOfpZOo3zczerDw
B/ZDGqoV3e18eXNfdLGRZh+LMzEYlHD1dXpQxuc8PnhGbeCZbcO8/hCOTNfoHiGP
8GHO98zy5TELhm3qxcOM+eE0VL1zHa7S/VIWLu7FPNuGW7Amtj2PZJndamuv8LqL
Hg8iKIxwn2MVk+js5TWq9kaLZpfyw8iYT2uomAikom2PD5/lvQelKD+wTzFHK+e6
cJxPFt9nw09hxlqEdg49bEZROy+Iunswe+xaZQhzPuvsiBXc1yEjymV4a3vHQ0Z0
MWokOALcO81IWc8wB2OEXSnC/WAzoFyNWp+HlbpL9Oz/Hc/qi3+Vt3zLrykqdj3U
CrUOZYwiKEWizKf+YPk6oLktR6BXY0JQZZ5AENMeE4yrgPaiXnHxbHvIRU9GimZx
Obxt1iCKdxJtG4ZF76khbEetXltF0GarZfUq/Ka3zHRck799Pu+ZQc1RhSMzhc9Z
tu8+fTfzX6VALCLWbbW+XjaYs/jAMHDnIAURGCzl0b0DZS7GBfK/KkCzbQh+nGsa
zroexwQA7T8JAus0tuLuofc1Hr9z0jWfR7i2izsTO4tP++ZtUra1EHrn24Ak1Vrd
16n5v1kUVK/+7AObS4h3ETzlfvYkudgOfA/BgXb2qjeF7QN2EDA6a070zRZ/aAtD
KqRfH14nZWEsQgewqCxU+yw9inBcV/x4a0hkCtiQ7+eOThyOYasMyFhcFr7/7mc1
WVTCLBtiWYP3RmavDC7avr+2wb8w8y+7y4Fz5R9nhixTDVzBNJ8TZUjeFFi9H9cE
ro8pXOmqMWAt/+zbJDAbZLV+siyY76Dsuf9M+KPzdLbEsd2egS4S4e4GKnn3kymM
cW1hNhUsRnQzOCA7ZUY0tFFACzNPLA/EGKCcDG5VjbE3BkbaR9QRdMuV1rhCifZY
+qkYMrI+ixp0MG4x00VUUf9L2AocQQbWuFAJZuCQDF0DGK44a2uRFdAj+QC3gXu8
lURFNgBuvaYZm8m3dbhR+cCjhVhu/wHRzTU071LiDye7rTk59CHxyXLtYBwJhnWG
07yyam9q4m0pjXwahwMIjfmRBXwhNpwwFYBirbPi4E1iCiaOA708Jk8d0IX8HO8b
VrmmY75/YkGkkWI1F119nPHWK4zSzVJ/lftYf4G4Mu2iNbT3MmzdGUorlFa0n5YS
ru/tUoJOozC0XF76aXLPzE3Hbhx0vHXffTkINYG7kscIoB1cUolz1jZAhHTori5l
Da5/+UzAMh7SgnacQTBmzzOkHK1KqSWtU1UdqY2dJ8Erur7RQeKF/SoTYBHem/8G
5fmgxezHfsncE9yfVxpxtSftw3gYyxwpHp7HIzVZWpwPUzWbm2l1dzNpvSuS5iX5
tTu4TGOyRAHQ2vu0SAFJSVTEPln5VVJtnXJmohJRnxYEkTQJ9U+6lDphd9QOsWwz
JNHh4EML1U4wwq+c1zFdI7GXvUNKfW+tDIVka40qoLRSHOLG/D9ul8CUCx37iz7R
JfkdXICgRSr9ZilpeQUm/6nzCaxGKOUrbq3+q+uJe+ehcAm1hUMzcYIaujbeyFZe
sXus32UhzPK3heFVRET2rc8NkJB1YGl9D4sD7h5LVQ7EiLjDeHf8wYYY0+PxUJtk
DrDV3scfD5fJvyCJwrdqlkAp5prysIIg3PSUqDS/PSp25TSgxlLQTfhvaQQxmAFD
ZXl0WRB/OIBeRsHTb4/Wj6lOavYyHvcAOyoSXQSqS8Va/fwGsiXe6Wuuqg+PCNGm
1ApCRvSIAT5jUed3J8uchce2BEyThEhsPemh1j60x/pcxHGdVYEdyjwUUsdBiQgQ
iiDOFXeRGpQC2Pn5+5ZFfhRlEVQIv8lFIhY3Vh7oFLVTeXYtGENycLwV0xIjc/TO
gJmNUn/i3kpalqd55TmlHz0CzdUCUVuRygO0c9lcqJ9/6mNDewBFN0FF+FflJ+jW
KbU6dW7lu/QAv3uPjg/vq/uhiExZhredOuMYYv57VQxCpadSMQ1YWJ88Fi/hs2DL
8Oj84EoJtritPr1HU6CU+b5ma8CGi9SRkrOfl74oom3j/jOhe95Y5M7hpzkHyHHy
Moh/k03tLQdZlWQUWDN6NJ6Bsp4euv402ko0UeihV6Yt9wK9F1y3DujieTawghDo
DE3axUXeFHSSmY37f5SvlYkkb/6XbVDXHFkMP4pJDvkY9o2tKOTqBNyLKYSoJ2hQ
obx9VoNpyxYdEm67j8ufnkedyCDimJdj6qTBdObkkRBAISxG0OjnfdjIpIdsueCn
7Wvkt1IrPml6MtX0Fe+bYBxU9M8ZHqYL7nynlusGHyciGrZ7J9Ckd91YM+MB6VJq
OQcHp+E0yqw5D0FSQB0/dl3lhEx5hQjTP67FhHtbIu2MmGcIrvuXOIsNGffL2GCC
SJ+giEOSFeEfbYD9X0ll5OTq4tq714ndir3h83NFGJUbo4RDodvv+NbJJIlR+SjP
TEsLHonWeyt4irpKbN2SrtX0+UWLL50gG3FdzdayWXGskDypmKop4+0FGADuSIUf
W225528QqupqBfoU7ovZ2i8BmsdMrGFAVNCokMpl6CCXxBsr/9Cpx6QEfGxu8FEE
RjgRQZh9HjZBqjsbJAa2+CcyKuXBvWJHHSmQE8Wi1Z9RzEhQF0+mvQ6gfxBoGls0
Q+ApZkSmdJNzZyrUygaUSoCs2jue/Lcwkv4Cud/ACH0RFURdfzACg99zjRPQFIEH
XF2id+madQ/KtpjMBCPQGjBEhcTwi6Y+2E/dSKqQ9oUK3TyWLt62SA4ILoFxaIDW
1i4qI0z6drnZvbxVAi7lvbccwewA+vPrLJbgVfZRapi5XoulzptWiialpx8Unoyc
zbVNrdpmphFiAkRKDQgW5BQTglhLMP13k9yptaGSBBlEU3Qcrc30ipZEai7l5rIs
ZfolFbd6daqx6+wOItddS2KaUEuQLCIsiiw0k8kz9lhoXUgsQEpglY0Uchg6QBU+
SLlTC/GSi2JaTZ3ObXATX+EEjA28EJnz1anMX7lX9Xgtfz7VRRS+wc2x2raAi5pw
Hvz3cZYrWkhUGCn560mC+ox/BO/oYUMzV4lC+OO0pxfxzJVKJ1wh51u2R17DyukA
TGO+MFxQv0a8TnE9IEPtNTh0nSIrrEgs+u6u5M03o9u3lDThdXTfYDryBhSO3wlv
acSDXyFmG0qQ2o1FBnbQp1plURn42pDtlmNvu3STyggXOUrZU8SGeEcLbgRmYdd5
Yfodv+6MANd6ynweMnTvRJXHsBVGNTtPn1uF94PoTMcjkyFjM4XslSeeXtb8omnq
/x2XXMtaVjU16KOFqjTRz7slI4maTAxnmRvZ3dZvkIoqAxdmer0tvNTOgZwZ1bYB
eBuToxfWr4EEP08L6p1tOxEPRHQ7wchnJnGAdACrw0ow8iTEFi6lhApUEHQhcHzz
vaRRTdibRHHX0nNtHLSB1MLGSub1TDVJzKTQKjMS3VgjOzVEHEIWk4gWdrJgCdmS
HIk5k5OWsYMWhP7IL58/eI+7mJFcV/qN1IDPiQml7V8/erHh/+pbrA7VJUDYWQps
uZ+lmbBWl5r20cVp2lBaFBatRwbM2hx8mcsoipcUDWmKhuKzQI8QYCEy43PfdEH1
CfC4V4207k3GZ8O9RqwI5kvM3leftrLnOItEDwnXz0ABrvXuuB2GZKDs6y7pg+DS
Ob9WVN/6c7IWiGs+ZXC4ldb1rRsTWgpcyzDM5tJbx3693ejAt0F/xMPvMrWsLQ+x
+LgS+cW48LDzUXJrBXjcBL4UxFvGPq6umPFgRartGK6qitIFBRWw4GtpYyEIe7UX
U6iAYHDT6eHyY+8KnTfPmT4aBEssW6UD9IfAnVjL9QQau8km5Z2Fhje/YLNC4E46
/KLRSkGR+lYhw9hmVN5tGN03SErDELMieY+Iz434k8SkiBd4NJHxHCNXZiTUpBk6
AUmeQ/nIbVfbXhByBwoCW7JK7vjbthLYdXuffecYINA+bR5+j1SWTYEoqgrPfmQp
TEymppralFkhTfU6jW4GPR1IUuHzL1LNlyrkkoqJbqF30vka5gUj3R/eKsA20Ykj
8zX27mrLuFwxT67YrX2nVQRGct7R59ViGWrtUeFl4fqbRxNzAbi96w094yzYcu8M
uw/ly+kB+05bymjNl+nrCPOuUf7PtXDnxQXg3prqB6azhbzeOHQrNyGZ6aSt7rzX
GdN6Sz1NFeE2mytf1spo5CyXrVZUVn31J0R3YgalZuIhGO3kE+pAf6/KKDKIdtqV
boN1vgkoZcIRogbeMq0ehOQjwbLRoBCRveYnzrAdlQy2TPhDzZsyuQPgYO7KXphr
lL5BGQzDvCHx8hLXfU/j3To4/Zc1T8PILsGCsHXKbpxF6Ten0+5BsaYA78p94APm
LHB9NJ+MngIQAuv9f3gEOF5BVkbp496tjOjc4FD+wHa/WNrxznqgh+RzCWl/yzvN
hkuBEkXBZSokFiAeS7ZfbcN8FRtN8ypfaxTJW0xtsY8rHtNj7CfKrihw+xGeGVFJ
OFguk+/rk/fTrP2RqVf3K90pRvY6cUHZYIc8uGzxtjmjeQcG+hvshJvz2xmeSKS9
6VLPgxBd1tCM6Axurg4oAXWeLhZ0JkQxNEjUKIzjJwZPbe0pJFwp4L98f+oGGLee
taY8y751DK++OPUjEMLA7E+4bAWaN0jn6m5q7HrJh51nQPczx7749nIrTcVtPhIt
M/4Gx7Vwmg4jgcieFoepmm44U35kvz+Tl6bwb8/uT/JDRBcCXPNs89Cp7pp0INDQ
fTix40bULeU9uNNOkVfI1bqRpMTm2Mfyihqb0Ser2iwVPeooqjSsknn3jqcPOQ2d
GwmhNeLp26s1jgJlVSNKOK8p4QFNpqbaT9Y3T7Vr0XBtaL/x3eBUb3/3o3fYBGP8
s3u0CPyX62TrKlhHtszhE1yML7cOzM5cvDNbtNLVBYL1pdtpqLDNN/n5s2PKhevM
GzrqrPC1vHJ81gTa6i6g3QWOk/lqnAwEBWNU4fFlJCtIaxqJsLWkgBVQmWNcfDtD
NWXpNussvrARkTSl6z5ljahmKERAGZli9v9LfMnh5TjJLLbODQLSThrrLgsqXFhZ
tnXpx2Kx0OOu3G4iAKvt9T6Xe61Q/UI2qf2EMwYW1LizOPGZW02Ln1+J9ed/2g/U
frbGGzA5YwzCvfFrIq4vyy/htvQExz38e984Z9ZM8n/vx1Ml1rLYlrdWUs2m6XGt
fS0VBQhsQ0N++VJr7nBcIVJOECqdKmptQPQ2GVid59Pm1uZ1EOEmuwXRv8IIYbq0
UeLMPURunCXDrBBWDRDTedHfPfO3pE8I4Li3xd60qYwUOo3+uW/dluoZ588FyKQy
fAORnViBrOqu81coiZJgxlmfLwagIiEGQKRAEyMla1r8g/FgY3YHzqmowmhbXt9+
zbYq2t1lK1JMkGGva3LWPkxUdS0KTajoLlh3jhq4WxHPhu0Ddxf59xIrfJtG/nmP
WtuFGyGvX6SC0920n1pvs50m6dud7XXgRm4FyEngYJTR/Km2Oua5lWN7fMWZK6gO
aYSRwVrAJg02m0ZraCmxuMXYe9eH711SmLfBaRJSnwcQhAs1ppSuIMVxUaTzz3+2
n1tafP6ljjd4AraYCt8vlwT0i9z4BqwDABwFxJ+9mLZVgrWgq/UWyEPdg0AVrEmj
ycEmJYP+ibs0v18tICe1clvZcfXyHCOvuF1U2LEzvfYBVcgcW0Pw4GlzuoQmSNWp
TFgHP0bfoFjpMcQzq2m6gej5cEWOnR6vIhIeYrJSe6NwjI09IPJI7G6gJ/zD3t4C
7VwOWAT4LJr28JRAd8/DFV7JjOWPhuQCK8ruFIwwKIj/Kx2UkHIyeLqpUjGd6856
x8gnp2f+eorMUHemF+q9eQRfgWd/mECbrgX88Rf9YwszkDExBvphJaVr9vdr9M2t
Xj6n1NkEuo64SGWQrnhVW31Hi/9mwbk0xFWx+lFhaKKATl3O1sG1Cf8TM8bsLdFv
1bmqqDuGCKLSOUceopH822mV0duD/KLlIiUOEKt4yu75ZcvcMjPepNrhCodwA886
GHW920dldtWzIC8zgoovUGbqdcbg9L0YxA7J3BoxJF6K0ce/VXjF5E3iHD0els+B
Vv3AgIczH5LJIUfOfDKLRdohWmRWj4zrxNZBW3DQwZ0y7xxprav7MR9asPXz36QH
gBBFr6xsF61dIgfeZMyMq//yIx89XwCCchBDTgw5+gKbLscxd9MEgeIU8Zojw0av
3TvaD7w6AoGg/g3vmssaMji+xQsA2xopF1wFtd7/4MSX6+0kuAEvt/suPIjHX316
oWAympUKWyVnuHo6fTLuMKkS1Wzq7BM/SJ+Q2K1yZW9MTAhActgPENI0PXHdt3Kt
DWowqbP/FgOGnk9lHweOOXpNC2VjBm/kEQ0BFnDmLJvPb+4/aAQ6Mo3xeJqJLSSh
ev5oe4B/jEkmSFg4gdBXLaOA9jnyEGnY5YvUFDI/slfDh3MGN2w4TwhP2xfG1Arm
twQTwo6N9YKm/OIIq1FP0GPds1XUJpg0g8tj9bfBDde0Ql1srdI51fIKQd/mp3HO
6ZP7/i4aLlyj6TZG3DfGed32jTy0lWwQimpmLbQejMnlnxztHUuj4HXroWHvvL0Z
gBpPmjt5HkwJ8AzFZtgxsykV9rPDMvR/sqktYqwqPUTrIQ3dFwhphHH7xH2mY5uw
gK9sgzBgTKYUpxmWSWVjHH+i6tlStbngvJNHIddIBQgzDl32T0KVThB0hIsim48t
L5aCBTZdMW9b5PEQ7V7xER/ysGVdkkRS6Fx3T+dEgw+9ZJ0f65EqBQ8S0jk5AXih
MPTHBhMs3STg17RaPLtRYtwCqiv2OBeTWNNEZuCEE004ei7hkNHaYAKdiX3Q88U1
aCjguc+BugJmAnuzJcYAUBJG6Erc84zbKeabxzLv/wh0QOi69cRW0Xb4yGA6xX6n
5ua6mVsinQDlHa1z2mgIEcGuZ2dOECgD4dVzVniTgAMIntNNrlgbRECfombSJjqO
qF1KjyOOPe2i9T/MgztzlEkbo8sfAFo6K0MHj5u8RX+3N8S13zE1D/2lJk/BDxms
jgmytaFZiIDzMcTB4tEP8WQ5lDEeBHgCm/k6zhJYfx0Bv3wbXrQNbcjrrGTk+3DG
ltJI5jy2j5LzwnU7QiIQPksAR1q9wcWndxvz2EfGcLSY4UPWYK80iGbVSkyqMHEy
6JMnA4/bbWL5XIjVIRoh0f6ljVxDhsWLao2hq2Aq3lHRtLQgQ3/Ob3l94U+pwWl2
httAyGu3ZTt58F0cK3Va6S7CncdySZ8rPhTzonNZnRYPCY5A5Y9PIMbbp/V9ToC2
ASUuV+TOip8ZfTD9uw/QCNXUFaNTdbgSNUFV3H8EVAkLJGSkIg/G28O63K99RjIA
YOnh8YvGaqlt3lYskawTuQMaxoKDhihfYgo37NqbHdKqzDfRLadZWbvlN+3Qekd2
s2VnjMga5stESpNBeFN8eyEvzDcnAMrakMbnORluDzN4+wYxnp1vL0YriqIBK4JQ
vveZaye0f4YMezVzCZfxl87AkiCTt00iElZVrRkPfsnBF7LoN1WPWYL2BbXCSOq8
jk/owF4NcjwxoVlTVYkIIoTJxPL8m1kU7FLhQk/t1J3/fPDKv3GPE+CvCVxyANCD
U0kGx8vYkKg+/iGGkLxLXujFXbhxULrcs2ROyhukMLekeaH8WAePT0Ud0d+ttCIh
XPEIyhldvTOsmRf6zArTVfw3tIHUafKRIQXiq2fyTFga3C/dH6h0Q86YStGz67wE
0fP0ReRcE+h5/fqwnE6VLmyts/evIm8es6qHzbaZUZ+/uh3nesnH9Qw1WrcNX/Py
MbqIbJakCuFixDSoZUAYZ6uwQbNeOTyy8xV6/CyzeUptcvrFIi5U9yi0h6UU1nak
LfCjTcAEWcuKV32DEgpzYYk5qNcick3ASUQn+YXmjvb78E50I7SwBNP/j4vF2Ouz
0rlH0y/4OhcHWi/TPFZmnsljBIhtjCc9fkQWVoTMdsIm8JAZud/yGLSobBV1VnJb
sNP5n4bMoG521c3x1Zf6SKjfyDR6CV7YTbw24ov4lVYEQLqce/FkzZ+bnF922j86
Uxy6nw+VqOgpls9TG4yntv4VlutmlVglo/4lr6nsYt4xkFCfgxELILS7WgOs5E5m
nhph8+lG+UbuUJrT26eWQEBYUZusJdoSztnZc34idWFEBVFGat5tb3XK7BGd5hVp
Sc1RwtWQXS2VZSa6fwIJ5okVWaaUzzTObZbp1Xl9Nylb0+AL+hsxu4AODk4agmj4
PAYpJ3YnnsBDS2fN9frQdPpfgZxkQp4ebhlGVtK+gb+IQ4XubO+J77NXEZuZz62u
yt59rHoMAGF11tjwNRxFfpvMAwKWhUKDzPINp7MEwLvtjLzRTzpQ1mocN+MNKCGu
g+qHrh6LGpWC+iGMBPpW59sivi56/+1vapbicJW2Do/5wD42QWRk9AgHq0AqH4L9
/ert0VaQaI1PG92lo1FeRAzaAGVYJRSvIb+yXyor55A9H1vhKXMwQnGzubb7Gxfg
8pB1QtMwXQghcKj2tJY7Y5qTAtOqtfizfB/kIZQ5svIUvt66vj0Upc9y5Fzu+dxh
NJoQ8IZooQNB3nqONz3F6xSwQKwnzq23iVp9x2GMFLWTvIt4xpCHcgt4iCiMlDkv
Fv/0M+8Mou6UIBd/kxfebMvbLuGtLiA98M2v8aBYjE2O52zq7Qc3mNlme/4veh4e
sxfv2JLnldg3SaeNhvPRQmc/McIgxztKt+pcp84pkCloP8OC8t+v5T+/R/hoAia3
S0Xp7W0zXfxmcZROvS1BZVDqzsX2r6Z0/GleXpc5C7H3P4nj6fAeRHeygLjyyRgH
8PRjMQZ87t6b71iXjc5Xez+hpXfrIZgkIf8/8k8nOzhoHREczWc12sGLdS/lFVOr
MJjm8FLmTLPrIS3OmX0NWYNkJ3Q5WKMbvXELY3fYVIzUZM+XWhKsVZ/OFdhRETgU
90rSoNLU78pXw++KQ5brXTVYK4auq+O7ecHSlRdfmdXaWgRdVzmlBBUVM1kCenBV
+2ctfioPkhaPVr/5d5245GjNjEU5PHK0eNv6MLMflg5FlePBND3tgqmjahshNzrW
iwJ/RyEYH16aKAGbrjrsqoJZ3tFhlmN3xqEqWoEW8m52iXlq98SD/cBDwV+uJ0aF
zMm969FVuXiYmvMyRjGor4SyzUee/NyE89s+bRIrIANqLFCvUDeOsbrC8mPVw5fh
+pov9Z2iSsCvJfwfZjQjT9Xk9kV4t4koW/xiJLALT5lueKV6SUFlgrfqrdOf6MKw
K76FKYqS4uki51FtEWKdX2vBOXr6Z+LO2NWcZjlaE1RUQ57mvOzY6SGSA7rTbnBT
ofkGxGGLFq1WdWJ6RwKloT/etsdNGzWRYD4SjeflSbRJAFfZCcNWhCmAUYPfClP/
U2mgaCESsgzCdfYTeIrmscLLnYmkHTTiiYgNy8Dl1O7406yQlqc8ATmTOYlLue6x
ozD73g201WJy5eleeE6VoJtHhuARdh3/GdJy/H1qyPfuTdqnW4hfGfmfag0CfvQJ
FXRgcecIzHvsaWJjwaPk/Bo/E/ViHhuTNsrL8UcMcsiGj5H6s+tm9NHXd/aVchSK
KinTgWSic0Fq+GzucVcgGgpz6Cgtko+0jJSyyeyQeSvB9C3+RNSXElcNHhamN6y5
CCIuyQb5bV5LONT2O2uDZxMGMTTyIATXD0JNgRyFadfEts/D1J1P1boTUBYgrajw
VBXaN2eQjxuhZIuqu5asn9GXDMTT8To9Y9epX+GuTEoYuJ00CED59hEjjjqq2SrP
G37BiA6RfA8TdvkYWZhBt8w/FNJY65YyNfM5HwN6/DjRhoRRRATvcqSqv1b0ceAv
ArJxlcaAp8dMj6LODV4j7BiaOfo8MDVVwzb60+hQ44XS8twLKm4cu3jusCLutMF7
E+xnV+ENXeV4KwEYW7s2Ml1KMw3cjJqCdI3t3im277UvEcH+3PZTGF9EvwHs811l
l3YYqNrubE36aJtBXqNEHchQC2AayXPhzUlPgq/fBZ0tuZuCOa/rczUPELCO/Jzc
5odEzUpQjqxAgbqJu8xD8MziCGEO75RSxgKLRMhiMkjJ2pa2x/H00iwpHuyFCmfm
S5LwVaQaY4ad44CL6p8Vnt3grLTfQUV3Uy8ew/6663EluiVkOKpK6rmqTMQbC6Dt
o5Kq4TiQUjl38/+1kNgqWlHYTVgPu19brwbD8Fx5m5alfLxl5wi6go6k5/FeZypj
zbN25hKl6dxnHZfiKUqRos8gGc20vCyHZOwZBulGcmoO7AwI/WCaLsEK+DdXe9ZH
ARb1g2NpMkVmBDMUaBgOLzEHfOhh224Wv4MTyJUrTK7M8YTpm4XaDuCPQzIgfL33
UzjLGjbferXzBQh+l1vz29mFvnoJNvCWTOc7FIxxHRBRrb/182/jmcgP1bN4hFFz
wBlQTsyZCfzo/lEDkxRojckEKBZm3HzFXijIVB/sEFv2j20TYSj1vENhXnyodhz+
8nTXxW+omw/72j7Q0mTwprZvQSu/iAwQPF5KizKazMAjdBChSX4XF6kmQh4OoU4i
tQTi4L0YeblXkttvyzChBI8MnHjgZTv6Cr8EjmRQVJ5ohPNzcDXDcOhzvrFhJnwb
ycsJsRn3k11pK/zxy9uTuCnnxrVMR1xGBWQ40GS09SoDRBYEVTB7sJ0afTxseo87
qeAwRDIXOpWaYXCUotL61EC2u5xw/QAlPqUUC62RyIhUljUrA1rVnZdcPQ9cMKXm
U7HhK6Mfz2JkPd7dshZItEgd3QwRAZC/EG4JxYEj7G+L2f9BDcSYn6B2U/m8BdiC
6v1viYNpLk5HbnPxhT+bTub10bcbHW5nsA873x/99VC5MRgfyoyw7HfCmP2WRYpY
BgMFS6wl4szeK0KmjL/kL+pyU6aig20VxPsxAD+dAfcChHus7slty0RISgF+AAMG
BIbOaKyYjVGcBmyI8Z3OiozRI3UNmc0KfDSDHEpt1FZMaDgI0/d8yX4E3SzPhRWr
kKL42Fe2Iqc27Tq6Wq3a5frtfjuV7BJA04sLXtMnlOmTM2txx5EfPu3VmsZj+kBU
jU0o7LU4G+8wiHn+Cs7NFmy3yV3QgXhqBtQBOYunq7sc3eao8gk4htz2jWGdUqUJ
qMqaq04q3A96ADRII4aaRIga4Wwd2VuXg5ssmvp756Q73yKfFhRbmbzDRaySPuEo
QdlwllMjxrAtM09fLrV5opl5PsdVwYF+WFJkSs+yUqIp/0YIL+goXVHVdWZIPOyJ
Hv5uOdzTpwAbUEcAXQVCKonWlUGpxkVyaqQt6m/E/88zg4FQmQd7EJNIY4IIO7oi
DSne0f3B2j4trQbnlbrKIXFxIxUzCupk+nehCTuYWZjKEUMUIDvn4HSwZDo0gmOO
XUsDA2mpkAKoglwNjMVIhlYOFELY0fU5kjbNf3Yq2jpM0QYZmrossZvKH09PtVEl
G3C7xkdIsrgNi4L/eAROG+F9RuK+Impk5RjmFMwZmnacDHx3zBTzA2TwJIA8YZ7h
wWbAnFXL1UhN3gfCK/YRBwJP6Fj+Q/liBitoqvdc4yKhw3Us9tgw5cJ71IDT7640
6M7h7BvicDYPnAYV5LMJG9HJKBYp7yq1N+65Z4pgEqbAPiU8outNCI0sf4Su4xvq
fqoi3Qr8zMsT38bp8OuBUsU3hhyBhs48F3sFBOm54mz6P5Gnz2eqIHhPNmmCmhTQ
yczI4qUcmH3QtVMcSSiSrkdYMQ7SGoxqRctaK0rwgrOS7UN8Q7/6mJPxdbBDRM0I
k9qbyMmxt1AzJ3tkBgITt7zMnEW27HGe3iu+ixCmTIjxIhRR00f3D5SzlHIg5gZO
7f7qwM2o0KFTisW8l1hv+sfq2R/P2lr0qul5jbcMtpM1e3m/ryZZIUz5982seIQp
qscG2FSLgvRfjzOPnKlSrnAI35HBinw1YF1FljKqb6QNbp76EwSR9ZKAFPbNk8Ub
q4zWznpr76YYAC2mHHwjzMbIxx+7YBhK+Cos0MoaM2teRd7U9E03jE4prPukKCr/
yLCm+PdUY/ac3kg6c4UUa/3E0NDNdGjnZZvthdksbVOPZU//bSDMAdcfZkYGO5J4
m2bkmq+0CsxdOUbRaG/Vxdv78mXnkU0JOJxWbZYCXRftHbhg9sMVyCVS8BUotLQr
3RAyYUH6BtDh0E6GGpLc4XQx8siLqJTXE8KpXzFuVBH27Sum2DhGIspEeYEy4TOP
+3Tp1ofDjDsaJ9GfPKTgfJRW0d6NvSMLwuCOloQDxSU3RJ/uh8SD9S9ipoK+ZNfO
92/DAbSLTilNCEljjsaCPaEYGTEYUmD3Bw3WzsMCSjOihUbCeE7C53ezYVnJU/8F
6I5u1EDvsnsmBcsY4s74xlWii4n3ui4ztBrfz4sa+fR6/ayVH25f+Syrc/UznXhU
gMvkX7YLQpjA7JVG21rSBEosqfAWEv1uyNZSUHmIiDKhVXFvbukGC1J3jvqCT/sO
pJ0Me0Qwk+3Rm80i9XvSswjq8qibCqOL48KnARuijzs8dDIPTGY5KSCXMeGkx+ej
egm1FcdX8nTkGQHNWvV+6HKReIf90dX/bKIKietg4m470KOaWRgL8Ukcf4H0Burc
uEJsSkAaiKI2LTgbSyvEH9rJBKUvx90HiHXsBaOc5QnDxlN0zDxhItJpAE4QbyK8
rMX70c5BgsNtDglBrsC9DDIq1XWIIk3Ss7t/AHexw2990cA8svL7g3YkQJCO4d7I
T7MzjZKU9LOCRgGlbwVU3lhsTLTYUTAsaFlpp0/ZaiuGJ53mWeXXNJ/LpbrPY9s0
XSbgJ/5fNgS086+szxpXqe1Q8kx8O4qefG76zxMgwfiuzMCXDE7Va6CBi+FQLHz8
dSWQO2QiMl4VBsnoGLWYrOQBvQS+06GRKIN+0NfrTwR7jX+AMJB6VjD4P7pCQHOq
t1/RonbVZ8Atdi9rZEWLXYSwZD8yyiGvo5+ApxwaDhhF0JvAlAazk3+nhql2wDJQ
dQ2Cc7Azy/z7z4SPQ3/CTsc3MZc70bu4Cqh+M2RONPbjUiy8abZ2ZjJxXmbVI0ij
eAYNWgnJ4uARQeSvcku9OVRBLNweBc/WMKhM9cLhE6X78LPT0JuWhZDS+DD04+iZ
zm6CLwn/Qhcy8kiUgmlhRI58253V3kfnC6MQ8Virtykp/zihRkijmY8jzytuV8pl
H/iCfqgAX7p7FdUQi1s5pbxunIU2e/hBZOY9OTaN+HtwFFxJD9lf+D3V7P//D6tp
+j8gn0RxwEbmSkoRnow07ag3SRWqMWC/B3GAwm+FB967mdRJJv4LtDmYCK5eVWer
CsjBIBfqsq3UG1xNc2Y33iimAfdM19vuEiycpCdTXCXWo7aEfGqVeCZVIUMlRePq
FK7tD/j3317wKVbQu+aMvhkw3mHpEXvk8i3MNY5t7yn48LknFovI9ZiehftR275M
//7SzoRjLQcoKK2bWzh7ckUPVRLDDuQXgtsXWp4aLI7c9RroTxEflxauTdxOx7fp
Z32uhA7SIdaCgzdNQE7BURHMmOgZT2CUhl1wc2WEmiHpPvD38YzFc0WEfZ3CgpXq
4q4J3mcw3xX2sFvReDkw26fQPKE68VxacajzCGM58skn4+vv0DRmeV8uY8xd+A8C
DZ/nphiWNq0LPuZFBBopohC1FzPGobKTCxhLUgsxlN3SEsTY4MXfnNkVLkI2XRMI
ty7r66gU0YLPHbmuWPGkNiicah323/JW/QrrxO7yKZCocf1Wc88oHbLAtMDSLPuy
SP7zRUEWDIr3+LOHby2a5dy2yjBka88QLLMmd4YLrr68Xc86tikGuztkJJYMQ6qX
KwwoSyxaX3wx7S4CJjwilFYo5ESMLBExbgnhWbOpM5oUAQdtnU5vPwTkDF4d7+g7
Mbskjhf0QpVt5h8FRN/QeYtVHUNut97gOO4F3RRS/LLks6tQH1SpYE4uvdussElX
TB24/mPESGj/v47Ksw+Rz5c/fKd+Yun43QxAns1lPHSgYmpOL4vn9/CMF62RhAb7
hNhBY1xTeOstXJHqyqFNm/UYzdNCCdbPLzcVZ4xw9Cv15MF4xpDAR4fmazvGn/f1
Xa9Q6mL1EncDCP3FkhZkCFTEGOsFoNNJTbNmcAHm7w4PdKh00NuWggoSdx7gDsoE
1CH75Cpfr6NkhF3HTGnI1yQeGW82rDYe9de9uauKrWyKn+wVMEjhwnvSv5Lh9C2e
JZg6SgKLAyG5vu68wPfAWYHlrLaCsbWTKkfxm4DICslDeu38YwU8mmmvNHLC91X8
ALMtXT2JaneZ3jjfHq9IZ54roh+pt6jFFL5LMi450bHHrIAQn66MkCYfPw3AjCoc
JIRn7M5mHPeUWor/J/a+GUCx/rvF/jxQjv3IjMGs/yCge1D0MfhgSpMBdzFzY7Pv
vl60PrywKkXnov2zu548C/dOhet3b5p+syQHF7yJK7rSHLuSHkSxJ+vuxXlZWCrL
tu3WgHzQnDjXdJ9U0LAwfKLQjdcF02Fc2KuniwNPe/G+kgJME5BdgDMhqyLzSxaT
dMxcK50Zhq1CSq9J9DSCKHrpAqLK/bsWHYXd5tEkFVcQY18Zpxuuvk+07j494VEw
b5RwMa7ui/7vwKJ4JB9Tslte9gPVu2PTeqDAVh1HpEe2eoNuVRXFvS9tj4vO30bi
ojVBdK1em6sKeFh15quyTAmMRqIWeP3K8gGRGK14Z0X/dYbR17pYkIbl1tgPexmV
JC1CIPLQ5yj1MSrApTjAZ/Pi+LeUK4plKP9jZGGoHtKMnR5SyxIvcM7s0HzcDHw1
5TU26USDEmlWLamJVQ2OqIlGxGFrOF/SRGlWQ4al/uSVFdjG6wTv8FNrviJAOInq
8MJz3H4itY/bJuKljzstRxSNdQaTTFs32H5skSqlDVpuiv/a5bD7O/i9WKoN/vRF
lfyeU+kigEzU/kxbEIy06ZzVgoaG2QIZmHZeXhcolsQv6i+6ItNnygXieIY4+HGI
OdgkmZ6wwbCrnL+6tuzMN+9UOTfVX2424LpA3KSDypOKW8naNI/h9X9y9nDI6SQM
TTQLVN5R+Fi6SOupfvmz3GuSqSHJ4gfiUhyznJb5nrC4Q0xoyHWr/iHGVb3m3i3N
a3nf4kzGTZEyUeEQW125mZ1Z4O7kmjHKnhd9WhL4IeF5QbHBVAa9MccjKBjohrnV
iLESNvFI5QKJ5tfa+LnvoH7S7NnQZzBZ5hicLQ63QceM5ysNhC32q2UnWLMPKUIL
SisnRTiqYLXyVjICAULOt16Nfl6ajFZdXfEqdiGJwg7yZWzKI2mOiwYxDf1sfjhB
bzZj2ShoMgINa6N4LclL9ChG7lRq8o3MYBWfHO8QgGettC95Yq0qmBKBq+mqdjos
qetEwqILb78oQHyivpD4UkC8YNxFoa1YTO2NNwWoO5NvCICuDWL/fkAYKqZ/VjWN
lFYiBwTZ2MqOyRdvBHfNmyY+hu8JMQV+O09DB4yahR4KM1BefDeE4n8Qfukg108n
TH5VQ+SQ5zNnNgVgFkr4ZEnGSmYL1+iW9+RqHGZg+Ii7FGM+AawJk5ixE96ooko2
yJb1rAegKA32GkPIRHjGmedudmruGngMZ38UIsbFW/oizvAq12oDHBZs9Rt0MUie
BMCUCl5Y+QBFM3fO8OA2PT430qL07dM4rgpnZp0NBzxfsCnqSlGUTPN9max1SmeP
SKcDSd3hLEm0a+apozFHzxGW9UEMrCU1VGrX98/YUlBpw5Kz6MJwsrzqFqZtFUSv
WdhHvNa0cZJBjWauYSELqZBizGiOvZaqSIB4vSwnAO3try+NOr5MQLhSj9DRR3Kz
tVHT1bASR5kvn1KQodYvdtELVtmjXqBVFlo/jd6hyTSt4em24oqEL16/T56BmP2S
K1QCGllYw5lk3lhZyJ9g/NOasD3JMu4ODUOhjrKhO32qqwy95GZggpUucXyWNbmg
A43snk86I3WvG6RmmyInkNY8xFDfupo7D8VW5OU0SdkEPmreBqMvjD74jWiYsY3m
e0IPPREK7NLR6+wHMtoEmN1SEJqMlG4cb7Khg4GZODWhO2nJrJ7tRpQnu+Shqb/Y
iYNI2SmLOpBbtlABrzEdCsnWtVDoEBmcpH36bHJ4Ey5aX3zO/F+Hq+DhYkQTw20E
z94GVdfh1RMxVKQdtFEmsHSDUmTMWZLmm5ywQB+/b6f+ex1oyeHSsxIwfAp8ULyZ
D9iXVriZjdRRnETV9AjhZYUb6HJge2dXfrhtKtbNNl2UT+aAe+OdlFMx1U+5JCaI
MFjLTDgcLcuXw86Zhuc57fAqaIt1HHve5VtwEpU043ahwDmUMzGkmhzNviKEJs4m
3OdbxpQb27ki0XJpG2KW9c5NzkrOksxb8Cwdxuw5ul1H4vaX04kmcpbafWEAlzry
P9eokPtExS1MQVoH0mXHSw9QWlxXG3OQe3YvaLkNQsWb62UwuqaFXhWhDrclxJTz
u8XMK7+bSJTiaFT3B0NcHrpfei4ScYsnRYSX1IOWdwO0ExHQJTyBYIvrzZLVuhNe
cQ82qx3Jn6Kj9YUi0OaKw4cDdBLicsZrQkp3B0ZQuQrVoIQg3g6BwAVY99eRlwQa
TiWhcLAB696TSPV1Bfja64KWD0YFXd+3gEcO7vMgqljjlaapwqicJf91zF3qf28I
MTdPdMONyf52OM06kyTJmgIlM+9EjPBUzszr3dMTPNS/HCGD10KGXKFPm5hZloaJ
6/bjGSQZ6ZPnJQAaPXhwC0FmEsrjyUIv0myuj4Q0Nv9gT6/99UjGBytlDDIKrQp0
IF+09fnhM5mXNOo6gYHzvx3Mq21NWd7818o2TSf7v1/NSQaSm8cg/0Yt/z4HzJFn
qly0aAkDloyiNxkvlldswHJFYVQdfyOF/h1xMEp8aZHWNokqt+0lqik0XPnfFIzi
3nYXCTbop36xpquS5Lew7qLg1i92uUkyEDfqYStwkvS7iPF1DDKzauSMWtt33m3c
LEtWmg09wavb5PW+eZD6bNWa0cGYBmBh/z4459ToNlO90XlBL45h/2brHThbR+t6
efB6CWj1dxcT1gDden6DmzAvYkZa0xVuVNV+AZKMQLBdrpwxYa1MvvuUs1/uvuHi
fDdHB3lDRqSJBcI4gozPLNUPjPjIcVXRhoLsd4srKCAU732RcC2eDGkCOCUQ/Qzb
o0dcBz8ocVB84YPV6Jdko5YiyaTyl/g0VMAO1KKw1asCl28J8KpeCzPb5XThHhjv
t5Hr9xJL3JvGVSV8VIl2/MTXDkyNcsVfgqZOQgHqN/s2N7q0Eq66D2qXBg7LY5c1
JnWDPF8+JS0RLjZ7ecUAle0wVpFRnQakI/7VFMPfk9b2k+d5MQASB4cdVCJzq2+h
CTvfu/+vprEJ94LodIBJlwGBZ7+/zqoIow7BV+kNvUGUnumLKBsexwyo4hH19X2a
u7Y8oCygaUT6DAybU/vdoAg/9l5uYN5M7As3ajk2qa7cLn/0YNTQCuxxkD6/dXre
BgphuRYJwCsq5bQug61ODVD+sHUEFvWvPnpUx09QrgJJk5elLUqtKnr9OtRPNGba
9vLJj/C8pzfQlgWz4WlnzwWkl13QykQeMRJ42KfbUcyK08rfmxYVqiWnf5x5fKkl
T6V7Ji3DlHWpbahLc3KdIf3T+1tM7zXsU/RIvAK5QQUTP4vdaRm3VsBY0chRE2iK
QI83wwncJIEUi9u5ocEh6axM+fu2U0Z1+BxGOfzYL83oZfi7sQ7dpXPe2OV1YVMC
mg/yBdV/7D2YoyD3Ows1/byzT502obhussN5Nimio6smvi9mom+2ZaO08K06gMmi
pUYjILhWjrecxUaf2U7HEByrQwkrZb3SUYoeWrqvl0IcR6CSS9exfGLv+MnboX4s
g9pnuFi1oCcEbOQLxEKyd6q80Nzw1KLTtxnhvf50q83RI98gEmhOKkXbg0Pq46+h
MnEa31ssB94T6In+8Im3Z89ILVctebsbObKsWZRbbOWpm0O8yZtEK1DqsU267F0M
1tWjFDWQxrzZU78+9bpic6Hy1yjvjJPwFSafvlQX22dFBbzJ3NB0/HU5NS6YeFRI
//ChCXpJRkKdoJkIRB0VxOPhqhoX1aaIN6AN/XHFPGks207XozS1x6SqpXcROJ1o
IV8OnBRklEcViONONNulnOWpp559ZgTTA3XsnF5FJfeGXHI3oi6kyIjW/stDiF+7
IDpUSRfIsolnUrkAaaBodkzgVV7PpVHrQOk/BSGhgKJjaTcH4YJgaxrKQWzyKMJj
M53KPxSpUddFYrPPSjXEO7JMbZukbQWBBZPXOAJMFcIctZEijeFY3U1AI6pqdDv5
OlBb4mA93Cl7TFsGfVIi1Pilq646I3FAbzEX8S/dN6QGA+DAA7TfjNQwXGy+lDhr
dvyuWR1Rh2flxSLjFZywhUGMpG8BXoI+vQh5+Tq0JKkJAwu9NPcFCUp+3mW5cxRo
GdoRI7GtTozkxoNcNf8GWhLB0Cd5CBwPPkPZPVwVV2Qy53vl9OfAkqoB+amFlbzV
itEHAhmoJlwcxWgKCnSJPYVsZjV+YMvfdtNJ4Ll9HokdIHtv9G1tsklwWxnO9wNG
TO72KxOeUGE/fvDgvBVi0q+OrBiJzf2Cnz+yNSH1Lv6wECnqSuvP0qmUmzLq+yDD
IH14+NYi/T6cTtzvr3o4cJPnRSa80esR188UP5OnnTyGrTMoR0Wht7FmcMdKQf+/
brvTvfyQrU9irEYfL8stpeOvHjJ5X+UbtLVAZqfB4oL9XtVlgYjHG+HzQFiTwrrS
YSebrs+5x5OFx/2rNXPhJ+4yFJGIZFftyIaGKkzKlaevvhVfiQpFGCAjWjACKl0y
eVokNT7sxHeKYjIIHriHRmZHsLWnKSEiK88Dsln5eUKHp2h3Gj949M0jXLqucgXV
9grxu4pMgpAYs2O+2ZsmrwLc10IRKltHiKOmFvB9vRr08E5L3YVBBf+QdFzWF8CA
ueHxe7fQdXDRlWwIrouqQ405jsXQp/NJ1vtiYGKgXduP0k/MKcrVrOmzvVvc6W7V
6L6r6NeSyW4hAZufQxXAW+8kqpXs9D+FnLstan45d5/6NsiIXYHZDVb2rNEqnWAa
3BlCX4kXi9IHhjq3fotWqvIWNd/jDCKYOjNA5ibAoPxY6T6W1z5D5dVM3wCaiqKy
CvYEb5SrpdAtpKqVxFtLGz7syIl0OXiBRXIwny2FQUNAx/cwVgy/zDb2q3jzIrtg
W/o46Cf6Q/i1A2pUSf/Gm2y15mABY3kn9n9GtWMzcvUq7fo+oIhs2q62MoLdZYV6
wylmr5ABXxWG0d+5p1O/kurbmUg0osG0Euloja5Yru4XZnKUmtuK3K5a06vq+m3F
5f4/VpVbGnxfVgFwZz2H/DcjyMvQ8DLsI0vjLQVn0gOk6VkRIckidZVAyWEm0SM7
MguAN4MMLmOLU0cYCnr7T+63o5ryBHnTqoXIRQw91SRidKt5Z/cKtANhD3i7yVBR
4Zaq6vxEoIFw8lzcVdAbtpmBzHuXCG6zqqtSD7Hf0a31toUn1MAKWqJSfV1fdvuO
s97OWdh9zrtaK9Cd1nw+b6WjRg1oq7k/Mgikej6OpPIqiiGj3GgdJ97YxbzimX5S
0EbjGAaruls7uXUarpNpNC+PZE5E67nLVXSXhqIIjPVL+9mIjUWXemAL8Jqr7D3x
LQRb75ArGV/bDcoGeJYeeC8CwIYSghLTt6y35O95/3fxAP49n4F7+/5XGkpuF94a
Y2lZVvw2WlSVDDLh3Z1/qXWsoJRMg+U3zlxopNg2xZ5pJuG9PLysJRYbo1eB3hvl
qfKWUYYODarTy33pWp/YLIi3Hz1jspnHX8HHR07KywLo0g0Yizdlby8COcZUSLRt
fq+MJWDRk3eVFakxXGtK4A8HiXEK06Pz1xpYpo12LmA+CR78hiS1RCpQxMe72DqV
mL/JukhVdRPT+eykUNiES8+okq81iL4r6eQn8ImBAf/ZOcXJngsjYvMWT45Q/zbJ
Q4mpYzp90TwB9v+YGPEzTmcdhh+LpOBwJu1jvz2t3BNrO/aj5oZ+JVyjUpIL2YuU
0Q9lKEhsWUSAqoi3KfRAGtT3hQbgZ07BRpjjji2A2Ih1eRDq+pDtkOPR+D7BNtIw
hyzXgmyo3WaKPQ2btC7n6JBfJbG+pSO1yBOPuSwTGlqJ46VwWfIqiRB0xEVPNjqG
Ifv3lEpXp8vXxodjzf23kIG7ZcOCVQ4vxR1KBmF8IJgXeprxzbvb4a+yc6qI54Rv
o4v6gul+1nK4t+nZ3NAZOkHF+8tkgBKMV3viyHAKBS9fxUaAjxOjZB7EBLgPj1eL
U8KcmR1kfmnhdimvTUvMWr53XvLno0iMKoCwrEWKEPnd7NQ0eCxYlG+jyLRfYruR
e61/uN4KsAJQ772UUE7Ic6WAZm9lRwYcG3Eiu/5CArF5USPnOlwhbdOb+xIFUYi2
7zzP9SBy0riZuk7JmR8PiHcFjj3pEm982XGyzRTIbwL3bw/+9bJLTMezTRfU8ukP
0/VVd/t/1yZ79x8HGGGJAOJw9tn7qlB1icFSQzV68HeF2wFSYrnkpAwgJlV1ZVeM
Oze6YH1JBUbSssmviLP0tbCEYqZY7E612wY13fSr4lpUpMzkM+UA0Z2BK4+CYUIN
PAyFFU6UaL8dTKTPuTSiFueEr3QCimV40nrYJvtkKPyxq0tagLYiYbmOdoLxhs1T
VvIlwQGigv9yFCz7gaR4JVe9++4VR0HK5diutUNt4LM87BKpoOi05/vGEoMPxgwN
i+aqStJkk6k8RrCWEP+pbtACqAHBkLp4QfFSHzkqkc0yt+J9w477K7UldxEAGRUC
YAN66BCrb8VISNW8xjnp8xv7bc4Q7r8NNBCjJukMBwIx7nKeXd6cbvVXNJ0pCziw
FS50x70H736j3p+gWSuqKLaH2RtaqkvRKnIo+Qi4lf/oZ+hWMD5Ikvsf92T3fglh
MmwpJG0RGouVp9Isy6kNP5QOJLfwT3x2ojxAGjmQFBuEPagnurAs/62MXcd74Qmt
7TuD6BbnpeToTEmlaesBpP3YM1kVrFxY+X22EPkC0NgnAQfcHkYdC/jqt/CBPdFY
eEYuFYu+SOrCX22TmOLRkDPate0oSD136Ta13kmZjev03b1R0KVFaPpnPn2dkfWU
B+/KZt51Pl6go1oqpFLKBvEU90SZo84ZAhLFz9MAvTW6kJobYdoWkZQ0RkNIjb61
bBQrlCeynxITR1Rlxd0UGo3u1Cr3AOan3Ms9bcqyyh58AxEa0f1GhIia3zVsPw8Y
2xrlZJDSA/1f3chkE099GKcPQ/mQdH75TeFkz85KpojdnQUxrNSK6xVxCJ/51Ti/
41LRiEDkuA9ZskwhOgvkUVARXsyaVZZ7ZeHC/E7PIM2kyabLBiSuqiTcbYFEE3Wi
CQygOV+5YW4gZ44u7XzEQkJeYwuWhzKBQCXjGy64m8MDc3yCpp2LCMOsynydhntQ
BHHI+YYv2iLOo1ZGrmOqD5qXTlQiESRyeasOAPg7/AF5iLULZuyA9rO5IsJ/NMrB
0Z1m3FhasN7vKvzImEjGkv6Aeo0T2t2OA55dxYVPEcEDFZe3pf/hut5n5GDL/2lT
NelPK5pDFC7ZfZbbt80wxZzAHrXuVKdA1KH6EL+LBN6XiIs2pjrhS4BNWLb7BIvr
EISOawpuEJ/WsAh4qzPFsqvJZpilUArza4CucE2w/eC6CJcwqxE0o5rI84DSVFpB
R77MarjLXLCG8xNrgjVToI9RuijEY4F7iiMAHNfZGfmaGrmx+nSH2Qkz9t9EBax8
vsHrT97WWm0aS/cWn8ty+V1gPv3XS9irW/rIvUf2yBAH9YCBLZzL1NBMWjzSrqUH
eLTdJPwho36z8QZuLFOCuy57EWKEqf6soxSVbGy7j30Tp/jY5iZlWetfl17nh8uF
bnVcZd3C0pJl+8OJ7I1S5rzY9siuAH9XJp8CqZiqQGp91BumR/xTVW2EYm7NvOnX
quqPy1tsPxBHZxRKMZy5YsuJuIGZkK+EMNSw1C9uk4kGChTvoIEit7l9V3BbtMkC
w6OcswOl/+/W1Qwi2j+uhIUFH9Fzq4HLYg0hrlN4WVWrAWdrNxq7y1xF+nMGovjs
VSuJaw9P59H8VZSAYZuBq7I0ecHEagcI6vypHphRq93k4q+DC5E57058QSb61AMg
CZ86w5pHZbR20gUtGm/H82GJrFYIUVb+FzXB7eSnW0rooMVq6dv+MnIj+RsbUPBh
xwtxwed6T7DtjSKi7RCrEfuLdaDYTrC5JtSZmQc3Wze/91A5xQw691F00fQeJGix
rNk6W/mnd0d8BUVc4ZBd6Jgcz7ANa3XVs8Bb18FEpqvrqMb+Mfaa0muoqj7mg+H0
VOZ1XLHlb0qFpN0fT4uQRId2x5hSGGNEsUw8IQtaIQuUDzEKtiP9qaBFIs/ui2eh
VQRROHKd+/cZfWP4k6vkudZVZUDdFBDQGVE7IlonqWJrEh9HteiBq65b7rIzMAop
zeqCEp6l+DiT7u4esvT2aHuBBAjDuxguamPHrWqSfcvT8+9H+f4lJDt/OjBEhcpj
JadQH1sSZYDnU4wJv1qmJje78+9Nc3NWAXxk7egey4bsjmll5aW9OwEoN+yQpqWL
TmnjIUF4Xp6uRmZHCSUxxUg3BKliZDB7fpd5PQurMjx6QH501VaYIr5Eg8MY9DLM
Yyj9XmWxbQvGXoL0sTY3yobhjdXeV8Nwap87CLH5QzrAvvBaULICGcax1rIP3Zcw
2mhwbZIso56FiDyVEBZYthLKrbKC4o2t0wu15QCVwzTnDd03eFkcYUlenfZy4e4W
ujW0mZR6nxzvAze3So7A9wMXxDFuHHQJms4aEK14IqXl79kpAy8ChveDy78SdkPn
Ch1qzUziZRsxcwuZzNq0j+9bM39fKK3zntnTmAfOb6CS7z9k4xtSrQ47BkkC+Die
RdrrXwiTRw3MD+3+itvdvfhoLMf7JBnV2ft7QCxXFIvfTYNjLBL60K6OpxvI1+g+
+8VX1M4V5Cd2QH4lreCg5wCOwAuI3PUDxC0+yLvgtDSXDIZKmuqnuuW7BCdA03O/
76LAgSXpktaMwFGI5t/uJ+kNWBbTYAdSmGV0sWda0Rww+LpIUPMSr4qc6xootIgZ
qNbXgmwqDxo6oxgb21Cv8CFLtXs39TEhMiY3pdHsHulvoKmLgizlmGHJDVQQVK+1
7JHjeZWvse3J2gok7Am+UnhfD+Wo3PWA3GTsSLkPpjBOGkx7RC0R8oWn1qwlY+iw
2II0wFbUse0Vt3BNQIHVdUFzYwdxPdOaQHL7kkhEV8lJ61SvilXsahKOnkD+WRPK
y6wOYptzCzsnbEs8joJYl9wFuHJWJEKnF+tLV572O2hKKSRQFE/dnnz9Wcwb+FFm
ZudEnqlICS9htAUvI3OqiV1XWC7HI0ugk47inoJlyXxk3UHqM/xskLQP72IuOQH+
PsgGTNxflQWQzDV2RsUt61C3/BCHuuS7fMcb9MVMuabC3C6mmjUA3wjpsefpPK/D
YwNzJwFlzMGxft/bkMkHyn9aEL1dgGFbiZy8jRF18D9UxweifxHlQERG3M3CguWN
BQgNta7xWSKGroQFp/wrW5oojM8zBv5WXuUVwJEMP6Y2848i5I+W6vCPRrJs9kuF
Ct2DhRRvqjuk9gBuQ4ZXMWIigMRsONqwtMSIzChCLE2qsdrnVagA4o72CMVEjF2J
8y6kX4ZI4TJ9IwEmkpdOVIV7LN2AQLtjQxqWmH7JMNndOJq7gr3Kt2r5KyNBFddc
OTkZ9wB0RgsLsMBK4dbMw72C82BFachj6l/Rjwi5uJ91K6VC0Gjms/LtQ8VFjEcF
iR3e3fxll6JCzcnLWAUgU1IOF8s3l8t2MMApCBwkyve+7EFAvwNuq3T4rBBt2ZPT
4hFk4nTds8jIWxVfAKKOEkRtqEcosPLWrGmpvSog2zPd4RMjkXHmcfxtgY7yDBsa
lofwKo0QFomD3izezFlY+bScgmP20I+AN9XVugB4+FzJu5IRK7dA0Fd+DiW+/Gkq
H7yhMGC8iFMZcovfBOwGDLZo24ken2CQxzq49vQlScbm2s3Hry67/F6D/C1JSsXh
vETLKfLu0g4g4mRFY/3xXc0FB1BVH9JzYwoi43Kx0NwPkty8zdtNZVH4c+5U5hgo
jQaPxrQ5xjA6O+X78pm+0+zU2ydtDy+DEVi+H/3/xDPTBWU5bupljor7VwOb5/Hi
F9coGAxHnW86qmc+Kl9xvsnjbJQ+IaLbg9XJ5OXLTdJFQ4GaTwbZ6WO4MUdBdjID
y9pvDV1QQVW7GU27xdjxjEMxe+6/zzNX0jBWuAQFPOjULOw89abJ0hD1Y3KFhrVq
am7+l8BY1aKJd+XUEJfFW/hoCCq3d2Z7z3itDzV9F3AlngYh3vCDvYhPbBgabAY4
4Zk7EQtgg9dDzfQQYZ9ASTPtIqzz7rEtPisqI12ERoBz0FGed6odR4r7qN+9a7vG
g+z9SnjJNiZck4h0vXx9CtC0NmTuMh6/24YFuCuhqjTIKP67PW4QQ0D7PTINsGcs
pJ7RBhI0eigPUo3M/zc8yX16O/ktSQX1hy5Gg3Sh5tpXdhRjhT0XlP4fqVee3iSc
gKlDppbxmytTfKndbX6L82+3mLn/mHx3d31d3g0mkVjVpuWA5ZRVe9sxpxqSj6PK
olEBNYbq4AAv8cnoe4gR+p0qClfrR8zRT8qaC7COBp0qY3AIJz10+jdT0Xk5ecI0
JXVAlqkdVhAvsJTaNDVgKnPG1yPFNxYAge46bdqG4wWxm28v8FM3r3mdNVbafyI0
hUTb0AeZbyMTIVXYecg4l2qklwwVcH7rUKrvm4GKbK8nCx1/yhWY0eCkXBuxZ9uL
4UaBYn0Kr2pk36iZF0H0Iq5ig89E8AO83BZolT5rzCNciVU5lpcL9yEXch/c+CwV
wrxw+OEGpHooFSzn/066bWA7C1x1oPbwPGxJGuehouXJcNzWyHSyol7MdnA+e1gb
jZzhXksmSoIAMvExchFmnGAMTmQXlinZ77GUFNoZyBNWk6wkQwwwbpSDZIfTcaK9
d4EhVRaSssi3MU5k9wsUkzLLsaXmyveMfbbGuCjDwnqgE1Eg6f9zojyXjPgHDdvr
hnaPv2W7mfhYBzdalKBGlMMyt+NvhozRbvctpyuDOmCDGHEfIc7N+pc0h1YK9Kff
/NfS8MOV5u7wJUMbScW8ca+mBBQp5KIOzOdwbfDfqcEiI4PKbEfngVBFn4ysSCST
/hzC34s9e3ua8yempJ3cY7F1I+ytS0fhRq8o9vJKeT8ZLqw3a1B8aUsqfXmBb+L9
Y17o1qE5wgee+gh5DLfd41RUO+pEBZvb3+eLWCwmFCEXpJMnXfdjy+21i2tSFd8Y
UKAtewmmxDTGSBfUBxvzh0EozIjPXCKe+Pmk2EkiQc3keHyIUvKo8XjKHNfuVC2m
cIEKNT9+JpcDY//3FyqrdQyUgflUpN8LnT1joYXBBaeEM3MiPBsb9OsuXSGWnbFz
SSxSghPtVJXMfgX4H10JKq+nwr9BluwkaWy9hhm+WIpW93O5UiU4NmXOV3RjFugw
f6ethI+/xkWXTUkJrPR1bE9GmAFxf83ATR63sjZH1JuSB8100ehkrU5h3csG8V/o
3vWd3dYZxesdp/K918xY7WJVVq98/H8MWWTl9zZHMNMQeU5BG5DUECOEDCQqs9hI
rnnmgz//19UqqrMO/++IXGoecfsHwuhTkLhPf6AG5Ol7e3wlz05KPK8XFJEJ+3vV
2FyxOQI7k22+Ct7leQNjrNMQB572KtI/gE5MG0d7+fba8zn44k8kkpvEDSBfhzbt
7m/hU6+KLMKnPEMQ3cSg5YQsddTATVe9ZO1LiRIA5Z9F56DaENFHV0nKVmjebl72
cANg+phjhA+hobDZWRlFdq6IvF40Hrx5NzTBz+19DoiUweA5kqPSfuLQYRzJBOPa
51wp0ZzmhylD1qiWSJNp4XcuX9ceAeAxfJLoe1vJ4d4fI/ZwvOEeG9vGaFVXHybf
baecA/CPOzdkFVhTLcNHY6/YPpRBou6XRYr5Kj28vV6XY1X53HvhX84W3C6EZ8Zf
YFAGfbDJZDW82I+jRp5gBGzekh0gKsT/uEXC2WaDWJ7zbeiEPZDtL9S+f+8nRypG
CIi7cPdeUXcCMiEwpa5mBx/ORkcEv42irrKv1JqTb9kyNZoqHsMMxJsFsc50Z7Ir
vzVChGA9urkD/lkVDpHY4HGNkECEIhdJ+HltWceIPE/+gv27p01+1RxvH39/4Xnx
U2MBdeV8ee70TnuWvmXCp/a0HvgHbz8mou/KGHuCpax6efteg5n3R0rjBYhsbkYN
P3MbfgdXdMEDRoA8SgaJOoU/qw+Q7T5Kd7EHtCP09PoMhzFDuF37BOYKEiW0MJ8g
lJndMuWRtcbXSZvj+asA0Owoi40H1ja1W6dOp6ZpDeqhK7PL4nTu0wf25C5i71Lo
NYsbxxJ012fhAUcuLjbmYsi6TdD7LxZeo2WEXFo1+cKkF1Hrm1SHXIi9zdShYeTe
jSQDED+3phrXhWaX3x1RUgetjh5GbmLpbFQnCjHRRC/Pjv3sFvTBJ7JXt7NlUwtP
W2NgxZ3qpcOTHK/dcMbDI+LMaj+Mjdx70rUfHmjP/ISJ9WdX0iwsS7a8Q4iE4m8R
JmdSEJnGiEEdO5LGp4Nf7m04bN1yNu6K98VKr0ZE9p3RaIlMnL8iHv0JxwybNuRu
hPflIlaFTee3oRi45CWhTCzoQxwV6unmilE+M7ybABvmW0SuiX1YswNrYwQ/r690
UlLgCXFdpX5nxuDDz4ppL4BA9G6DkK4xsQfVQYpapDNe55R2hQxMbMcykulNTTz/
h5rhbnSwX45lMiJxNIdnV3cVZqYlmpXR/4uJDuWFRlgRNEZiw945apQ7l53VhFZj
FNhlHa+FkTFlyKCV53SJCNKPZZlQA+wu6JL15iLgDvI3WFE3TdWFkhNZR3ZbvxHc
wl+WY2OrTwhI4kBAw/7Al0gCKXtRACSS5zFDFP5QunJWYWrzdjM87TXIghcle2XV
vhjMXJo+MGKbQw2glwQOza1c8Y57Vzq70GZnpXtzX4QUWTsmS6HnsE0vLQBrbavE
dZM623s/QbYwTO5ZnOizR8cIh49hfF5Ihxk35FqD6P4F4fYKc9ePs+qLeuPkMqPu
39SOxASKtXeCuXkYH0piFw7+WFuwxRtmhqiysRRsP8Slwewm2l+8q5k1EpxhQ8iP
4T/WROHcv8BrK2XB74GqmrYbhtMlI78LvtIiSMUuozjsNUS0wRKN65B8GBqem2c1
X/R07kn08+OBVA/WlsVENAXYoyP5HJDa6nekrch14/WdmqzAb4kK3o+PYolDN9Wr
a+jKmaOG92xcvvhrEDa/sz+c4KDq/X5FcViqVsCOgHHjvGIspA3WiHImx8riC6MR
a2udZ0l7cRXnVzqmZVqgRIg8Lp1kkIfWcmi1+lW0EXp5c1EqDGysx4zQbl9NdlHz
tcTsi9oh5386aD2yvM3rPulbqY94jVbSFTewime+taF3SoTK0wNOjw2b8Cqcp+q1
I6SDY+JpCV7WjDvFCcoeXfg2AuYpv13F3jaBMkPs9lVydrauIeXXFFVFTb/oaxn/
/TFmAL19l0Zqd6urQTECddkiJ4mJy/ZpB9ale4cvxVrXPNgbLv+yd36cSfkJVSWg
xy+IBzBTv+9WKtzzKrjzi7mETLWdRnVTua3Hix7K1hWhwIhfYj5L++GRIYFxQv+I
2hC/f1iwNFagB1iDQWkO93K5yvLiym5FufewB7NomiTN2RcVKxxKUBBvzV4+C0d5
jXT/1/v3bLYJQwUkOtedDO3l8aJ482n7eLN+i7M9YItPDqhm9jneMkLQSsEiwMpS
YTnyGclbPIGn/PYZ1kTyoa1ILmOYqrSSbGboaeUVfra6wDreHPNiYyae0yVK+lag
wl9F3Ft/Qv51gbIuZKAzsV5VgY+/xzKv8V58sTP/1TGLi+SSoIJ+akclHuJRoi2B
ttD9vVaRTvY+E6hKmP0QKujXD/cJR0FUGlPXTgQvHkjumv1D29rfSBpt1hC2FVfG
FXh0e2Xa8oQQCzQdYwM6ZcI2y11byLI6gvliFemRqZ6pvK58BfHkoai+ywLUu8JG
XFd8b8Quc80HnmIrIJkRF9wOPxpH9F0Q80EpLD+kngNLbas8b1dS0yeItvrj/Geg
XAwCVxFtQV3jSjz78rGKTP2pI9moDWFG8RS1BHOeTvbFDfWYxxdN16IOoAszaZV/
/4stNMksKwVy17Kewx26UBJMSGF2rIMuTsDtQyu/HKHhvdMrqVU6sqHsrUvRWM7z
SMJ+AgPK54YFv2D9CJsO8ZtfG3HPSJpYzbWBO7lSX8/IW43u33mTcZLDOEHV2tNh
YhmO95qPrNuhN40MsS4opcG6qMCxXyf71hpmMS930y1IdD8HGlqJm1PTW99agABn
Wfoma5cVkeuh2pDFtlXMUoDDcjO2OxaI2T61pe6KlOvWYDkJwh2eDhu9DIGRAl7Q
yjlsiYCA70GwdfLXs71HQEX8Fa2i76kEOyBoKL32BOepiu7nWdvf8SeUS+XOXgiS
ZNNEgjpkgDo7LChuhiHuaodjNaBh6pXlaG0uo+pWaphKCwkKzTOCcwSeo4EeY/TQ
qCzJp0jN+VYf4FqFmzkzPoc27amUqOLfBOmignWdNmtfiqt6DNggskDgaTt5H2Kx
1TLUFDAtE8KQ1btaK1vvQV7a8kHgPHyDKtiJIjRkdH66RVg4vX5E8EBWU2D62p9x
QdU6/CrWKhV4zPj6YpwohTBa58cy2TPy5vNsYonbyi90PyueEF0Uk29uRXFh9qJo
wMLEFBUb2m8fL63ZrCLMZ9Qx64oMifVDTEp7oEm9vSYdkBbbAaFA5vnwDCDy83Lf
0kxprMFgUCHyKeHZznX4xXUkDMfntOoUZwMkAZMxA71oKQ0Uc/Ks+8NaTuJr309m
VVIaNWApRj1YM/JcpSsXGGcC7vxb3ziTOHrNLMkKHtVFbeGaTLawrhXDJvbn4vzn
T8DP8QfqVyyoh74HOAOeC39FhzFsX9ZP39lT3C5G2wBpofRn/ajUiPC+iqYGXTSD
LL6Izi8l44FKjdnkRte0qKrkBf+6S7jlGOTKrbLX8irEJdYYZvAIc09cNDLk6WIJ
lx+TLSxp+tyjgx3PaWgZTL6L7eExwPVvvylO4E260YuCke8GE/aw6pJ05gno2Axe
3lSiYc2KwckJbNINUgXyBoHqRJpBFaCKSLc5HT28+4Z9M2hfpGojd56NlS4W8Q5u
6/sKCxvUfrlbYXKuFzp81bucVPPzFqKOJcX2g0UjVNPIeD6+GeM+LGo+B7JP01iY
guPwr7wiPJD4LOTSKMfXXAJz66OtGKNTa/cGXJyZC+aDhxSowDAOj9IPfl7yG54d
l1HkehAElcK0ExROM1akYS/JjH/lyEycM0Un9MXP/le3qZUamENgFbNXHf/MAqrB
TMkkFFBE53Ky0HaZ2TfjJbjRG3Wpaot78GccjIao7RHVpLB+m9Ya0Sqirc8m1tEt
J4vAmKJMn4BchJrgZfCweEL9PR5TQIR5WQU7OrzX2pZWaWjKv8dbTh63L6AUBtVt
r30T84aPN9gPPZvIRtUNu56l39xwjsbaOHbF58pRQqeyIwPuXaiVOBamR1JscjaG
DLopdfnrGX0CG/kIAzJxooBJwNj49ltSHWrkdjCoFS9UMh0iSAbDJU3FesWsgzo2
KuQfoxrDXDbJ3k8RbQtqnUl0zvNNVupcHbx4MqJQygL35OlIrjjlv98ZxJ+G8usD
snC7vM+Bysk9/u9ugim9QPXrKhUjkpVU+08Ma9hjZcRsSzyyNZjFQrGooA9GKYaF
HFTvZ+rzZ+m6C8OUc85QUc8UfnDGy9FBXLKHyx+dblThES+nGk0s+BcbJwXx+bxl
9UyUp7NComoKSuLMhJGCMKjGWN3LKV5ShS5Ke7xPkwl5nI3r9SrJjyqn7HbC5FOH
/cRDrrdwmzNPZn4ATetykw3VuqsqMcLhXBs8LLHmLDDkk/gsp0SuchPiASHUeXRG
kUtQ/8pkxzEii3usf6IM+Amz8NT/PeZLVxlIVvH75lqffLRsJDWBSoSHNLmaWvhi
54s0/Z+5YZth3+izzhJW0fkjFfptHDb+Ppo4cGDRNg2Nj5UNNyKhfrzp2aSbsEA2
Yl67H22j3oYXDgDqPR7QLFscTTbtmpiduAFIaH9QpVZpVjwFszTse3B9cxjNJaJG
74Uru6Ke94Ip1jEnSxqOljvsCKAa5yRpEpcZVuoffJTFSCe+y7fs0SncNqBPc2I2
rmLKrbojZnxFnhRdjM05W1pbfaIc9IYBnCJB5NtXjcPwkj86Q+Cu2+65gFaD7Fhq
r7MZvB8vdh+qMkYjmHkUhqugXTKw7uAaiXpIXEfhKqIL2pX5kqMG9rw4gOORzVyy
254xcaAamBbWib0FczMWIfMxYWYYMKV3XP5mWI+eci2dCe1KGyKk5ZJEJ0nvGZNC
yW0QjEL6w+D0qxZY8E1BBgpQWDDfyqjJ2Ht6709gaM8z4LxegYa86aZ7WjQ2SrmY
eVZZ3evPEii0AhgiOkocMkFfceE2yQntpm/VYK0z7SFmNGozNz91TppsjkJymXrW
EzN7YpDV4avN06opZmuR+yGim4mslNhKvqcHZ29M07xDU5bUn763m7PcPADFXqM7
r3ZKAR9/n/xcL1ue9lPUGGsbZ9tpoLRcgwrpVFC1JxwiktBuvgyPe3Tfb4MRei0Z
qRXqZEXbq6fUNkSkwGjq6REQC1aXuR57G64izGpk72fVIOcYMYePMr7IJvhhTc6i
1lf/viv7FCUU4sT2W2lFpm0AYwsXvmzUKchc9wksREVRu8zJm0J2MhGWWBSGfj+a
uqnsaR4BVQm7i/cOkr9muiep+yj4H4DMpHkrwOgogZFMqI5oGZnk9n711JWXGt0u
ybXGRanp7w2CF4/MHseHW2eowp695LwFXqwmyMvGzpWkwnBBHTQu2nc+WAMsjCcW
fU5YkjYSwQ97Mr48+rm0r4kOEwWVFcHIHDzTcPsD0o/Uw7OnzkBbXcyleoxd8ziZ
QNIO75UkpLYAubvELI5wjQ6WznphbJ+VlaaqWh2LlJ7w4ngqiJjJcUhFqyuloMMT
p5cnALJYvG/jm/rwWxzWDclItDTIJ+hzmOQMZM+HAd2gvkGZ3gnsG5P8LIBdn0yf
GJsZKO5I3XF0Uao6c8yh1syJw6CyS2sstuXr7tjALich+hRWmnm5VLGwn1HomG97
pk18fVLXplGgVnzru4XIpQFCbODFjxuTMVB4WvLUNTwKdEDbUZxml+gbMg8yCpb7
sY8MgIn8MelTwfbg8tErkzh1ZGOmLSb+Vzg/xuwTtAMKQE2+sRKn1ghw7IO3dx0l
zF7F2Janpp8bCt2XVFXWuXBeR5YyKkEU4ZHwJSqxQ9WMhoAG7P/UfwFyTHsXwrlv
Yrw3txjqvYiEcjVdusCH7IkRaEaovmP/QcdnOGyA99+NrSZLAgOuo5esL8Uoh4+R
SRv8bOjhjFVCRU3EDHkX1EX0J3rpI71g6FQRks7c4Ktzt85TtEbDIjV7d3sS37rX
ycHcFynRgLQW0ci+Hv00CES6OQ+jzc/O4ipC7CB3Iu/0SChAvobhekNiLaePRz1u
S16QTZmLv3wfollaxwa8i4+pN0O3g6WV6cl7peKquEjcEjtXaoryIIfk5hPZj1TV
V3q0s8lBuEZqufLBVkOVmz5X2oHz2RZkKBXuw9/+4LD9SEW2ve2j340pSyUS1E0H
tdkB3DsnM6IRf3xmVAnUp4DdvwbyB33NabhcNiQ2PtlqeBUu3NsTEepI/pV/AK1j
vGmeZF/Cl2/mQblQqxi9zJ7oSmoS6ylrpJBV3adzaGfr2A1tK2ukfQejiyo80fdN
hZDgRQp75qADTfo7/m59ZrS8tRwYACzfrQichrVS04qXGLoWxo815sORII+a0VFg
FI5N0Maxwl3aSWJvRqrl6tRoo1xFKsqlQyzjEXkzVv+JCkXqxwh4uIErImE5GZlz
5+91wOHhTE9AwOov35+9A22nH0K/PbUvKzOPe9DaocNjaNbO1mSMoNVJm+YLBaNb
JRxSWSYeK09c6E5GwILbQCIQar4BULq8A22iq2Vtthp95NwEn+bDpZc0DRfEiglE
KYkacKsBRg5/yM60S2lDWkCUPxEKOCCXyVFOhGg7pP7b/vwwQYC62MIqR+/XzIGo
gHECWIeN+r0YJCKmTgNhav5r4kh/3KAT1iL59+ids2U97ftBEMW06taXYTO6oyFO
9SI4tClJK/1XZN8/KwI9ulM9g/0Aj96G2X7NrRMb96CSVmeMl6xSdH6gD+upDvsY
nFN5xXYzu6KXzNamvSaX+N9dapj4SI4V3ZaSyF3j+6hA4fh9mj51Gafmv2txDUhZ
MCrgslqGCs8cLcWvx2qMKCwaLaJc3DtjXZj3UT9iSRUN15IcELw5m6RymDxHi4Xf
1TtWtuuw/ChTI13uO81EISpbASmr0rZEqqZx2BerUCRgnNAzMLdm612hIFaXt8UW
lonc0MIqzYSoLgjDOmx3clFtdpDWV/+GH0x16YRg01Cs0m+HYcPUP0qNRnbuaC/R
goeLLMG+dp2KOFjmiFhQtW6AvtOa2gePebckhvqTPqVA03GPN5EMuNjY9+hl+/eg
AIAWlNFdLKtKM9D0S8LG62rOm3sYDBMDUprWXnJjfv8tvnWYGvXuE695yR+7x+nV
iHyjlX5ZDPzsoalmwiD1Ub+3u5hiluRLCp9laZ1mJ2eeFueoPBJnkPtjZH7L+k1T
W9cn0zfZIrBQ7xlWBaZc2Hvm5g13JBHRhzeZ9Tdsz+Yd4hxegn9Pc7JriofRqX7E
aDiX3yUUkCjvYYwL8RIX/HVHumQ2xCzQ8TqF3rDSwHgkVW4MqXl2ylouMs00juCX
NIf2xWMkNGK+xm9VngIRzTqQocufbMQhGM3HxBYIeuzDiLTImccdt/IxLWJIlEwt
ewOe5HrA54BieJC+rFO5GvXeLAfiTu+OYJCwhe1MpYNt8yzS1YUhINLKDE010SGG
/Kn9+NuWxkFDlIYAjKc2WUObnd6rZJX5g9Y8ogSzPRjM9ul+dNp4okRpIVJrErj6
mh2Xackmu9lWt+vXWeInrEBJO4KU4TVeKxWVAb0toCsbyZBxpcubui5Fj63uQZgG
jMbN2OdcQY3yytUdh4eNhtFiacFoEovf5mgP5WlL2ACeU7HqxbILfl47m7YErHWO
pKMGrI2AvGpW8rZe8TW1+vogxvLyts2pCy5m0azmUA48QXboX/NuKLo9xCVtQD40
lfb0Aksnlm5w0WjfAX3RFsS1HCexjuzXQhWbuDuYePta3dB2C9jrf77CVaQWaqm7
gMaJfChg8vW4soS051cviU0JrxSmvor+smFWDHYg5iAkYGIsZ1mA2g/+WCnYFR04
LEwprXNrOOZj6ZwMVvcvgGUcT7I0yLgtueU5Dfd3zNp7xK/L1cmaQ7hGEsoeLrSQ
3CHcURrbXUs5yJW+mbPZth0Ckn2fMo3dg1tCNBsv6OZxfxA2GcLfpnvyYzNfQh5W
nQfEK0CYYe+RfT7Pk8vgvW7Yc0BueTAH1fd288s5k3HlsVFLl9uZRPXBfWB9TyQS
GWQWw7wZasg2tjQCZv7BVQUikLROhensF84eHgRd9JHf3BeKbpO6RyyD6ISojfrg
1B3QbWXUUrsONBWMwT06JbM6Ov1a6iZNGVANZzOkkDALQoMubgMPgPyAA+u6S67D
DZKtcDYuxy9CLKmx8GqzOjL3dd0LGHDVJHsbzm1VEZYgmJHw0DTalevJv3ySr1Kp
l5//vMc4WCaNX55o88v0yG/Fqqbcmta0XVaae7xZ+ODHorwMuCG0lCpDqqiOrBWZ
4WiiB17GpZODK5tMtfWB2OFZ7FXpO3zgtPWUg3N7plsKNrodBYdUQwP01TOD1czQ
A8Ht9jytyA5u+uw5uKKXTXr0zjOVca9CrWHA87j7tKwfwbDKDOO0tLiZKYHedvT6
lnA0YTowvk/8i7t56KRQxZ46jIppVw4T/A3SW36XZp+mbX96psz9yRG4lmEbD8w/
dLQd8JcBY81+s10ii3zsERKyxChEn/7pwPNA1qM+g1FAfF69FGA83QF7BINlWYac
0Iisbih+//C51T5nZcE/JuReNR6F5X/VWqglFuSRT96SqkQGDDewxAZ8dIcPaqLe
jd8AVQUBUvWy5C8K+HKwCE3eELSv/+k78mOUfRKNLTamN5H9HFj2DDEEj1AJ88Ia
dxeuS/qu6WdlQDNsSzPvwFWiWFI2IhDjHq7bKzjZp5yHZCob9SIraNh0VMxkpt3a
VLLqLli8EUZG88Rhu0nWcNKKk7xlhxv25s4EgQc/dpYyqP7bQRVkW/Sn/PPFqYHZ
FPUSkQH5+Hc2KViT8TD8sppRGsNhpfTRlwieSds7m21HggjGkpc8Q9Mx6DNnwVPb
SxT40DB0ZGJ+UbCAxfR9Ywapw2WCiMIz0ZTm84SGo9r0lvE//O6jMRmwuU25X8D/
E/GB9LpH6qd5HLBRJM1MKj6gjuvbGSWaGVATvuyyVqnymHCsIUQCBfP3auNs2ljC
Wc5HJTEFOSbqoZree1X3o1V5R0Jr+uhMnjfy4t5ECofWxIQ4EqI5TmM6RBIh12kR
EQsU/0dtRj9Yq/o/bOu7T9Wuq9KRpE7UD9mgk8ItOWirClQEA5X7mgZbCy1InDIa
3tHiWHiZzOiOCq/Jt5IzloKwdI3LTgrIHvKitUHU5n2T++kkFf9CJhq0DA7r4j2B
S1As/dqJjrI8NmJbC8SbWt+CZ7+84ZbTOB1KhJKQ2J3LIn+9CV+dDam287tQ8vgs
FbHyaiBLIl+BhLqsu4XKh5pM9VNW+OegI2N8WedSOMTP7Mu4txQqCrh3XahzK2Tf
0WJ50DgIn3wsRiBRf5UylUF/RwaA5wb9f2b/oXFb98TJjzQ8D+DzVA2Mn0/EoD5Y
SaQPJdtGzCeN126Z4OprYujPWC3SMmHVbvziPNF480NZDelGsFfFSmL1iqAraxxR
eTS4YUK7n4g1U/4L/RHh9H8bwN2UO3L/baHscRwVslL22xyXJ7mCp9yisGx/NrdA
bfhj/6EagpD4rDo1pFbiGPtrx8WEf1qufumQLStmp3coLBOLDSMwhjtdZUGfffgA
Ihp7taswDhE5TA7pQDMEj2PNrr45T5nkUBw2YEySt8IlpFCERTwnYPpUCmQUXE80
z8aWQUSDbNQMqjEY9g6EMXFnlC1NlWLUv2mlQNet7K8I+Cg4/4OQetg3RtVjX0Ue
Rf2htFtjw21h3fLC/LPHLx7JYxN29gCnpwYqUT0rx+u2adKpGvi3579hyxVjiY2X
Sn0egVZnK7nbVqDz46/eTpK8EoT0p7Fa7ZXuTMl5DTblYIhL6WVYxJU56mHAmyaM
8gMQTkYGAEd/kzTrDLDy+f/Y4XKXf+g0KcCer1Igamu0U7c5QBQBGUh/6PW7wOFo
9YQprrFkWGCEwJVIa/zaj7nHutts1CMXsZAo0dxodQC5/h7EIDinP1uPfYHsgPlU
lpQQz2ox9NctAz9eNDA7e0jBh+TdeIgAua/wEGsI/YTLVsRt5nEQaiSFgN/0AfP7
ieDK6/9PRkQBoDVjLvrfWo7FxLGI9xrhhSeRHjZH//++PrEFbGgNC+InKa4qyKM9
2dFMfx+631S5aloAMd3tZIWUPGsEmK9movlsram2vtxGpGUSQho73V15DxRlWVB9
o6WGOVoTcvX+jniFZ+Olb9fxD4QfgOED/Y1kTezSyqhcBytfwlgYo5t2+Bj7TSrU
2K6MN3992Gl/FGUYVj66p7dhL+4L1M/C3B98+OytzTS0cohg8EnyGmJkYGw2HA+4
+01nFBtq0TtRpuecQdJAYcyPCR7mPEe/8gmMOJCuBQYE6siByYn6bXVIszvmfdR+
1hy2yGBDGb4rFR75Dyyz9WOhT7hWyPq5LiA3Iebcp4nnsXhAedIVaBkBLW1Rl2eK
VDWTtsqSWUz9beYo8HdyyfcPD8zYOSR9FUQwbpQJ3eO+rpgreZwDAa9AoOgwmU/6
sNohXpsukYWCD5Rnvqfu4Z0m6OZWXTYvrtWuRCn92vFiWuWHc5LGcyvgvrLUW2YD
/6r/EpWNNW1dTOvmzYv5MoI2qKuKV9p0ccmBSwaIJwZZ2m3rURTRux9g9Pnx5emo
nw/8BwBtTc/kaQHW2l6sZrfqPyJqLjmvEbeJDNKTZEQrMtamXSZ9jen2zGTMkQyu
OmieY+WBvi5rlkUQpsoL32lG6iZheSrgOErRzWy4m7ry+A+oSrPTuu2f/XgusOEm
u0tMuUfAqcRW8jLUC2BUexYRkwewzzgrQ4onwMqiZZAuFLPLIMh/TWbdTVOlQSPq
m4oPatxnbB7F7iEisw2+O4lMZydUPrlBKvNyttbeZFXyrm1nt1oggYCPnRlx3hAp
oezWwxcVe/DO+zU8N46v+30UGwFIfiCSeovnr8pVg3B4hJIM8hjXUdBau/mKnhFp
h8F8rO7NvGm7MSeg4V/ZsYgMGU3b4z2NEf72rLM8giW3ZpdHS0rIAoKyOZqnKnwt
8xtf5epJleKRqD0HVJvHgqdn1Qplp3RG7zBWDJSjke92eEKM3jfuOxwI+Pzl2+HF
LLdF/DZrOYfihwy9rE4hWR4K0b9hlfB8jcHhrI6XKBevPZwiXCt6k02WGaKSaHcj
CXIWCIl9MoMbMcHWpf0dbafKD74WG8M9+ZfZ9ov/hh7t0+plrcod/48uT3xVt2EZ
gb1RETe7ZUCupDkq54/LKajR4U3EvTLQJMipLNEQJbVFjrqj0KuJzxA+OzmG9Nei
TOLRtZeaqsEkiYt7+xVsguLuO3sat75hhxlxNcBdspVWkKbTLVf3kfEChtlCYU/A
6k28EhU7tNDRdvJLysBthrhdpxdh7DY8pFAFS3LPXPUgmRC1ZwwxDXCCteloGq7d
+pqxbrTBTJheBPzbTuKSz7jSUz2rVm/lJfJMaIW95p+6mC0WP0Yoz2JiqeoewkIb
OBCFgJgVPSL0QsEQEUoPsIfknBC/y9XZjmIKQiLSV79o2tYjmEFPCm0TkUWfoLX8
NdTUKSuGxBMzEdupiBBkZTkKd4zUg+n69JHvIS8gLjfpSM5d6vCKVYlXQAfvKZsx
RDUJxlYHYXQDTPx7t8OqwMlD9Q3/pX4wcxIKsmB04sGv3O3UKXLLUvBTlYMaH3sK
plFKU2Uq4Cu0mRNCFyg8pZYP4d5muWxeSIChCYq9vw4tzNLYlHdT7ic3hBgNmsvK
wv612AY/IO2T6aregoZ3BWqr05tXNG73euyGYS+kTBk6bN6IA52LtAtv6ywcIQQO
siiBn8nm/7Z7vujObdiNVnMiQX8VM22Wxuj2scuzy7XaYX7n/Y5ODxvdFMJrPOxR
57tk5clNyHuvvHgUOSc73al1Hs4eosPTcbXvn8wfkVUTtBRJH2P331OfLZ/bseq5
z8wnseTVe5a5HWiRHTjBJmzYOrsekq10WHC9R7bAa62cgKAE63VK6ZEnr3pH5/fl
ariQtw52fnAqJ58IlBvYIovGdJBFScZ7cbHnwlEOr+fTSmjkYVMIsEEHWIaOgmMv
HXEGFPk894aoD2joNjmo3H92FPpv+pCxo0mkbIOu36OMa3G45QdeGRFsRcpOe8Sg
s/uUgRWPluEtqgnSktio0vaEONjqabofPSzi/HZoipkf2sK9nPZCOhmAWP+5faUc
TCnnO2YlHpDqEEWHl1bsHxXIZJei4H+sonh1K3a5SuSJ0338vkM7rH4Q293/fDbm
mPHa3M2BPRSXrvV+Fe4BOUY3L3MQbd2XjBDm54Jn4/o45VAnpeM61kZ1hMVlbhss
7HZTcYjst+4lvtKMMUD1MY+mHd3zRTGlOgyE7P+JoDDfG0rg/1Fp/jDGn8OKhxlS
yLPhWMD82y/LUbekfAeaeelDzxKg1WYHX1/VyVUAJza7q52kyNGPX607xCTGIHxi
PDLpUX2hvzgOWWXpKaADqG6cQgRSHich97WE+UuUIK4yD8iDnkwcN67bNwScE9W8
gHoeP/efrc6PTk4Rs3k+jqUorFGaBkbPxjQe+E90sFPnSQbQbsXT7lclwlGT6zgI
fR/IC4SaQuJXlws4+uWS9Ye7i5d2Y0461iYUNr445OeOCEk02LLGlI9UBNESjSKd
SqsXm0nmVSnOJ+1vBxmaRrYlX3agrLuCM6rMWG4fa6GQnOwtS95F9KCVZoJaSc20
PDdEatC1UZcQhYF45gZPYPVP/hwC0pWEnYpbqT9doPM0fjwW7HOlqE7ZPn2E3zCj
IMavaLsu24vSRR6CFIs9lJXOb+czoAmlATzg5j7R2kinWtIMxUyuzulcNISOV8c4
P1hVnFRv2VmoQNnbBPfy83tFXVV1q8Lv/0McWxPCkFt8/Ax7h7pxteESqopa6zLe
b2dXGalnvHw1b6XpcoF49zrU8htF+6PPW5vBRujvjEWyVMIV+CzedgdFQ7Q705uT
+e16Yr4IohDByCHKxQ05RAFdmZy4w6QUZTrlPO2bY6znMlkiMNJykKXUZBkj477d
/cY7vwmABTBvdPYQRQDXjAC7fxMbY/AJyLiTPSwDuXPIXlNJ/7YzGWbkXP1PF50T
wYmTQGD0hY62B3YL7ceYRDb+FxkJuJPvpCagp92HfKmiInW0guCtI4C2O0eNrhgb
ooK5ZbWJFyQJBfNV7ZxXBOcSiJ/PX9ksCmoGb1TlB91h49LjU+mAlD/OwUx3VtWf
Ei0WusgXRjzW9WMeRg3XmrvfZMZ279SRDa7LjxIpxm1Ajk3BHBGzCf5BBdmD+RM0
/sbhRhuFkuIWysm6fZhGiaQFX3mPThDXruk7YCjcTlLkpw7K0dxrJ1jVmKyzE8Mt
DRqNI3CWUZ/z8rz8fb76Zt+XFq6QZ+0XlupzX+9Ch7EcyzDvCj/ASf3+gAeyxklB
PKGI9ktDSho7V/NuOee5GTAThBYgD9WDNaEaRHRf+FDQ4c5/uAX5wb67zHZ+GOGf
So5y216x0WfvnzhLN+PAAXbRSXrGgWdHlnohJmPLK+Sr1gAuEoEDsep8hfiaTJIi
qn9F4wbhvhMrlEN2/MTNvhY7wah+mNbhUSnoKj/9T4xLp89IdiIFIg+sQXWaLg++
1eCc0cv87UNfJIJ4K4K6+k3MH28szKohd0npge009nH/UT44VDvJUuqA6baeh/Pi
5O3H+lAA6MUGSWzrOydeEL97G2Irn7fmNNgzmcFtOmqqaWN55DkNd3kr2yatdfwj
Xmo6t5jRgcqD2ayp4E7OIrToUU2GSLJZ0qe1yC5+1/bEMk42ei2hsG42YFOwbWxo
tqE/qOXPNVpwCFa8knGenmP4XlqobsBQbkPfHKBjcEnpjzIIno9LXM3FKUrau5Jx
D1jU9qIh9yqrxbZRQzjs5/+67JjwpejFt1Lqx+4/HFCYTdccoHrfgG6S7RgucRGv
WSKsN27jQGJZ7KBhHOA8lE2vB73PNztkAw/I0XOGlgTGAeSbuDMMgx2ppY2t07aI
xK0H4TftDr1EjdNyIY6Nb5vinQFfh10uKKNvERoj5RTIdwf2o3bgTc2TYmF75Ifb
2aG99OJpRJyo4ovZeAE8XSOM1OySa3iS+jZ+oaJpWWzg3XME5bgHUV+ZHKfP/kuX
1na225gqnaZ/9vaTauvXJmGwoVyDhX3xS4YT9Yc3xTUDN5v5ZjhHASwWv07UgE51
2gAvtCIn6it0feN74jACK6ipCbakvxlRFZyheA7J301Vc2WbPkCwfZJtepO/kBcb
0v/5Ft3rKmiZfcDWIj0pXve4UBgm/LXHfuIGhMt2SPbA/mNMDgSm888LLQjYmK3l
6R9mlmLQlp/o6TlwEnkwbFc4ysiLrHD61C5HaZHteoWYjPQdj2LxgD+SFGByDmjy
Jywc+m/3ZGDbrxEsGAFR2L90t4Ox4xcuGNabSB+zpJq2wWBkAa7Q7jZWsF34FRir
M5OZNJvJhM88XhVFwfUj6j80FW4T6KOQy6NXOiozIrJsyQ/s2FLJitwZYOBR2XaH
FETOXdPk+Eq1MapliKy+qO3rvN9hyxmMdHn+6kuNVwPT5wnJCdXqBFkaEwatvARq
AvRI5IVyGhKnLwtfnruzME/Z+NPDzeZHLniA+LZxIpmgudC5EWhG83TMH/fLhPX2
dlEkmQpNbk7HhaWGlS9pa/8RokZOURxn6F8hdEkyTadRbT3DPgDyzW4TjuF2I0Cl
5T3WGK6tIWG0x+sl/BcJthjJGHlQvvyWJU/NP4NdF5tb7XovmFzjsMd/fOoxK1pl
MnslDFPQWpdyV4ANQ+aIWOj85EJZRKfHyHi4ZqG7HqYEK1v2+E9Ji/UGShG0XMUV
geIf2VPZsFJDkoEWjCH8P1H+0MQva5/OPdcT6FI/+eB5sKm8wP0zQUAOr8EMaErH
HnK/Bq4hrZRV721YTxZxIF3vYk2Ya9oYdZxccjpwt6G9k+Rwxk/70rcQT38R4bl1
Q64DF5TGyVW3z5/0fwtz2caT3M7/pWp2/uIdlK4979Q6L4EP4nOi7XkEHZPYFTpE
JcbEnjBLjsCaMwzQXyYEnoCq6XdiF6xhPJ55S+15xMj/OpiViebExifFUfzy1RBA
1IVMXh3qdW1rU4Kg70vLDYaNx1kB5Utho5MK2yIvvcYSkP6GaE8D3uHVaHGK8FEJ
CXiJxVoLzv/v9P+H6qBVINR2/k82w/H17NFFT4iSRqKb9wZUztGDoJLeJWba/0v+
kjNJxT3UsS1j6zdAovhDgRFpmAjap+u5dwvoObEcZJxsOLYRraSpUK5+yax8Zks+
Ys0Wv+gL4+94STEqEcTvkoZHLaTGgCjXL/yY2C+CN52ou4s6YYLw1ySzcC2Ya4V/
7QYy7E/gvuLdWqNgB+vDA45OX+UR49t12WEyo0QtlXtHjIeztVoQnCSD/qDzuq3b
ieCTaP26bMjnrLJrT/qwFPAV0I8AyaZlszLFoiNTvH+yMbyEIZp9iZqMUD0QlPnx
hBOntMV0CA2qiae/AXqcHjfYoKk5XOAIVr3WIxns3WeqwT0pb4zFzbWznA2cAoln
7ciVhTKMLf/2GlKuBH5Kq/U6UFzT5Wnfc2bMTGVV88sAgFMoV7l2golfe2meldRP
GTy9t9Tt2d5r8Uv9+Zz0futs+M6ArJ5YSeClAHFJUOn7+YjNnjtIEdVpnFIO9NFH
SkuJsfktynwiZWnW18pktBuUCDJeRwjTVhIz7uvUDD4TIV/FZPllIg6WOIq2SZ1V
UuRg3ZwnHsk6OwJMEPcVgqGqQ6lmCnMGVIphRYNk/oJGvkAtlwJ5uEEKz0DfrdIX
UOeheSjnUzSY7GpzarNfA2YpxOFcdkUxTUFjcpK/avx1fKB1GYQNQ/4Nfdg7b/Ni
x1Fy7d/KdiDeurp2sjyga6OMMzcSI4rScfwC9H1+1UlSTfaVDrOCtDLFQsVFyOmf
wJ9Wy2J1A6BDOcQCrIcEE46bS78HTNJT44pcO9mVyAL+fxPtzFZeA2JiTHEkA0Zz
/53jZbqLhwdv2nMagWgvtNl+rxbIIWIb1h0h59uI23SjtgvAsvbi0C4FaZ5Psu9D
S8IB6Zg7cDcpdEEwLiX8wfmqFGI/CyZIbJJFxhhnvmvlkvh3Zj0IzXuYXdAZ/z3K
TRFNpx7WYsZMCoYhj/zyMlogq6Y+ddqfooeT0N5IIljcGj4exK9Xj1l5jrS8twQi
zbkC/8TsutszJAyGUdLxDK+qIcgzzY6s8rC3jwSqYkOC6n6tAMPtAJ2iamu0kcQW
RmrPTMskYj8FwO3ov8xgkRnvs83qXGg/tNMVriCCaSJZRkXqi/l6nQEUsHnbUVYd
aUULhyIvmsb6e/Nc4LhHfvT3kqaqDX8gOP5+I0mGqRjEKRrhkCacb0fzDOzdUb7K
SHIrIC6hBpXm3pQ+8cmP1+OM7Q4UEheMYyjlmozruhuf79Vsaj1XgcjouwgNjMWF
Cb8ZZavKfgfgAy0Yur5IGz+7A8dTb6lEvU2LxU9NficdVD0bjl9/sI22g8Wfnzq0
Xsf8aiBxLxMUuEMmgRnQ4TVkQjO943bQ02bv+yqlZ9Bip/3uGxRfX4eNaBrbzz3H
GO88N/rET0p7bKrAArl2h9OZ7NIpHifa7/gFLnHmnZktSQKTCFWDM+yd5bFg5RBw
H14RVqyf1BbOIXTvBZ0V8SavBt0YzaBnZeESUo2r4c62JAssrXSoemPbDNQwPjpD
fRkQXuw5Vvx7wInq9pFDPCZJK0ML5ucXVvoBaQBOT0MY5yEbFYbYOfXHshATDNbo
0RxiLdEks8pqiJp5Mlm0lLDboynGtnXIPcyy01fRERWeYuJb/ogzQtpo3i4uW7yG
Zj3/JZ9FbQ6VIPJSAE9Z/8dyk0UaE6o1FU1V2mRuwN1v6n/SOmxrCYC4XjSVz0hY
r9Q0of+1iaF8RTCQS8y6h7hjvpNDlMJQ5ra0yXaeUfxaQXWpnAE2kvHJefppiKAH
VAcy4ncSJxY0W1B2dU4tvlxt/kyhAPafnFne6r2NfNFhDHZiQeXD4y8Jw5kzhpL1
ARzLsFWZF1rDS7tdmwkn/m21IdmIB2Ra7AKu6jm70pc0JKyIIN0Dv+J3qJbBc7c3
vn5DoaqIIJPCzvcyjF9CrSBp+0YxD+oMA5EMJu2Frf1Sm53koCf+epQiV/v1VBgl
Yw08eCBfl97lrKJZ2K3ZuFG25sivcIvPDM9CjM189BvhZyek63COgjzBzxpgvI2K
tY5JVkt+mKvZVs83GDZ3L/SRC9GrpGju5JAJ57CPLicvS8+4Gx7yzmtNIzSca9ZE
KNupdB5RZdRiVWSkZ4pHv7FodR1wFIaLApuZ7IrkRatuSUY+Tl8AYXvH32QUKPH4
wiOSiNxAKQLHZEo/3ktsopMJgtKkjJUE8CaJr/RSHMhb5GvwPheX6VhFNwHwngsD
RPP+3cslGRwHTXHRBLhW0mXwewPi5VoXZ+nTFpRH2gYwtKJNPfreI47UAFkIGry8
M9VvZpuaw4Q8WcPcbhYgt8C7YprI9qEbEA86IdktslX047GhXkWbfAjCS7Dl06MU
j2pcry9R8MCZTaKB0jAsHo11CqoxOOBx6Lz2A5bjMtR7rYCKhjdrkEwUz1EPhlCV
fJkLs5PNhyNrJugAuh9m0BXTcYtEbzh2TjchusGf0OrSZdmw5Oyq79k3snQIL6xz
XrV24OQwY6Bmz34brxiQ6DrXYn7JQqObWUr3x0765UwZDLrLM4HdhxDNAr3jCiO7
Iu8KASGY1j1mxPm5axrIfHk8yZa3kV8sDEDo2zXeCksnKDIo2UEtRo4Pxc10AwEq
ahO8Mu5n75+twfTWEw9tgq3rNdItF84LqqdL3AkribT5ylv80xweclOadORkUWKR
8zusPaOXoHLZEcxx6zs0YbBVa7Kg538u2NtXv8FrJe4ZrXZpF+MaqunoWA2bL282
PxDAEQ3RfrphlgywUDddx02d6fdvJwgiys6LJJ1QZkExDUa8n3N+Nlil4b1w7HFK
gQv172shkYk+Aj2NrComtPnkoEamA+KJedtfzjeLa8U/rTJdcEJD42IGywA5srdn
iyD2fVH9KXHwV+7e+ElBSlGdyxOjQ1tdoJm+4G+GbomtRrbdLdP+l2W0i1TcuUCq
JoxgXlIcXUckWrPHMics93QMBspHz5K1hzIPQxPEFNREo1JLX1cGQcmmzBG76Njd
B/FEa67wmweWMpUCkYm6pa0/BQzowbOVBlKVLSybktNaybDZ1bNWDOlq5gunhnHI
dzL0kd4xjvTygNRNBtpuHSVvfCDtCnt37YeTMigm1zVrCOlqclZxEvkosOm/ibp+
NgmFz0NF9bdW8kYwhYahqkoolmRnWTCI3SNryWSjBs4bX3FlaSg1ktYfQTKGxSi3
IJCyrkbvVOB+lpDLG4ec07DUQexG/yVmfYGl0EJK0vaxV6i1yc7g71+lpaB63jKV
RMKxoBTPzQJTmnzr66o3JOsO2MRWHszo4l2KybT1cBxsiodsDnkfQaJwx6tYm6cz
fbY4Ju0PMfjyz7/fLbndNWS9f8Uy1ueFE75MZV76kB2dIZz4po9XMgBRzxPoau2O
W+ruqmt4gKsHPiQPGB4eZbfENG2kFBJA0wr4vSvPY1ui7Ibfy6hJQ0i9q2U0brCD
FIUYt9c5rAAhTZNjZwLk2v1Z0c2aTd40U+CVVn3YngWn7VznPBay3EqKd/UZsNXZ
whkvIrOm9eJrwqGPUTw7Qgig+NBA89qlVSjXrCWZZ5admhp6evDBy/Yi7787yFu8
kgOzC2GxGme61TtwK+0icB7Muiyp8mXmkCUMrrhxpKJmrGdhpZmlIuV4GUR/VEKL
BEkRevB1B0FbK5bMhEAzaDyGLx3WF1Qd83IKR3SH/kr+vdjRTbxNqk0yth7LdhDU
ZlpM5aDdh/HJc/gxjr5GiKEx2QSE5fP2dChES6igBvHZWmy13MULUAP5qOxBswjz
jQ8B61R7pBQv4Mw7Lb2B0pqtY4Bi49XnEvcmXFREoHIWlVM902Z4dPVqcdO3RwOB
IsydEknw6BbAu+4WzIyHfqus+HzPC9/f4TyvnYzFCQ8LzsgkjakzRChHnmxjMv16
lBD/WMOXXmAy9OC7uRwix3bL9UbC6E0Y8wjQcEZZmp2HW5GxGAyrCr2nj13oiEbQ
WRetUCJz6uSOm0SYo/KBOQz9S1ZfpcTD4d84kJO3O59rvbao3gn8HLniy4YTtbJx
0nE93xZ532KMLj09bMHyLvkZ0778zHHNgVPUBhNaDjtyayvHQIcKiAtVHicMFwXo
BuDjvuZ8PA4u+AZitI3eJEOtvZc7gbxlYZRTes1mVjXA4BGPYu5GgaifcOIe4HM4
jPE22WCMrG2ut4yYGC1Pe8rk3gta5y0qpwUcOh2otDpiKjl/9v66PM3CfhpDDJTB
UeyQFwXrkWfRmW9TStJmeRnLOG/wrAUuo4G2lW4I2+kWqaUvMv8LvGJeWQ4+dItR
EqVbiKPPPg4Tidq5WLTXQ48nX/6xJitVrXXntm4Er9EoNPuyyqaUAUMRgJ3scuvN
bgeb3mOkLk9tK4VpC8bZOUlu21tx+QAXhX95rGcTiivqTR+zxW3xDMFpbS9QQ9lU
BenTat8Mt6PZYh85fPOepSKaXathGQZ6yq547ELIysBKqLuZf6u3gE0mrsDu50Xp
QkdxsV0N4COaYCYCiGW8gsdv835L19AtpqRXw84uB8iTDWC41QGJzBSNPZhZPGd4
e1Ar8vaP1OouGo+hl6cqrTd65vfSY1A6+4NI+IK/7M9yIp2oIoPgUiC90Y6DfiGl
JiLOs/1wM2B7Nep988nf9VfUPMDscPQ1q/HraPUnVpLCAP3KPoBIs6w5T/8v7/mW
eqIOkgOvdIvg9i5imNetva6QrdECItr+hkKQ/91HChGqwGSoOSkmRqv8cXSR3yz7
ier9cPwNCt4FQCf+PqVW/EAyqov7csm7MQ1/jaVKA/DGWpCn479fuSSDYgY7zOgo
EpmtZjw4JqGV/n2+cFMk5AxRbzZbCgqBnHfPb16Py7PHbStQnycjBCctD/vZ2kww
x5KfK+0Jc/gCLC5rHsnbGbfkk46RRQmgkkEqDSH815TqNTEqoCtnZyOF9+PA0Z9E
ZyFl9BxulpvorxQR6ssiuiMeaXaTcH2s4wl5hKrvebrnZhxxE5HMbcDpr4Tdz0uS
p+T9WrTwl/fJEcUD/oQ+GQSsRxI1layF1K/e/8FjvtvR9Zs8XA036rH9pc6+gg+T
f1MaLRO6jukwwd4llzpw4I269jSSzjWNhPnA+Sj6sKMXNuGRg5PiSY3Wt7itoZwa
5Zkpi9Xhbptq4Nt0b2dHFq4lYNx06D9jvYv2f10FREu7K3y4ruFhWE+ShXf0XXv8
XHlgVPcZosp4hs4aVdb/f+baJOxa4LUeh7GTN+zDheA/xsECfBo8cGKx/NhcGEkD
M43p9g0vsYEItz+xXw14NZS2Z5L3KbHxBXPRWNgIod9sVMcVG0xE1Xey5rNxDWoT
D7AGlulBcWgaDVrbHjaHCoP1mk4OrcE/zOgriRSiD4nunlNejZ8i8t7CSaGIy8sW
/3zpw17Eg8O43UvIoQ135xi8liZn/StxdYwCwaQVLx8/dJ+dCh3h3O/Qw63bYh8/
vySW2yy8tTS7rgPl0gLEyLNVFytJQl5ykJFrvYcHLGmsOgFidFKR9MBFJ3lQa3fI
8HSpiEIzhEe4j8sAzcQ7AMqp/Wfy+8MbBMbxe39KhAvtso2934OziDsiDfxpyC4D
bJaelVgoXCCPMLRXdt0co/NYXIVe6SSG+aJbsMFMsv+QiVcyHKyboIhGR2G2Yjc5
QnhH+TLn6XcUO5BfHnR0X2JZWfN3wDpj6uogoYSlOIDhLuCAq3W9G6YgCVZ0kxJa
TcQCZE3qnhUKcqgA+k5PvSNNjxVBrHrWlCPZvQbJySlVfRYQcDH2hM+kvxzFxXwD
ej0lUmguVh/TR837EQXWPtAi/7AuDU5NkHoW8N0R5c0FckH/bj/1LtpBZNiPmYPj
xmfXY068DtIR9sqILbXnqjNm+355rqoBNhyhME/a78yLFoDDaubCavm6zGo9vXzf
dfFP+xW9aSnIE+SDGytgB73ObQncEmSo7x5MpXats+Fsx1fKjOkufCh7Pf1tp3yR
YQG7BQxPgDXizIa3y0XPCiTrLzkNu5jDiP1DNejAuSlO5TZCBz6nIBN35JAHZ38k
YKcAaArctw0BIevqkxLSAKIGC2nET81r47BvOFxFxyYL82Jela1562xJ4988m1iN
QuqOCcmSoTYqr0tsUT/BQfp9BBoKMImPmmPaIXZsljl9vvRi3815ql9ldypfrBfF
RbDJAKJXSR9iJt8IqRqc1DtwHgBBnqhm4VjzKCR6otP8ISSJ/IvXbCVFRkiKQVbk
eCU2W7yCMkg+d3NoBjy1aXkHZYel7EACUiq6mF3v1Df1EDx0MLn5hO6LA+i3nF2K
SAdMxobN+ASXmlmqtey5/wdbZJNuKtDeXnTdm9Z00rDd8V5NmTgpuCP/qlfHcjcM
3IKdTpd3XzG7nem/XypDBbHd5yosdBCQekIkDLDOhSmZKfhsHPIDvQEesdLVPFth
KGoFsDiX/KQgNW+rG1SWJ0JjgElrMZJAkMcGlI+vy6SDQAADM7M1NberVzbvqMCo
kOmuh43fIGyqebAg+xQ3Tu332FdXu+kYdPa3efQr97sLNkUTkANzKaST+ffIXAVJ
UaJo2uhLrBIBIazgF2IW5ft1eEL5S9JHQUlu2aeebgMaz/dH4hzPLbdKUyCwm3/X
oTrIklWUqdovlwT+gcQl1ntgwUJocbcXnF+T2FsiMUmjCPTjCqqBwijYliOxVflD
bnYcSluV5zR+doD1mP/YST9/ir7MfXcxHQWOqUrFTYOPjcjTvecdigObDxTMqIqN
+7AOFlr9YJBmL7VFiDQ6SGItUlMnTmm/ycJfZ3yJq4oJLw8UH+4mq9yH+Q1XMduU
CjO0xuycjCGcjYAtEvS7mqLeH+xroZFvrC6Dm4NlTGXFpiYMprvSGaaty1b4hYNj
NSJiZKhIXR8KZjD1pqcEzppCklyQonLbfjLzAJ9lIVCkKUDE7r2sgBBs1KWQYONK
JS8/Q4g48U53LyUXDUHeNlxGnheWClimPNCWbsh4IElTMVeRNlSUR6xvK0z7UU+Z
gquNM4+HCBX2J1ucNn3GYo4+zaMCHGJAWzQASe2HHZgD8v4Cg9a0hCcslqIGujW+
oJzOho8mHpaTMt2JgTkPdqHsXLT97+84oJpVBxpruXkQz9qMHZkc1Fk5ExdkyW1x
i+6RKfqp4+WLOZgImtSF2qru1VraAF8waWo1qfv4Om4Sg3nQYEnIKo2WMtrQbwIY
3JjbTg1XrMo95gKP8u4XD7unzxFjK20etPI3EBC7C8ZcohvtlTBdAgIlkdfIm3yh
wrTTLiCkmhItyl7AwJWXnbnnFoOtYUCfsMajIrY7Tt8N/dN5yTQfbUzCXcTHaV/5
2cdpPVJwHgzbWy6rw2EsqmPztOT15rgMy+eAjAcrjXISHWKBHCAAqqNZIUDAQ1B+
uOo2Jwd3hs2RDhrXQHc7jySCCeFQsM3aa6TR0TwQ1Pw0sBNx4G0/TS1FVyqlZ84q
J1Y7Y1Njk2KmRIowN88/Y4U4wkre5Ycg0wtmGa+eyr7/UhIxDQugQzuiBkHp10Sa
qCx51AgGYD1DV3mWX5FiXSecGm4Fbxy9QRmWe4mC53TgFu83rNv90W8HUydWWqri
0IyN0iVH88QXlHzpED+QIPfFXJJcpQIjPJndkulBs5fmQxukOFOWlQctpxz3917P
flgnjI8f/47snfMXK+h/lRufNH/jusEUcjtJlYyK32d0S1x4R2Y5Nm+kNKP67bNl
eIXu6EQ5mnDdHdUJJ2a1skqpnX3RjkRkuhF8D2N6OEFyDegXqtCNk57klVpfGpvG
tpl+/lUw5tVG8ri0HaMlgzhE3+iIZPM31NWFjF0kwnXUR2o84aebtMST9Y4uwOjg
oIi4oZistaT2GwMNsFyJdlCK6wyVaKydYMjHz2xuBnJEOI4QcGCSRjInoPYxg2/f
RQ+2hjfGgye8W6xuA6+Vj+8i3K/kWs6Tz6SztXY/DuxZq0pzhlWkwjv2j1pOWLkY
nR2k6CkfQpn4smW8kl2WyeUcWQ5hW2AX30wnstc1dkPOc/CAezbLYK3AxKDcujAJ
2scuQcRcgxrBSrwQEzB4sMYz/3COl9Z2NcRfCIW1HddyH6/yPpEs4S45DuMxYw5V
+aBpbn4cRfkpOn8AAZQjHjeui252GDIYqpjYJ8MoYfIuelfYHvvnip/6kAhUUCBl
Ti+EELT65l2hq1q3fqzAvAUfrfwaBjsA0MFr5gK+NfbZGSAMgp60MMuxkDe9Dv4C
sJHwKRBcjDI1q+Q7YrhUvixd04Sl+rKRsnuA+mZxSd86Sl5y1kduG/MpJ6tIFGOp
yGhyvVAUaBr89fDeo03THU83wBuMfaomNeXRPEsfiR65qa8vFcQ/kcrQTpDb7ppt
7V1ymDZq0sYCj/JLpXqopKDgJzPYTzPNIr2JGkvlcMFIo53OL+b42AH+RWFaj6ba
O2gkczsxiAuClMXrTZrbomPqxShF/SQn7DY/I0F3Z3oN5xohD2gxT3sMUSS4+NVg
swsa9q7cm6Xwo091+ggKtqv9R/QyKdJN2Vp6q/SCrzJPL3oeX6kIXHCFpkt5+iIc
xOIf7amEJ470sPyc7he6d2LAt7O8w0Cee6ZxCsbTwpwkjhV+ccg7JquTC9l0vW9c
IVDEsQLuTkSlvLBpP3E4EYsJT6RIWxAu91QPyzvCQDiUe6suDGM7YzXPcuuk7DAU
kwmFk8juy5cxNa3xDnQGqFkpZMk+8aP/oiMT+1EkJdvLDsm+SJ0v0qiSFxDWXVKk
rTzGQsndq6hpt5F3If9zRm73kF+Dt/x7Ojgu+GnH1Bq1F4F5CplCkr7gRUZlMUQk
nfWJFwYXxyhXX4daMUYzAKaTEcurs9BMd5nyrgTvvI1soGQdI4Ja3xOOs5TdzlqO
q2zfvPxBIC3d146yG3Tn9fXOM5TtQsCiCSrBwfGbkslq99R0po379XS+ZeC+U2Qs
qQ1S7LK4qcwO33gy3sWT7QC7hc4Pp3gMEJwUxtcmq5bFJlpRWgzPDf2TfVvpfHyY
dzn4Z7rXuPq+nuxP9xtG03kbGatnBvVJ+cBWQ8EXvIgWanYAnqyxZL3lgZGKH5tO
PqtE/75t4+TR99f6eqJqJZGNvlONeYRdgw+u626u3q6oQpA8KNcCo0Et9FNGXhUh
q4pVgxtJ+5fQm93dnIEi7nHg+8eMJlUxzhhg3EsUd4oH25Rry5Zz8RuYA31veChK
i8abkAkbmIiw82otUEeXF+iIJRvGwPANwSakP14yYXlvxCfqQbB4mkabL1MS5Qw8
0JuVXA287y8yE+UAko94HaA5smFLBUKS8YcJumzFO29YdDkeZn9Sg4J4p65+RXRr
9TMHau/RGTXgvCM8pjrVa26C5wy5jgLYUK/MgccpUw44YdvsRTk1L8v1EcsjBwgx
MgI3EvnATyfXznMpyeiOAssnOay8furVJ2teYx3huWWQdaZMYjCB3Zp2N/fytHuL
LUBZBus+ZaFak5wpuYsP2Owfxpb4DU/p7/o6zkVwsyy+wCotFrtgaggH7BcWeSFj
fu+90dXEaBpgneXEqdBBGt5qcbaruTVbuM9T9QgxBxkFNCI6As12D3tUD9r2GOzT
bOeKt9vmT/nwjBV3Lxp5nMdGHESIZV0DX+kzIloCyxyR4mLGFwLVgRt4dcBA3EVg
nWf14v4SPbs3o+J7jkJxRajCtBCU2QQpNcDl0GySie8sYLnVh3yU6hEwrE+3qTdM
j4hw5TF0yrNYyCRPblmonV6uWeNS8fDE+RbKA7uGVPm5T4WM6qLvOlQWIVecUpTH
OkQUb29aNx5+t9uzJ5J13eX9ZHuqHyCMKirBueGsePXAbRc+X5RoonmsNTyvROGi
eEmICaoyxICBU2KaWoo5jdQDHOUasRIPhEEBGBwd3ZfVeTjJPLeKUmJtXLcnJNpJ
A2/xtm81yOWu/m/HAstx+J9Rl2RJZsV+fCUSfpHdfNp4/qlgvAII2qehI61K7Ydg
5zVzdTfvdmtR6PWnpqAI9Odp5bHxUz5SpO70dIWZZj9k9tD7VhI6TSGCmRfh+cam
bBzk8o7IPlKkFOZJOiR/yT+XwlHTMqYU+8GjHihJEbrMQfGwfBje204w1Z1hy2Ku
qb27+MPMcKv9nUJtxLnSTZszN3tq1sNgB0T71uS5TfuqL5Be/gidKXKkoWm55pZL
7xZOsakxHc377RlgRMHLeOxEqx2SZ6iqtLi4TK8+syglOIopYMXpJmkjmyzN1qTd
R5Ix5tte2fXwK2k8JSnV8egQ8XnoW3QHWNJWS/jidpxskc0OEC7KCjgSfXwlG77S
4Zf1looyhDBEqUD24vFtJ3o8YJ1IcXwCRlC+6P9TAnwKe2Qa0j71yUomik4C2MzA
rTMdYsHOwaNcyddUBTMi5cDf5ER2LfM34+xgGpEg76py/Dp9PioqmcfHOqnc0awH
NRCXkZR8omtIvuU+GkXzpMjUtbLRj+e6wDvW0dKqYqnkBCVZWRmu/OHIX15vVzgB
v+UnHRQB+uU8bq8ijGCvmBRWqvbbzEkMMOLOzBoXSbBC9iNdit800orwkjVVbnBk
fY7fs0jdKtBrkThh33s2ueM0MPFjyw5ulCDuwQG3D1wmp6NRK/+Le7VJbmuiZTJK
0Qv2Ern3NpokGqgl0wMraTgMPZ0eIFewUBn5OCf+MaqovWbl22uzb8yrPZolKHvV
ZCFoIGX0x117Z1k5jWP1HKiA4uOMw6xPq7FpekfOQDz+DUfTqiw4ox20HPM5L/T2
wUykY+vn5JQ7nwIR+EKndNDzYHaCoDT9ZAzk3LuhBzkFbuoljTM9z88Y8ewJ9az1
4XxPVtlo614t7KqILyFN1LOKleLpAdN4pJmWhCRyEkQsQekorfJ9tr1eD0raVwp1
67HqravYBoEe+UlUZD8qJKd+7kz3ZwuZMbwXDfMOCrF7tOpcS8LbDdEt+gLtCpuz
OFa4jHj0RsRGnHpvZdlS1qcErpNFq9cm94FTUcWaDQIx7UhuVy/f9FBUoKkNWpHm
SrJGKkxA64mkOn5BfmrR4ppBnp5aBAiDWiSM+iaBSiNg4Is/UbdT9nxCt9KeHFv/
koWy+M4z3yCqORFd4XXcTY0Tp9q7M5mspkWEwjyLRPGUZrpfqmr0//XXPb/GNtl2
Lq3RJxtOO3QzMRKDmddSqm/jGtwKI1ZjGIjRlo3bYswGj1iVy6qhZsa+xAKsfJz7
AOVefuaGPLBsizj6a9zMBxqon/C7BmE03s5OfUt96F9Q7akngMrmkbTQcIk3tCa9
F6kiJSinpVBuV7vIptrbzDiWoi2FqYtebTyMFEljG27sd80Eaxl7be+UNsSUYOvo
ADFcmEsOmrkyLJtTUznQ/BwASMpqji7rcBCBkjRi667sxSsV9tJms7m+G1AYv1sv
KbWPpbKZbxQM2Oeh0gm1/uBwPcNAlNDp2AjzCeXwmnXaMQMpk0FD3PIcC+8XKxuM
lYMjXplugYlIzuBnZPlyJuHWt1zNLp9GPu0XhQhWKAfzuutr0lXYrzAIi0L90iFv
o9cJmOABgSFd4uX5GsVKnuEmRi2kiMEaP2o2nD0xsFrKi7bJml9l2GPVAXBtz3wT
WWGyfD7FFozoRiHSlI2GQ7nA+ICp+xaxv0NbFcCniO3QU7CFEFNNZtGKK8zH/Jqj
8OlLEym8/JOaZlap3QtG0LS3sYEveXiQOmNNgW5iT4Ir0g4CL1M+4bez/BFcT6jJ
oYDgePU7oAwxlr18cQgwi84DnW1AsydBew+hfs5Pu2GLC78C+DYrEqQGlizh9cnd
WUMub9LII3x/GwY8HMMkPn5JwXNavODcvFi1kCBhMqILMey4uMRVlLB8Dae6Cn0K
BXnBMRr+ns2yVJE9s4uZ4LzKEFrzdXYxaTd4xkzVISB4ZIRRt3Z30Z9+MDKHNbqn
B99FOwzM7e0bbGMgGpRDdsW6jxF8BZfwQ6KLugYOLfZtZlJU5Et9P07e15xKVNQ5
TorGJamkJ8LDDy7b3BGqD+I7grdIflMsa0z/ztr0QUopLZAAlmINDaW5xJBbqruv
UYhuVWrzt9hJOqBTOt9BvZrektjs0lTHlWrwlhGnIj66VnkPT8hf1Ks6cr68QdWJ
I0s1S1HDw5cBkQVH3fOxVB1A4yZOnnTddNBdlpTcWZObVOA7pZk7BkCLauv5CEMn
yoLoEeKZNHbn21AialZbbNs6q9Xw7R+tWwBs4nfveIYrOqCZu9lZwb75B/hlwtSh
QLmoKgITkJKv18psU8PZ8cYRrAMCQAUTdAIBDtNnxMSm4B/FwNd/pbtOI4lI3Z1R
UfEErzjmoBO4Kr/2JCraiDeoGrMn9ZhB+cPghV1fiH9mHvLpz7WGPli4+P8tTNIp
A3eeBLwP6TjA0ocXVxm3OU3dlklvjNpZUZ7h047tU5sceu61wQY+Oj/Rjw1ciZlG
wHGbYq8I6ohzxPK0gvkrX6dTxPF1m4v1uG02JY5hevt8ct5ZElxx6LhmFvu8Dggn
WgyK1bF7di3+xDR6N+yq93BW5I3fZVbPyZQtcwCegw219Fx832mXeJII3FXZOtVF
qcpgcNKSTMHxmB8DurP9hQ7eSRga5KuAAuEAXqFwIemohbbgr8icyy+3dgEZlYFY
EBSD1YuSYmJP6RYASVhkVBBSfSWheguKDWHW0kCBLHyMlZUxOXLH14I/tHOLbsf2
CZj1ZV2g4zT/Ab2SpHoC3GshGel3v2gr7dvLUi7RP6QQjrrd/bO8vuxenK0KuE1t
YRbbjQDAegehQDQUshxHpUnOerHColKDTWxJ3LwUpD0ai7KGXpmOm56iEmo8hKxw
87teIkJy7bM/opL4QXN+a3+uvm0aZP3qLeTTHNPbTGNNlK+79CqYXgocL0JOIrkh
canW8ddQj0DZZsAx8ZhS6W+Qg5cFwGjE3t9Dv5aOU1I1uY2nteuE2V4sGMyS94W7
bldd1WUoAhs+Dpt+BiIOne1BlNPA//nVoCIxzv/QKyNPkWr25g5WtRBj8iehRUxh
Y0LkKrNS/zI8rTMAXanyPUTNa89eYfXuoeLp6XOEEakGLJadxp9eQ1uMEaSUw7A0
hcswbxHaTk942KElqZUsOn8TFg/CrBLiDjgr28uBU3QN4BWn/pyNFel9qFA2mCiY
9JfQDQVYv1w81R3wAK7tHqa6SrbrzSh91L2zPoxaEVphS+0ofkev/dV+aa+fUadA
7b34xzPzGqOpwL+u2VCD74D6wNu6ZewrECIU3fdPkLPRLRIuHiuh+qCAbZzrRNh1
K2DxLG5ga/0GfRsRKP96Ux0ZuQhvKGq+5ELZsezLs0daD/RUinBr0dWzgm1Ft0s1
AvFFMM1Rzpnw7zVW0F4x9RtFJMuWUeNR3Xvo9v0GXsww7u/2h5iJvHxvnSuFetrU
Av1iCHT67R0mQtvPmZq4r5lpbiTxX/K9dIa6BChjvGMuOT1dSdsZRZXtRllc5NbB
n937/lJgSM1y13bpdRqrAdOYjFF50ev4vXbJRhy8pK78TWllzK/sdlheAO+BW3Sw
EymV1IMljMZ7aCGjV/5mmflP8SjxyuzgYqG01ROWF0z0EQujTO4TFXI6wJjyTpI3
rN+g9t+fuHQcsWCoevaVD4C6ix3xZcA9HRYYpdMvDeeWs4FpvK2JMnJYwIm+wV1W
ZdILf3uF01LzwXhVkBgSW8s/pu3C4i7ukeWulRRhiZSV3uLpvTpiWX8+CIqRBkGM
NfluIAyY2x30hbEURb6yPKomWbNyuC7zhrZXazXfccsP7EUKNpyz1t+uo5eQTPZx
eZ0xmDMlMk7AZeP8phUH//FnipgFxXcEJvbNmToT/b6tfP5WO33fTJMW/wn7wZ8H
dK3j2Bscoe2WaWgBZt5GWessUX2YYpCzb3BOrZGmao3EM6Yq/n5MEbPH5rVSd2h2
MEQLxLxxTBYqi8rQ+iYUi7XKscBLYwsGFJRe7jExFWPjFDJkvB/HBgrXK8Jq+Hay
7LJJ8jA5vOllSUN8FGFBsD3VhRfCrt0xGB3fxcybS3YMUnkO3ohE2yq9NJBF0oUE
3W9EP/fQn8duQuwVRKgroh0HeNF0tY0tPtVJSso7YiAYEwvIkNJHrkZwhLX9hXOm
HwBT4I32Hx6IkvYyftO0oe9higlxOjEaNUrZBA/xXPK1xqyk8jMyM482sr6qrSCe
SwxgURhXIive1S2bcRDtU7yfIXPrNSRpkjp0x4uYtShy7p6HcKut5QjxTGdprOqW
g3Aemm/h3hVQf+JWnCl/o5bQzI6MCAeHS2G2fW411ee94Fo0WzCzu2Fof9tZLiXz
ETzP8ITP8A5Zw+B7L6DkSpJev96Gc0ExPG256dN2u1s=
`pragma protect end_protected
