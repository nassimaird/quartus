��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�APq�lG!���h��2�&�M�N�5�cµ&�z[հp�F�/s��2�3�%ȧ�4�U���G��V{��K(��.�r<��W�$?g0�f~֢�!��oG���{�p�4!�����
�D:ෆ�iG;�m��2 �¹��J�}�?�����s��@Ź6��h/a$���pm�P��FF �:���Ȓ�3� ���z�W����A	� F��ǳ�ԩao��Y�W��ubu�mW� ��(�e���7��x��?� ϋ5^�G�T���&U!h=߬��sNuo�D���g�=X��Ϳw�:fK���53~*��d��>�ՙG���e;�_V\�Q�]�8��?DPc��.��(f�{�|�r8ϯe��ƥ��&�l��H
��KvD�r6��ҁ<�����'Qe#n���HU����o�%�㾤vV�4�
A,��  �5fie����G��S�9~>�p'*�xZ��rp{�Ă�܈mq��݁�+ڗ�Z�6ZE9��3ᓵ��]��`�d�5H�^ىn�����X�[E:uuZ��v�p#����Vq���c��*�,�jܳ$�{�z`�9��k��mE���
7���l��=��U�5��P�T�	#0r��)�<��s*��A��(Q�pTų~��m������~2�%r��8h��A)�������ٲyz���u���;d�k�S���r������-����/.R���5S��%�VsO���A�rDw
UF�L�4"9��:��&.d$Ш0�g�jط�ߞ��3؀��ξ���Y�qnjo"d�Tȕ���j������j�CR�HJ���O4E,��\��پ��v~ B!���x�mU����H��F�x#��Od�䂋 �LU�%R�/8��� �Ź�
��,�����9��4����y�fh�:'[`I^h�����y(�]4���
�hD���	;o�Q0^f�#�x�P2�z�^�O�@�j�MA��Ogv��{N�"J���m^�4+=�%5hc�va��!H/�AKF��m����M�Ӻj5������ ̛�=���t:�MNݓ����k���v��<#�1���MW�r�����q��%'�zF*�p����&s;��`*zB�m)F����r�Ƞ%5�~����:����(p�LG1��׀N�Z٦q6Z��xxTu$ 3�u�aA��U4Y��&�$��c�-v6Z�&GU5H��}����C�O�6�W�⯖���.@�Kf?�H*�r��6�'���l�KGp�`C��ʦ&��/S��-{"�>x�����<nE��������Е�hb-U���ˁ�B��FM`G8�����g��c���0 {H䩚�8������8��,�զ1-�s��:�9X�f[���Fl�o5�S/e�R\�������N�Ə�$�4/x�'Z1W��9�Z2a����G���O�2����l�t����ѓ0�#.o��f�����eFꉱ�P�>���̘�	w�6�Y�4ĲV�+6F+Ы``���P�4=y���D��P0RL�q
���j��1m����h�O[�����_c�V��1F��\HH��c!ms	�j:'��`��٬�if� ~�����2
���շ�I��a�M.=V�	�����^<�}1�S����� ;�A[e,��w��K�+v�)�.`�S(*�u�΀�xS�UB�H���̘:����e��Qj�.Z��]vU�:(:V�T����(#~�QQN������!���U�o
z�*�B:R���p��
�g�$r�`c�*\�ފ/���p�xz� �u�[e�W��N�=JH�����<H(fO�0D~p��اwa�ʽ��P�-�GG�|���EϿ��vޱ�y���BV>��NN�}4��a7K�Cw���>���kNf�e%q`�BA���5W0�k�0�$�;93����9�v��,T Lg�0� �ԓ����ȡT������%���C����7� ������f�[>Pe�j����������Zj]U�h��eOsqH؜��
�dQ�[J+jt�0"�8MUch�r׵���J�<ZO�
_4cu�8��)����&<ע'�GK}02�^�k ��	߮Q�KRirF`0�{:�Gn!�Iy�wF����Jy�X;B��y�̈GW&x�oc]��~��/ؑ��X0�(eα�H��؄�=�ul��Op��[Nrx�&��$d���B͓������nڸ���y���	����[$��[�6X��L�q\�ŭ�0���Y[p%��5�{m[Sدf?���0t����bOg�Pj�ͩ��E=]7u�8��-�A��U���*�*y_L��7�f��OI]]�^��eNQqL�Q��'�rIOI �7��u��T�G0)����ì�ū2�\+�������!?�p������-�����r�%��������(ȥ&C�d�~��UHT�Ԭ֗rlm�b����,/�:�52�0|n��N�(�E`����x�rVp;�
�+�c6sqѵ�_�ˤ����@�_ã�o]{6,�[h��z=�1�:gmz��I<zm�����-���@�C�-�˕�����<��=��P�o=��q�X'6�,ʑuH��o	�{p�=j��]����a)xZܖ�*��`�Y�_Shdp�?o��?�@W� &��B�\���3�]`W��W`ҕ{*�G��{
�BP`1�� {c�� {� �C�K0^�.�3j���ؑ3ٻ��N}ؼ�'����r[,?��*��3�vz�[!h���g�}����	��'d^�2]��~ѼȾa�>�m�M�I�HPFy:P���
N�)2	^���|�<�N�3��7�- 2�x�#�y��F�� m��y!���X����clf�����7��]UK��s�iXchw]Qq,:F�ܥ��1����J�-H��z�fL�\���ᭌ�g\���&N�[�|M��F�Am���3d�{��m�"U��F&�=����V1�i��|X��h�n���\x�s�g&-� 0���q�|-�K_��d���RA�䬁%��z,Ǧ�QY9͂c�S~�c����o���vlv�VMN���ȟ�H����>lsȉ:_&�ho���d!��5Ж&�u�֏Zr��pa����+I���2:��&[*����
�]� P�3��Z�^Ċ�4��\���G��4̶�fڼ��PW����F&�^:/�N�9臩಴:�\�PZx�r�:��&m����5c�{n� ol����V��_�T���Ƭ�>!�uZz^bxd
�/6��:��7��hzN]�i��t8�&���>W��)�j�>޹�
�  p`�1oQx\d�ܸ׶��˿�8�1@�~��z(���&� !:�1WE�ύ)� �}�C0a�� �C�pO�D_]"���a:�_�����{\��De�\�bH2Xl��G?�YU���`.��Qo ��5��b�����7�@E��"��:�!�"�4����ٵ���Za1�U�/K�[��w���6e	������#+��u���}�л��9Z���C�-�W��N��ˬ�t,rFX�C-$rX��� �'o�G`��x�zm>�<�i� 2����+���ͲX�Jr���o^�p��,j7��
�{�by��u�÷�}���EsJr��p�a��n�(�N��+�:#���ηڢ-���\��r��옺����F���|JVlX��"��}���t�l��6�>%�ES�.m�:�SA�{�_L��<͙Xْb�+��~�G��^9��^�����7�4�">��d0M�pOh@��}�k3���]D�e;�l��y� D�fi�*�C�U�`9v�Y��z8�r&8�[��Y���k�@6�'��c핑�%'���9�2žd!�	�Y�Vz��S�d1ހ����+�ǐY�a{x�zf��Z�^�us���M�3 3��/���҉�w4- 3�8كoN�T�U����+}����C�{\(?���6���z{kK�D�x0�臾Vc$e��ݳ=�7������+;�V��L��2�p�֨+�h30&f����!��E��9'��{�1�e���|��x!~�i�d-������&`&�S��������d2qs�9Ԥ�̉��b��INCAš='�[B�8w�
�V�a$2�!��2����$%Z<�'X�`�b\�C�'��<�Z��������xK�0	��:�������� 'F�{hY�:IZ�l�:�Q�ڶ�q�c7G�`�x���.Q����H���nu�����z
��LUI�,O�r2T
Lկr�:K_����L�T:�u�O���U�W�B��X��)4{��*Eb��?�.�,����5-F #ﰢ�!=�y�O��mir8>���A r�e���v�"b	�Z� ����>�h������C�e��Qie���M���Bm����Ү^�YC)�N��gN�R#��GF�9��.�-?��W�hn��^9!���po�R�b'^����.���q���y�m��ܶ���ۃ<N=��$2��ܤ����d.W ʻ���3��R�M�4Y+��-��=�� ��]�(g�y�xEL��kWL���J�Be�周�Ԉ��E�;��R�i�4�ݪ����Uˈ�==����~�eB�Ňn>��C�~��}�lL�4�^����E9d5�1��қw�D�
�xHD���Ĉ�QL�
Kʅi��D���w�m�^�n�M,���T!:�K�ؕ�%%���I>l3S*OΉ	�:_ᣯH-	��|	���["�z��i���%*�Է�Zy���ҀNEkk�����]l�=�//�$�2�jh�Q$���"�d���-�o��B��SY�X�[l�$�%څN�'@~��|��L��q�,ќ$�F��Ee.z.�
&'�)'��Ε�ZKM&ݬ؇!��ϊ���Y`3��X�A�42���7Y���H X��PJ�A��ST�A����m�?�OI�'m��x���W7ٙ�AЕ!8h�HEc7��io;8����Ax���"ٞV�'�1 0����/[,9jH>�P��kX�;gI,������ᜧ�Ā�Q[�L��L��bt��o�}`H�(&��9�py�.b:����$�(%�>�ӥ�y�-Y,�����1,��Z#�^E135��A�Wǩ�J���w��*���n�<�����lr��N��J�o[Eז�J���U)V}:�3����� �O'����q�4�&����4+�&���~`��c.o	<�B�;`����վ��BP6�#��O�H�
�y���;���������Ю� �.��L vlXOb�e�`�b�)\�wE��u��Hu�D��f0C�*H��>�*��:�����B��v�{�J+6�� 7�s���<ji�� �*jX��CJ����ة���~����	�rn|�ŕ�	ۀ��=s�/�,��]�|1ЬOÿ�i�������fV���� ��N���'�6-(km��JF=Ő1�Sh�٫X�g�PY�`(i̢��N���|w�܂���  !"g�R��&����@�Q4���<�Bk�L����3�ج�ݜ;
Hocγġ�@YA-�C��]��F��5ЎG�ufWS3*݈!���[$ʛRM�RJ�T�T�_֔�-.����D�zh��wV�4}�U�y�+�|�E
��Y��G�-n:,V�~��=n��elT�`�/�$8��wFԣ�MO��8��A��c�s�����^'Q�E�3\]�z%wm���j�s���/��ju�>��/���|���0������'s��S78"��"cȼr�cΦs�k��EޟĵlƙU�
b�{�P��"���3�zV�L*��PV=r����B�!���$��>��~�m�0���Y���*h-�}��I�r��PK۠O��.@"��R;���#Z�,m4T���F��{�<Nai�ٔw}<�*�����j�d!Q/F,i�����_/�U�2j=����(��o�!�K�	�7�0okn�Ͷ�0�p8#pi�� o�J.��7[t��|��YDV�a.f>���X��������PSv��g �Yy'lB%�O�>SO�ּ�]�|�������)sA�#:�J�P`�����z2 ��W�No��E���<3���qn?���z<���!I�����N1|�7�Kg��M�9ۑܪ�,mu\l�=����t������Ŷ�
�Pp�Ε���[�y �G�����Z�!�bӪ�]Pt�� ]3..��I��=v]�kւ�|؍�jv[�)���M�x��X��^yHYD���W���}MDhN��h���H��BC( �r;.��<R�R�Oc��B8,5��mo2k��p�#�:JnC�iO�8����=�͍�'��˯�>K�����*��%�7�V�\��:��@��9�V+�}Z���>.jz����7�����i����>0�R��$)����dM���-p��n4���M9,[�r��k?Q̆��e���B���������=���)0�H0���ۖ�OTm�]�N|�d=&E�_�5둸;��PТ/�E2�^�������y �_�l��(������N�OLi *}��=Y#�Yt�-ړ�g��x�A�<Dif#��sc�Zy�eM�N�Aĕn�{V�o;�J.�|�<�؟ꐆ`xܹg��m�ԺK���yt����t��ۣ�ޑjB�t(�Q�ڨS��U��i�1R�S�#ty�Fղ�������O}~���Z�kOR�M�=��c�<3V��>؂�ϐ��[E�9-Id�Gj��Jؘ��BR�+�'Z���A7L���!A�+��G�akꌯ��miW7�͸��)�/[�X�a����(�aϴ������	��>5y�K�S�c,�'���7��㎮�T��<[��2��*nd��n~�K�.���{Ů
�x�M e�ӗ
>�8?y7��\H���5��y�SKrR':�5T�����k����S/�)~ٴ�`X'�c�o�����[����)��q�8v�%Qf[�I�?�֪���RY6� l���1��i�PN;��*�����
�;�`��@	t�F����!=�5�f�j��\?�JFU��Zd�?QI	��^Ń����4��`uM�wd�|N�J#��'&f�yM94���X{�p�A�J;z��x<Pw�aSȭ�N/˄��~�Z�^e�E�Z�穇���R0i���T�e���7D�N<'	�UL`e�4�p�,����ь���۽�H�����39U���}�||ر/��#+��?-B�8Em"E,KunD��Α'�+���Mg���-}W�G�3-�~��ѥ�d9���O�a{������jo7�|�_a�@d�����j��-��X1 ��) ��v�@I)63*��-���Y[e�ڜ�w���-k�X��?A�
��8Y��nt�'ZB�GE����M�Q�^��?�D�y������\ã&���L�`���-R�D��<+�d\�F�DH�&���ԙ��@^6Y����w����h>K��h�q� .�!��R�?2ˮ���Y�W3��#i�yX��QD직��1�E�AK[����%�x8KVÙ�,�&&�4V_(y5Ж��3{!v�Y�LH��Xa?�%kOv�]F��d�cen/o�D�8��U��%B#p�O�6�����cF�"|�ʰ��?������~��
�mK�?�1`I�#v/-G�
��;�,�ˢ�F�U��:�C;����w	�y����c�ׅ���QM���Y�<��^yj���o9i��Rs���7���R������F+`�᫰�)���o���sL$��D��&��]O��a��4 �{��`��W1I�E�_�.���y��4"i�i�-��$]/��_���ѷ��%~�P�3i'��TV�5��4�P9ߨ����GN���QL����EO?��蝲��=wm_�@�s��X�cվ�����&��+��U��#VJ�p_R�TZ��ժ�.�J>A�(rF{`�������n�'�T���w�k:K�I{��h�j���3�s��C�.�������#,��O(�o��e񖴢?�d���!�9�dҭ���Я��~<!�Ne!K�[i��i��r�8�P���q`[c�(��IB��TU���������b�2*�h��nW?�P��Ω���(�6�Xi�$JO�n&�3�c�[�݄�|��Y��g	����J��JAb└`���S|KJ�ƲS�,>n��7c�)q52T��]�2�+�o�e:�s�pu���9T���Q��#���?�FG}ؙ��}�g���/`Qyww84�B�/��K!M����C).����֡v����Ċ�$��!�/��j�e�w������,+W��!R��E�Q�7���Œ<]^Ņ%�c-ޘ,�ѨҎ�hҊj�a�����'I-u������p����/�a�)|A?m�����C���[QD8������:*, 5f�$!�L�"?�����_����aS�q��)�g+V�C}�<}�Z�m{M��Pjd�"/� �
��*��ï�j��<M��$@Û�(�tX�����P����_�s�vR�̧d�����8H��"������J�i�u��J��ka���/���@�����-�-v_���͒��_wi�1��
�L�����'����ghg��x��A����s�ob��wv,|4����K����#nH���ˉk'ػ㛂���Q?�	�KK�^߀C�Ǩ���#�X��wk(;~��;	����_�74f3� N��}��H�=���7�P��4j��{�������AT������� e�`:�R�bzd�ѫ"�S����/�|�2�=\%N�Pː����)���'��|N�'r��#��0��J8���J|��qXׄ`������o ��x��e�mƢ���K���8j��z��S�UxW��jT1��^�\-��:�0d>���� �.]�Bb6��\Ua-Vz�`�8	�_^aM$F�m�c���F���x/�8�r��NV�.1<�)�} ū׎����,�L��-M�j �a9��F���t�ڇ�g�RHY�ʆ�.a���<
�R`�bA�����evt@7�Ϋ�4��P�ߡ��P�o>*i�t7jv���k�%FO�wgzc�P[�<�Q�|0J"Tu�$����X���c靲��>�G��IB�b��'�� ߧ��S�UuA�>/{�n�vVa����t����i5�qkt�w�Y��e��h��Z<���&����i Ԡ�"ΔXideQ>�A�1�O.Le���DV}`��`�E�����M���0V���m��5 �3�n��6�O�-��#a3��f�k�I7���_��Hd�g��mj$��<D����.冿H�j&M/U]D�͘��6%�9(���s�̩��
Fۛ�_:��WR���CaM�*���Th���X�\<}�K�n㚱ag�]�iЇ��Ϡ0��S����{�Aĳ��|v��m愶�&A��̛��őL�E�v;��K���Q�4�6j�X�_��+����j�����*�LS�>NO��+$i���^i���Z牄 �5���|^��x�[�tN �&�_x����z�!-y�lQ���$�#���|s3����~c�~$߈�Bb�R�eg��9�zx�PS��U�#���E�=7:�DU
�!��V?T���h}r��'!q�07���}�"�
�Q�a��A�S7ɞ�"�)�<c�>ܿ�Hk���k9Q�ꪘg,_�Y�3���,�� ��X�����i��1̌��eN"*�3�@���N�w�Ѹ+6�*��Y+����G��~���a�A[�rg���3��\�.m`�^R���:��J�b#�EM����}>·5��p�m�t����/s�Żm�V\}O�Vf��08!vʨ�����&t�p��A8���wl�?�y�G`�y\�9y�4�������,�>I�n�?���OH�>L�)����b�)�b��$�H�2���Y�Q���ٵ�ٴ�ĩ}0�����&�>[�2�����|ȃ��"@ñ�H6e8��XS�6�_k���+_�5���Y�-�����"�B���n%f7�� � 