`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RpOot1xyVWr7TwpVF68Bc5RlqABytpdy7J9WeCw3EE5TJLOZw9yUHDJPq1d9bC+U
oIN5pu7C2iLj8dT+6LpHjYHyK0VWYz1wrN71boWyEjhzVPdB+vH1CvNTP1fZa8ea
oIHyvpxF8lgsIyzerAlkwZVXFmpOzC997nZBNl7bGc8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5648)
kP431DrSmIUSIP+W82Uu2GNEAv2Ns+SUPDFOWlN4GgemlK5DlsvyqGHak0SgpIu+
Ljkr98MO+8cajcOYt9P/3hqHeMoKy+3AvKB8swSBOYGhZ8Lf4tqzc9UlVjmsDJfa
7eKz6DCGv4Gt3nUvP04KvQFEw/HMJh3Hu1EhvAjb7yvU6eqItxINjHoOFzIsHGMe
/vtb42BB2P18DNg/tkFp9CgaD3SDf92GO/Ae9oUvrXMmaDgCf0zmuRiMrArgJR+t
R8HXhgOXxdktR36/VX7VPYtnWN09spu+36HeOxqc8Cx9CMLuAk8zDVVgx0jS+0Aq
SzPpu4JjOhmnd8+32v1ODrg8PvsPCfLCJj1R/f51nZTuaPuOtDa0YKXkIx79P+/x
0Eoa6Ti+fi1drufi1ZWYFRA3QVaHapJChnUMQVGo+MHwvCOZvi9n3bCVMWvU0xOb
njbG9i10hMQ2usDvc4VT14ZxP4uF2ZfdkEiNndRcZDJh/8EqV22GagXzd2pwqUSa
gv3Ja8ig68IYi/Dy3Miuzg3BtdYY7dEfKuW8bcnT3BfTgMRrKOfn8Sx4Iq7W+dJ/
c/dLDX4fU/0ByQ1Rb2TJf+yao7el1O8/GceTeyWmoyWpvugBjVISfc8n/SscbN4T
aRI7x9K/FtQh8rTLol/zX+JXF3KGsB9hhTmyio+LYAiasiCC31f3Orz6THe8QYGY
1s8DQ41fDMg+qoqQhjaipgGBXoJCUpA2s8cUaYaiRQSNvJLqwfyAAW4becpt2QMg
fvi/Wc3rSppaQlnX2QVSg2XGhGxPXqyYvKwU/PwPqdvEKuoEicww2RLTlMjyPlKT
0FeP03uKfY05bh1UdCbnMLSi+kVEUdmVnbyYK6Cdb6QjGzQNY6D4R6g7FuxTAeka
bJeJ6muL+CH1njd5L0dZy4F59lUzPBg8NysCAlWFrJNluIuNK92u1VbIgr1AwJA4
1UGvqm+46Ha7fG6/eNX2zpAwk2uhFY3fAe4XDHaUT3l6ENkmYEtJ35b6Cl6VYHAu
+v5N8k0nChFMrvOjdXWFGqJGhxYhtbJy34pHCuMk/70NiNHrwe4ZTSyDkmkhVRvM
1OX+KmDdyxqCNq1jw1q4eiVEDA64xqqTQUyfC0upZ/a1dl7Q3DsgUvpWLiNMUQDH
BoR3uuPnmf0DuQZxGxcab5kjeEw9ENOacL+n+uuN0RMyfAx96527C5+JsIpG6Uv4
OH+q9CP9ltyPiSZ1LKZoibaFkEWSpuH72rUx7y8tACGVKcBMswYu7niD+ORuYrUg
e/2Rr3bUN1JVl7asGfUdcVXcExCvoL3lKES4A8dGTKB8QBSVoNZ/NseXGD7/gEVT
+AZzrKuyll2zWdU5DAOjpzuc3WUmob3w6qqgNNALeZK2dJM/0sCl8362ir7WzG5v
KyLas/Aecs8JC49X0BAwz5ll7jSry+Ix1856QVtnPR9GxmQGHQoHaeZxY2k5U23i
OXxMwgyKMfxBGAq8m5PdvibV70nhE3JwgmfXriQT78Q61Qh/fW/NHYazYsuPnI17
0BF7phnv05TJMt2MnqbqEc8q9qjJ1qW+nrOHRaM7dZNdLl3nulX4yTPOTUkGflUo
gbAeZZgV9nlEK751J1e512UQlVatFWlDsauJZDVeZJXMNQIrXcFcciZbaei37Idu
XS+P8ByLZsER3NnkIZbP+TcLmeL/SQPIssVfi9smle0ivREpQyen+GsouswwYxhH
97bILhkO/7l1vQNrWfe8kP63xG7cj65DMir+Ofxwf5C5HdAHxPSqwLPYl8wnB9B9
Iv29ZMPQJh4fMa8Bv30p8NGN5UMFkaEZbjrrVAgh28T5gTEL024wCwOVKuex2GWy
pc/fCj0TyMpknUCFZOw8xwX0CTl7xmHE117FDGe1YJ2aArMaD4pC0B0RhtqdHUse
UesVaPLnFdx0bWqF8vFM5yCWdCJmnX0GJj0ji5jXZ64COuF1ANNNXVBmOtWEua5/
uRFZ0RosrTQ/gqGvl5K6IfokF940vzoU7ND0NFqudwbWK9MzPHpSwjH33ZFwho8r
z2gBPG+sqTiF/afZMj/Ba7RcC1j14wLilS+ex4BuHiH07H8gWb4d/e9sqLeHococ
qnoawv8knyv3LojHwVoVKwxJZWaWtINMm8AlXUagU9Z3J08cY7u/NTVC4n0GHMWB
HyGYt2sRj7PEsA8jy+ma61RUHQES2rEE3/GifXmT07t/xkU8v2f4E1gQzys4seJF
6kb5EPEmR3qFmzQ8fi8pWaCVeHxW2Q1DB5R2tfYs12tBuXLp+wGsP91dx0L5UEyv
WSF3CGccb9/w50tDf4u8oeUnqXQaf3hTX7p/X/Hh+6PWv36hYnCxtWE58D7SY1bJ
AP9fwFwOc5z64A3ys+uBEy8qieQ2UzHM4DKUugzG+HNPEzdvm+ZKH8Su03hti+W8
pbZEFjmEOAaBsmy2JQG4iyskvcCVXAq997Mk2oo5M6m/PtW6xHqOLwMdldwnjFEp
bQJz3DABm1/KrdA79nDLXWX7varengFl1eIXptULXRODsSvknN8nAs0SfRfD4ByV
VhnrUQRPpPrqcZl0MvNJzJ64h/0+tF099i6pfAfB0ZmODeKhmoq625l7EqYt6qcF
btb8lScJNNw4wk0coejFSbQde5CctP+Cc3cm1VQbeuPmliCQNNlx4VMCWqK+h6Bu
efLVkwxhYTxa/5xVTM8yTpeNjDAD2W75D9FbRPboDaQrb3HWOeXdNM+iScsL/ggU
F+j6Eq3y0ZNl1e5aUsrTUgsDuACCIokDRWoWvpnfCbzrHR5msV6eai4u4bROg8ko
rPx/crgmW7LSwZqhJjkSQ0ufgC14SNVxGkDjYHoEiKzOlTXr0tuQFm5TBSt5qfTk
LpxpJDmXlh3UbiRPSLibyR8on+YTyDIw9oTiMSweH2Qh6iTGrZBrnZk8lv4ALmEY
jkX5r8lm083gcx4h2HNXHU/uJTsOMp/8bqDZt6zuWz8LwrBCXdNkoyWVCNyRmX7I
EzQeAjN0x1Zuz25h3uUoRCz0SqCd7HRmQSJtI64kMOwuB4VR+EoUpazoce65jHeP
G4jSlvst2GBq/4H3ur/7LjKRYObCpthwXfHOGumFvGkpuEq4V7r6+f6xJ6wUoA2n
y/aBuJ55ac+dsS7PDYcMjgYTkr8R+alTO2Yh97yrarVQO5Ki8W6EmnpNrBrg1B+y
3T2sYMwE2YhSYji7dQCNv5Co00vEDy+FwyykA03bKAQ4cKgGgvoNkXuqMpU6y3tA
gdHli5aRjvdzLhaoXZbA6726v2iNzPEYMtjoi4exLfn4dHC6pLzylVAtoAaxsZXC
mVjFNgfFDWFJp4YEwabLacVMb6RMf+JJ7HRUd0/OZuGL6NUa98Uw/rNqHFc5ka79
YWISnj71pJJXeD979HEoAihE8BqAfWpmkjvpHQgn0yzGvWE4ZFT+K0J6jzkD5UXE
ln7YItpVW9YGXmD7dMyvvRHcdt0BMlJwlHAewt9eTouxM8rIYxZrItzmYIvE2fUP
57tMQzYzPVKl5Bq9bTysfPa82M7FQX2WybAwXzvHHwBdWdcR7JP2EAfykPaNgYFC
A26+GSCHBT5NapmHvWvJksRMTz421oET3tkJMauuwEyY7IaYLhqpzo1XDHooQ88k
TlQx73gSy1MTVIwAAaregclp8GTapDWQDPXKQBG/9GPrDWEaYsz/iLhUbDN+o1Zq
mFNVldT/J5DbJnVcBRTSAnRm5YVj9p6kr+s8xnLKSa6qwv76s5yDNzzaiXZhNDRO
ygb/7UqPqPtkv12i2H4mMsPMfQmDGghCO70JbLfuLALpZn26l2mJWxvfhVKBy+Po
cfO6F/eAZdObaoJwogFJ7DPqYhb0M2tGdoDR1mgzdqOeCXDrQOcP1DOKel3TmJCH
wsKBFVcLyMlsYKH6oZN/ReN9ufc4XLnXpnuc+J0GSGiSlq0LHn7dD4P6FqzoJURi
44TeE1lhW080PTOBu/Q4cbKZcHon8L2yst5klx6nVtb3ywJ1l1URgd4M4UXwUke0
d0k6XxTTirFP77eQuj+zHCH5ez8wIWHyyDkguPEO8n66Gzuopmwl2QmoGYJdMC++
tCh5uxcGjM3zalFp+4UU0SXvXgPYs3sZVKOpWrMLSwBltc7zh4o2YdOxT6QQcWZ5
5r0JhGiYgpYpZ97Lq1MuF314YR7X6YNChOwIbCRTBH+ohLfPZo4TjRLTBoouRjyg
/fcpDw/f1VpTS2elEiHO/5byIJuIsvUUM69v3WSQl3lEsWdF8rOMQDWGUKq8vwRJ
lTfHzOKtzmV/RTRjxKT6mc0H5lLyEelGiXCDfhQMHEFNyyPolWqo9piIdsUGY9tQ
rHkizebEozw78AZ35R1EuobrWqLZNH9yb5ZepB6duF8Ogn1ds9qvR0cyXwORA7iJ
JdGJ/E+Y2cx5skVWalhc3sUZQ1XxBqbstHeFW7a54pAirYrnQc0nH4mOo7tHN8RI
0Ea1QGemvN15YNki1uU4/m7s1j56jGxnN1fckxPlo0eTENY6h+5Zuiv2JMX4NUgj
LWwqO1ncEDub5juVrWURYnMANTaj2LL5umV1cpZ8uUgw8qJoBknc168ozXNC1z1+
sN9ab4E70SnFx2O7tdSMDE8JMQK80uDMTClnOfRA6WXIIiqDo+o8a1LCEp3mw1Cn
K71oqhjuDuvrMZI0pm+mfDtps1Tp8CLZ+bCrRFJ0DGCDTMx11QByxC4kocCElPdS
lNlsyYi3nm2BAiLUEEYmoqAqaQUOYQ/OmwyCODrVQE0/TmyJ1R2D5oB64Al4M8cs
/+MVa+IcAcK0FDZl6HmzmwfcbBYyKHlKQF121fPp40P1jgWux2ShzJkiF9z/0AP0
WZTmDZnfJ9vLIV0gwc7t0MgmD3thwb80CmGSp4egRmxHW0I/Ci0rWW1g8ggWRt08
Gb55Eb/1/PZ5EZBpy5GfvBMuFM3qls779Ptrhhq3LNkxIV1/IDxfYplVOwOjW2RH
dpC85CSWNz/qIm3bT8tibkchTkADHWFTd4DwTFgPj/p8gOs1Fu2p08RIc8xPiSf4
2VJF/V3ri17d9ZOh1RShapwjyBtzsDhrN0Oxo6CCIWQ/tVFi4JnBDKh8QjXnuo2W
/Oa+8R2C7yNMP/qSdVcjZ1i3TFU39KUzJhUUDCjTt8JHDiVfnVS6wnwE+2XOKoig
AAydT85obgobJlNxk+Ldrx1QD3m6akGloUiCtH9Ms4rKyq0d/SeUCxfx6O7tkk6O
JI++xxTY+CnGLCQM7/HwhzYWCzp3df4+3B0ZWKYxlRtUO2wWq9s2V5L7iO9oUAlW
DSjvptJ6znX/3kDARt7MS4KApRrKnQTZVN2AjC2Dz8AR1tp5tY4PQhPDTbj8YqbT
pmcHYorJCsQ93t1xphTSDV6fskTAnrtmBV1IbjPqRtziHcNvbwMfYy4GE+K3BH0h
YDaA9M/01VFiyl7HJu3Xwr0n4R7cp0NP+5c/XzQmsZ1U5MAwIsTqTFvbRljGcFkq
spP90X9Ox+cNB9oE9qTUyRu+nWXFWRcM0oOlURxOMbJEB5frM/5ylAryGIMJn2LL
ShOvGGscN0f48YPCs8fcZgI+jpwHN1iEuGqfjMO4amdHusiIOShlqqtMOKbkT8jp
0AKI6vDUpNRfjpdXf7TD+Ovv0JGxXwn+snpN3eyEMLCwWf8lktMuUzqe9uPCf5Th
P3k0DJxREMlOGMlvIBV06Ajc7SLnvZCL9jXd+VeJ/dS1r/AGsfyiaVK8jpq3EdQX
BmT2P1UJqK01TDY9RG7E/Q3LVDrq8xXAF7VZpldnUJ1zz8HOutE9GcJTdyUT1hh8
yoFQXoJP2SYHb0zCtxj3p/6Gkr4RlJDaBBwXESDwKPrUjIMeNzjrgA0wn9RxAzzc
HfA16kt0FOSW/jCYmOIgQ5ya0QzXzhNoqjWC89qS4wl0QHhLhk+SBFuGILbMUPdJ
PbqA3v0ACESe+ceJQYypoBqtpdB7TrYgqDab8UKosLNQIu5FnN1hLvkTICN3rail
4TShVdL34ucEqH8xDLGdBYitFT31pQmfT1X9zOxGTvlkFxWxIA/4uYwPoo2L9cuX
G8fFs6JoL+731zhC0EdwHwIzkcGBIIMqd0BiE0oq0CqG4vIFceJdbfNAtpWotbgZ
odmV5yoe+5SBnEklpTNhztMZDLnmlqCqJx910OkTIncDc0WhrKVqlF2v0FCGC2DD
EVmfR5ZEbP2QsNsDbXpAYsdV0MMdIckyDKJCgoE/LdLryiN1+6zAupOIkoMXiLJp
vXm9kv4L2vRQgaWvvt2KyiFVJzv7HeuiX03UfFJlrnJK/+I8J6H4knlVCvWu7MXf
M49w+LVrO8/sXuXrdBtCMUBE69xbbXt32QVBjBjQ2FgbNzx+fK55+a0JRq1jIa3t
C/Ewid+2hRUjLHFUtKj2v4MwevkEF2CSIVWPpkrEu9bFLCG1XEyOxPlEwpmew1F3
/Z4r4NQd+/QQGcbReJoZ7wQpckvhwYpZOZJGWOgTJQ19Zp7TPcofwTG9pDZwOT8y
BaNaxiLjpAs3Kv62Gt5KA0tL5KsBrO+A8p7OFHztktwKiODg5DuQCY0qhHXbo4zn
LPvQkTYX0oywlVB7FIfm6G16lyo2QzrgEtOOSz6nIEuauVRjL5b11MZnDUXfagmG
62AwUigi/rH7jRdW08tTgJdb4aiezve0JFYSlqhesBbuzODw7kYOxCpAB/YSP62z
2lw3bjGjoOpSQyKOScMeF672NB96KeMOzRcdleV2HYFH0YqD4VW1tKhfvenpcwmF
kIpTLMLrSOARfOqXDTb7adG34CmyqVuI/dZTKnAA7IYX3zHCgDrSx/OOaODS137I
SIWFd2C7RMhPuy7r/41GTMXlJnleme1u7NSZyka8DhuofMzhbTRCjXD8C+xcUG0K
8eCID2iwYh1zmPpRIVNUyunZqh1L1gyBWCKbhChg8eXvkRm5o3U7Y9lNrfoDREAa
oON6FjmnMTIfezTEqc1fgtKAcKAY4AKO/2oEJKDuFGmsEzlSJDmRC/Y/qv2yzeEo
FycgCiG4UD8oHIMUSuKvaem/ldlhH1EzBD2wJxTDC6BhRNoFzBbs05mHjg0Sfz17
axU6JK7u+LN1e5E3s7zAeKFdM9YX4l1sdTu440rfvy9gV7GSPqk2PEVDWfvlIO8b
bOVbMONAqvxunppyWmDDdkbiPGq8g6Wdgccme9zXwQyhJrk5lKtsVMSU2++bPg7C
FI997UOCZfnQUf6Zb+6rtqvkudwG++PGsZoLWB9t6y0B+i9aobWTlFLyfAnz7VEB
GKzOKGCXATiYvXqhunJz9gquOxrE0wpckhBQzgkhBcxlqnOCCSp2zrpiEjhzO/aS
lQx6P76F3YVijEWwWC/V2r07C4R2eFzxbFpU+x+GBzfogqiwbKcN9zVby4dpQnZh
WHOpJN/WpkGkCPA7WqP6U7EC7Vzu08v7zyKDYLLomdkv4hnDXiZ19QWT4nPK0kW9
FS6HDBPncm+yXDuB5u37HotM4MT1U0RripcpJclXuYI=
`pragma protect end_protected
