��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�2�2�*����Jdf�g�4�c�/����RR�
q����(]<��
�>��B]��ɚʒ��:
��#}�h.��4�.��ӆ�Q�y��;+�����-T��Ҵ��>3��ls��ŧ�l��j>ߺ�ۛ�~jz�g�F�����=�}nqR�.R�B)���Y�9w���}�F3&��2�0ZCkA�뀭����S�v�e�	xW��.iD�؟܀XI���wc��z���@x��0ku*�7hĖ�á��a��|V`W�&Ȃ���'�a1�;���O-� �+]kR"�;�GY!�T{�5,�' k�-�:�;��^�,�^��R�;��%.e�^}/�Qz��=�����`�Ne>z�XeYu�<ڬK�24	:v�M]izH˛SJY=�$wS�枷�_IQIZ%�|�LKR4��JB&����f��u�u[Et��$�����
��� �� u}�}k�(3j��f{�a'i��'��4!�*a�'�������=<�_�]����C�a����p��c�U$��6�G���O4�O���@�(d��W����:��z*�7�o�櫻'H�5�I?���+�ۜ|�;d�x;�U� ��JoɦhV���c��sW���\�dPd�r�S8�ڭ�4�a�&��ۀo���0��T$���)�p��)Ǖ�1�$�3#��s��Wr\j��A�C�o��=J���@���������h�-[�{- Ԅ��p ���ȭ�Z���E`;���Վ�Q��1�.?PM�4+^{����WZ�J�_=�m���(���,�<d[/�����=�j`��E�����svT8���7��o�����~Մ�l~�dV@D��{.���߉�"��q+��l.��_�J|���S�E�P�P�����!M(�S'D����j�*PN_�ǩj��9���&eNf��ľ�o�=�߱GX�kg�ݸ��q�1׈�p��&�WbA��ݼ�@F�E�S�:G]$؝�\M�[z1�B��V	^��`�s00��	�cA�9��|,�D�wiV�����(�����-��|�^`H-�X�����F�1~�"pQ�q�/nO���ޥ	�^]ܚbZ���AgTFu�#��
�0�n�L�YN3���/�!�Q{Q�U�D�ܟ6�q]v,w��RH��� ��LP���n�0 �.��m�e�k�ă5�i�!]����B�{p���j��$���BE��5��4+�GAD'cpF5hV�\Z,m�)y�?��,��Lo8.>\��S1t*;*���DC�=�ݸ�U��HM�����g��-My0	t�?�"���j��q�֏�!�gU"#��<ȄbQk�u(Bp��cm�H�O�+� A�tl;;�}�dB�=M�L-l{|�Q\�ɠ\�OY�ٚ%~k��ǖ�!�:Ǡ���w��$������C����r��x�;�oU��>��ܿX���n�}x�B��s��ekMS��e��
�|����y��S�vC��X�L�R��>�۫����I
�����g���@�f�u*-��!��JWL�kzU�{��O�=ܠA�/ڤ�IJ%�����/��[���/�.�}����L
�w���~�ppQf���~[57�"0R�T�� �K�h�X��ۄ�
=�gء6ND�)x.C���"��%�����pyٺ^���zRT��TYH��~�������M�S�[���P�2�J�id9/�^Zj~>#�Bq�r��B:N�SI=��i�:��2���Q�3(��7h���s��FT�2m̾P�{��+f ����t`GK��3�<ɰ$�81�~�a	�59��Ť���;���N��ﷴ�0�/8�&	k���:�$��`�Y �vys~k_�Y˘�hn��k#���\�@�Z�&�^���t�-�����}a���A���k�yD�lk��^}��.Q!�[�3���c媻��� ���?�J�"loضh�e)f(
�ԧ8�'9���7N$�బ����;���3�P�~j,g���� fvG@@t��i���\�Y0����O����|�e�&�_8%��b�a�%��F-O��r�i��XB�O�	 �ڝ�g�3oeY�s��g��R�n���x�t�Z�� B���+4%Xb��i5uE�b�Y�T1��JL��:�5�Ҕ�~�Ql^�\�t%�3��J��p�篖l��N�Ht!�	<ł��׫�0/�q79���P�):�*�N��59�m3l���jq�ŵOL��72�u���y�M��V�AiɈ�H���3�� Y�TJβ`��1�x����d˧���H�A�uI��u�LU��M�ղ����]�@�F���9D�տ���K�����j~x��V�@�,7�`t=\RzZe�P�u@J=���W�>)�
"�+�Қ���w��e8O'�����2����e�?z(���oB��KUYO�t�J'6�|h����P<�/��r2"���{��߂�G�����L���1�p��ֵ�}���j{���[$�'s�i���g�)j�"���ja'�س��3~A{�s�e�h���W2�GW/�G�v�A���^P�T��r�J�D�:�Ȃ2v&�W��J6�Sw���&��6��.��P�΄ݟTR��/��}�t�$6⣼�w�)^L������WԮ�@wt=�4�͌p{��b8�y�������= L�z8r鲹�����d���%m)�#O2I�;���!u`�Z!�	�I���,��"r��f_I%0N��K�h�UJl�':�&Ȩ=y�;˅4���ٜ~΅&�� �ǅ��]_y�w�y7Ata��
��x���x]����9߳���D^�6��O��2zj�g�+BIqwex+�q�<x{���xk����}c�,��"轫pL��+�o����Zby��)=��
���'vtE�_�"����	������`k�,��yh�E