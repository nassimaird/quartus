��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E��,�׮ـ�-�(,����9��_�8W_f��U�"�g+f��'
��o�/��^!�ݬs�}��"ޝ��ٝy�B����i��%!���UA���Q�� A��a���u��5��+�-��b���0�+�6F1�!;Q��_��Um���z:���ZVK���\�z�{�fF��"5+{a����m
ß@ԑM9�4}���^zT�4t�"Bl�׮{��ѠF{��A<��))��\FM�:��d]yFdNgTz�%Nسn��:C�g�����a�c����m�/���I�o��ՕW�V�󅴈��[	4;>�c��N�K ���!���PfD�Ɗ"�H<i��v<�4����VX���,����V�oÿ�q.��7	�Bݙ��K�4�Vm�H���U������81�=x�o%.���|�7!6q��I�U��^-w�KM��}/}���f�L\We��f�%t��Y��q�4�B����~��~pݧ��ݷ.�8��	�Mm��!Q`�pT���<_��D��o��x_dT՟�1�|�>�gΙ���f92��/N!ە��?r�W/t�Vl�����7�hr��V���=� ��7�Y')�\�/z�V!�D���Х�Yx0&������� b��s��k��冘ȡf[��^�ox���W/u�\��\d"���,��æz_� 7N	�g��I����E��<��}D߫��N�Boe�jeG��ܨĹΕ�K=���R1�
W��sX�TSB�C��P��񷍦�%���)�c]&ٜ�]�YϱH�
�]c���ǎq'̏q;�&���G�r��J��[������I�(���Ŷ&�NA�6�{T�rB*��`tV)����z>����Z�칛Fel���,,���
��E��&H�4��j(�-��da���-1;Ĵ��1�)��Qߟ&G��R��ƎࢁH�c� #���q���d������#���sP-�������w���h�Rݭ�O�s�\6�s����̕ d��f_<�,eTΆV��
��^{��DH:rC��L@蹘���d�KE<�_E.ՠ�U�Y�|n�!�<0y3���5#�mT�?���� r�X�!��G�@0���wa�9�F��3{P���(˱�i^����L/�{��!ڙӰ����C��7���	l:��Ǉ���/ꗓK)S�^�F1b9�+{v�W�Wq�����`�J�0�C�g;�ܿ���ji�&�QZM^�Վt�h`��f��=������w��)�� �J�z�{+"��Ӵ��hK+��I����:B́��m����I1�9R������5u��Y'~��!2�M���w��>-	}�mG-ມ_z� }��o�n�f�//d�RL��jې���u_�R3�l ����wS��P��P�H.&���Q躰�qw�ﰨay�\,�A&�h�H+?Tns��`�ښ�X�18<~�*&`[!�[࢞��*,l�'HhXP ���ƒ�nΞ�fl��^��ݴ�@�ҟ�A����ta�p�Qp�|���� �]]6 ��L��T5�tn/��\�K�8iw���&��1٨�DoȘ��x
.{NZ��oo����*B�ɫ}ء���j �+z��c��c
���L+uɅ{șe%�P)��A~W":v�S���]�!npA���1���>^�mm�S�R��1>7�.�2 ����Y��J��S����׻_Q:��X߅�v�n� ����Mo��� 7BC�Gf�Szc��?Ղ)�L�CC�`�Ӭ�:Z�:B�$#��A�s<qތ`c���_͎�>3iͭ�������6G9��Mq��2�(�Y��y�$�;-�"���iWd� �F+0�̇&|rc�=����SoĪ��y��\V��%��#*�_�(�gz��(t�g�'�UE�}_�!LJG≳��7���y	}/��4�=���~T�G��o���;��]إXdab��H9Y3���U�c�'&B��2W<_�}�L��(���ó9�5ޏ��'t��qn�ٛ��~ �!V�	��e{f�?�۷zU�c�V����;���֥R}�2���賝���m3d�N��N{=B)��B�덏I.Wl��׃��T��rU� ��P��X@��� C�%XL]+c�rrW��������8���	�H�O �y���P:r/�6!Xrg)RW��*�B�rϽ���'�/ʁ/���#E�L��O/}B5:���ۈg>S��SҐs^�!%�RTy��-�ݵ��8��],��n��tIbiuƬ0�/��q/,���y)�wB�l�Qr��b�2�(����a��0�����1�#���B��� �u�$V��4�Q%��T�a{IWa�oD��L��/�}�~���3S�p�i�O��G���Q���a '+�,0�Xff�Ĺ�o�)Bg73��r`�C3щã�g쯾˯/*#�v�
U�k d��3#qFI�]d��0���1'8F*��$f ��"�c�b�'C*��+t��";����aG�i�O��;��n������\:�j�/�/�qo�dUKU�G��j?�t���u�����2Z��+���la�
���y�<M��Z(ݡ�BѲ�KR(#=P�V��$�,��?�%�y�����]p�28B���-��@�W������bG�^'Pyg����T�m`BH섫��B8���h9�+vբ����|F�$�2>�c�Xj�ԇ�`t>m�ֈbF)��0���OL~��xNI���̯J���v���#�6^U�����x�l���7�Y�h�%� vd
��(��o�#*�?�:��3��5�ҹ����Qg�b�|�,��!��[��4��������Q�m\[�XK�l�V��(�� ��a��� ��ȏV0��I
K�� ���H`���<\��?���^��J!V�]>�Dx�|�!���g}��X����Mg�]�)�+���+V����٣8���֊�7�*��ode���	tWm'���P�����G}�r�'m7UZ~���t�X�N��8K!��栫�]��r셐o�щm�8��A��%�y�`D�+]"3���=�ZsG��Ju��0�{r��t�� _iCӄ�*���'���@�
mD,���s`%s��]��)V=ymW�q;4�ʧ�lT����p�i� ��5�Ir��<';���wu�N7V���PP��R����4\�y�dz?��l;6V�	����Z���Ȃ�Ϝ+tY�'A�+�i����1#L�_�r����(V""ov��.��`_g�	��a��jQ�t���\����Yh2S�_ź�8�&�Q�cD�����֩��n��`���/�NLu;h��G�k�IE�!�oF^<Zq{ ;ђ��ߊ�uy�����?J��q�s4�����r&��F�긠ʷU���m[�[� '��o�� �����$p�>ٟ� ��\]������ɤ�Q_L�v\�� `dڒ|��w4�dC[��y2����-��n���sm{RqB�Uș�X7���~"4��h�.�=�`b�y��j��p^���#Zg)��t��P�ר����7ɋh��)�.��Wr1��ۻ��Y�*U��kB�q"Ӓ����j5�.��-�Г�XeW\l>5��U�_I�̵�yd�k��n���5��*6T� ��}�E�TJ�U�`W��
��܅��א�ҎT#�Z��K�`T�v:��U n���?�g*�.�H;��L���+��n�`��Z��:�1�(�����`�3����ma�,�	j~Q8�-�d���}����1nme���E,�t~�o���X��W#R(�ԼKP�b�����פ,��>V3�N0W�0��G�^JH��@������*�pe4�^]H��:K">�=�7NɗώC������q��xO��IY!��a=��)4�4�O�<.�M��K���J)�������	!g�0~�
�5<tSkQ%V��4���:���	�D͈>�b����ϋ��K��* ��(C�uW;߰�+e������m��U�4�I�>r�0�m�M�( �/��cO��@��8wX]�RJ��]		�֊��Y�]�7�[1S�U�$��zAaCKCd���`�W�c��M���)��ZE�cJ��؞u}��9����݃dM:�ٌ�B)y=`0�21�Cшj�Q�r܍��(�8��"�-��	c�it��I>5f�����+�&TXR�~y�\����E���V��(�N���S�oD+��.7k*�w�xB�����k�gr�3
�@O�Bw�y`���L��7�v�aܓ:��X45�d9�xP�UV��_bR]{��Z�(�Y$�`Zt��xe�7({ ��>o<,	7��Qf+��n+Y+I�я�TjRj�lނ��h����M_3h�=����G��_�y�u/Ҵ�pR���t�qkB^%�¸p�2A�<o���~�~����9Y�z��]����p)pTMӮ�6ڐin�0�i=��dҕJ@v֤��Π9�~?�����7�`���a]E�;7�-.z��O&]Ń�g'ɠ,J*j�+|�dԛ?���hS�hZǹ�]�������xUL��ܒ��A?6Z�8���6���7�#&T�C��=!H��?����Qtꙩ�Z�I-ɳ�&�آ0���.t�Pm�,Ђ�g�/o\U<麄~2�oP�50# �
��2v��,�/����t�H��U�?f�M��s٧��v�LI̚��u6�Z<O��H=M�|f\hu�[����Mjt[y������!)>�y�����8�]o�sW�k,�DѠ�BT������^(��f\���I�T��Y��kQ�x� ���,�i��[-k$