`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MQe7vD9RzWQ/d8sScZnX1yK3Ryg7zXuPOSLiYnZGIWQ4rA0gT6EQMnxXc6zQefeF
0J1iD+64TCBIzKYmmsaq2XmLYN1cU3t8rBxWrdLEfrfFbb1nw5Nfr/EFG6sHdNCx
WNibzf5H25J+aHBIeeGpzJrAdLxCaQSvutvUAs/qh7w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 144992)
ZYgxdEGW/EpcHRhnXcyFpnxESLK7/8GGo0oYdpSkrp0eKazIgx1LUR+Bfc6wgivt
nibYeoGY0hQtRuUbvA6kvq80fnGRvZ4Sj8zcpaE0melILaFKd9cRxDBq4UYGfY+d
quiYq1gukniEf2qfNijWuuogVx9vcEsSrHmTAxj0dmnptt4SDtyqKkLHz/GCT5y+
Wi3Wb83OywBzQCAOSPFiKnv1C2BKaQQbR80Xs9XD3gwr0v+y2WGGdVgJ5ZZiiYtG
qkTAw/ltwbZu/pN4/ubWsO+TbjevFRIr+I2hRFJaQTtMPI10pvYCcoZR/kO8a4TX
/Vr8xovL+zbutlOkQRs7As2J2kmZ1uhKD+BJdomuBGoX3SkHwPbkPep2+OX+WAoX
nKmsQA+Y7A1pC435IUdt3rDJ9XiLvVW9Fr+R1a3q+Q+wjo3BN6T9lRqu+y/Tn6t4
cYvnEppt3u9Fvbpdb580sxO4ifOXuz4o/CXWzU1H1ICltxIEGisJSTfOdur+g/DU
YMq0hcevMVS3+qgdL+IsDVpxXAc8qooeIn1jGb/0+61SqNu3lrlELNhv91X7ecLK
5bLm3JXttrmKEf6ejhnjVALzUkPfhBWCwQeGfWj6S610cIkmgArmj9Y2yYjojjhm
yXTv2P7nyGDK86XRZlK7+oEJXsWmd3Ku0/PEPuYEj8bbjP/yNxtqk73FKtFTLvxy
+Qi2fL6/bI+c3QmqQ7pPKrDT35CTtFB3THwBYW7Db0k8vq2i0LG69gFinjuP4VcW
nTWLm94Ms8/Z0iLLWHzDIQhAgcS1DyZ0zaRlkUnnWtX/vD9AUurf3HGZBaXS7gtU
yr4GxCau/RRoqKdxic7Ji8z4ya+L2F8uDJu6dTSEV6TWfBJvBCxZHd9Fzoz7hbX3
qgsxlLWdAxOTE0JGq0UXJmIehcY9WUHosHgva+w/ivmq7AztG6kkgEiJLlM46pqo
eVz/Y8+udmu1Dfn8qKJetXuufpTztw7i2SONU7DOIXdQHO7VXNucx7Vaz0BkhTSV
vJSZ7apFgYz7mPToZ55puHo7Gn6mjUpHXWXVaqgc1+qtlYQAkl1JIvRJem0IAeHb
Ek5ugfizhZLsEXLE0LfXf79NVpMnlKQ6B2/cZPpE2z3NwThg7zbjnVGQCl+Rlh75
21zsaSzPsqmfTV6NhxY1XNy7pgBuBrR4XCNijBKPoYysQ6SPkM1k773+7Ub7AgfG
BvuLNqjMfO5DxfZoxf58nOItG/k6U1mNwpKQckEmf3s6c4TqDfaVE/SXXsqrBwIc
f5MglV+QDOCBBJCNjpz3GrRXsW7z5RJBNrNoaQJVZVhQIkuQnMrPjwxdrNoHDd8K
88i6D+lNOMgsmjSARVIMOx+rnP99ni2F+zZxDK9+uwTz+/fkNwDKLF3B9Gk+TJj9
B+jeR0XLX0rdHHL4J5bFfqNFew2idoAcNNRetvJV6EIBiPR+wPx7nty8X0QNQ9kr
HRMFHn1d/gsWTgBiqP0hkicZg2Tt9KO+lpPh8aVVKFyx9XyZvT/S4iTvw6BrrkTH
1+vMCF5pDsqQmjFZWfrJTwGYZ2Pkii0P0sM7iJsd+YNnwrykX5IH4IzTAZq1Ay6m
yNmlEAdXQASDoAqPHCYPIQi6ufIuYtSPsyUf/Rm64niwiPOWoWmUSxDoV7WTppNE
qR2LJtGpVJrXXPVdMJT0wD57SO++PWi3XxfBiufE7G4esLabvOnCky5XR3z3MLaT
4v8AR81WQlIekpM240+HaNLiUSd1TC4Nq6fSLtQCHdwOLb5CdwPGNrOrP3aTRWAi
wYfemFDGld2/mME0DGlRH2MKL+bGk2ARw2WBFm61gYpIEBZAudATTJfi3yaqvpEN
iwKAzioh3CC7yLDuQuoxX0iktTL8R+SL47toF418ukfqAyfsqjIEFyJ1vpzZU76W
wXjQoaB+WNrJYaMZ7sItE71k9a69fK/Vxy/BqIt4wWb2raGXOLEBOGphwWT0JU2v
xhAbp1Kolcyuo0m2uH0WTjkT+tjxrf5rmenbmGZ4mpe3tfP6A+xezXyhYq5q/IxW
UQOhZT3nNVVwOi1nC8UXscJP0bRkHugKdpUu/ERLeUnDc4sHL0x4R+zwwj4QojQw
bgzX7zTNeCnZkkCiPu5A4bzKUTRu5kPzdvLD8vmToBK8w6Wx0dW8NeF5V7Nv9AV8
HJs7TohjwgOZHig81vKE/HSU6ooX5cuuPZuYzoifmHz2TV4y8WQrurcjyIPMYwyQ
gGo06e3kB97sddC2i6IKcALDaxS1aJtyxkJgrWe4kl7A9vw0H6e9mSWZeRKDXqb7
PW8ueO3R1Q/IhLx5sKpVFRGKP5wfoaFj6SzdnuiAledd2WYNE1JcyKKpRChLQFuz
jP7Orl3w5rwwk3kJnhhCVAD8Bw2WW2+jb6SbywHq8jNGnBf+T/JYnD+U8iDvsJPE
ImnVRaQDq1DftSHxOC8FBIszq6FgOmKtoOCX/mh8ZPVYVsgpOJIOzgsE68jiYfWe
2ZpWF7x9V2DPMRryuWGA8r6LIoFVxD1rZvyh9A9V3zDjzLjlXCjA+s8BUbyPrtuz
oisM1wE1h48oWrgSxHtKv0OHuMhbTy6SaN3PrXq8b5LIo9Ss2BRHE2s/SXvL0xYJ
TDthk2Sm60oVglgTgl+GxYQuwu078aeIvnL7HqiBSkZs3K6KUmAgk63L7tslox4L
PPtlUKRgp7jUcWH53L76crTOW/87oCPAXETGFwAQwVIEMyDg011jOKMMIuVa5mJp
0qC1APt5CdnEtU5mQpyZZ7V5Ud86DLQFFf76/TSizbFoASRv9ekwD93/J1J023ek
sxkKQmJjZSHPs3yPi0ZoHWyaGzvr+mdJytzmJRtTIh5fxwrT2fUXAfSwI/buhJuu
vZxJT7wGdsOpWrJBd2T8eucSQUOvx+ovfenL2YFv198I2hPWOangF+kTrox0wWNR
SD4Y9TW7A0ib4i7AxtRDsQxs16YQ7l1IN7ITlqZXyG+xctUPq9DKmn2jxbRPq42y
Yrcl0aoepTNv8ypG9S439D6PkFAGjF9G5YHrRnOwrxZyazVSvfrqamk0PdOEQC1D
ygerY7HOccZHcLaaVWUxlCAkQ9REuL13/pDS2oJe2BqdGjXt71ObtuW21TUksYDq
/bMybvCzzS3uBkqiQ4u+1aPVKlRA5OMAHTEOYC6TLcXGcC4Jd9/XtPPDc0pdwCTz
ViG9ezwzC5NwV21h+DCC9izQlLcTSLvIyqjw8GmQtrSb5XR/y6XowudIDDaMz1fN
QBeCBJFaXxpJRsGOVwuZGlwAwqhJdN796X4rKmWfKurCNhWR/jfuekn075Yj/Hw6
9w9maanjYnwj4J/INxHasH5it/ic6EY39/WG8t4Rx3Ff8UbIaa9baSDcSHhADYXq
6Dg4fAvutrsmFICMa55T1xTT0vqlTTFTMaYpA0I4gW6/PrtpzCpRKKVXwJV5R6Tq
Azw1xSdf/xCrwnt3IaivfvpRQHUf0xl4ibE/Jhq0QEDXLaY+tWSSIcy1ZBJw3o4r
KH3woqK8+rARMqCtXiURaMa0OmoyOqvvF2EzGlUrlWNg02XYu/gV58+EcnT1B/gU
Xst/tZFOVk443a/YzSu6F/KWgDuoSeZkBYh/3b+U4ITwCQeEhtb1EPcUPO8iC1Rq
lZ6NkRT/Pr0bLBe7asOWeGXpnHrqPDqnrHTg3/TVPiETtkZahQ3jMT7nowXcLlg7
VuMpfYUlBsZwjEBbGn8vtTSmkv4zCQvSKSAOTseped2lG3IXoHwh87ji+0VRVLhw
lu9C/MtFDcaW5aEhd6HmbMEFL38i5RBqYkgg5nYycdkxBDiUUg7/XPDc3UKhdhtQ
DLsyV/FNriKHmP1JYVaPM6lKORSvhYhhKRDiONxkFxaetCKfIdVraVAAhp9P54Qv
ftGFVKXJ7ii4JF7tHdKqR1G3oC1PECigDqOoXy9sfmAs+Y5gwKJH2Fo+YWX5ihQx
reP8Z4QmYTbHctFF7HfpBgsIDARIbyOpiJ5o/v9puj63r6utuXNgCTeA2UO7S1RZ
KK3UzvN7kKUUOQqlOEaWuZwFZqNw0E4nSKdvx7iuS4KcZo5bCDoggfPzXbh3xaS8
hTKBhD3ndeK9twEfi/2AU+v1Ldit9q0FGsizABjMkpNTATuSrciZEk2PtCu/08WT
gIuLbESbWTHB/hdMSDij5nCRaXuTgbKdA5h/aQO1lM0IDLgY90ntzpDX70Jur+fw
ddDHtQ/DbzyH9bcvwEie2OpER48a9voDxD1rpyCeX9ZWMKVaYIpl0uPcuhdSG4lu
j+Z0WoDSC6LYXjHn6DspG7TLLao8SKYX+priGMQ52zP6adJ7cpACyu5UQBexG5K1
67VCltSnIZoxme7/KWk+a0hxtcebxyCnKZFS5UQicuVdtNNuOjGVg5aNr123Ehm6
GQvgP24HeD1zvLdclJLdLaIOqQNTNcYgfZuEriAezPcBRaMemQy0WHnUfJnOGkoW
Gl9m927MH8fO5OBxtQebY3XEaHWy9izVBbeELxaaOCTbVtSwnzmnJQC84GfBT9j9
Ho69Th+GXmwch5CRTRq2jE7W/SDsYY3ouX75GWZDuHUkXCuSIzmre6MaLPM1LKZC
U0EJPk/qNg3rx1zJPPIOsIQZCghsbUa6wm4kSN7TiVETanjFf0mk3XB9nw9VSX4k
Dl69qzutQfhWRDwoxpuajkhIm0JNHP8sj6zs2MzTrEzgZI157apZJBmsiWqHRD3r
3xXRzftVrgz9D5PCYA15CxvbxSo4ex8dLi/gZw34ypyCeR7iltyoUGXwUzRwnk5o
cP6lgpbBWBDHSSgDEVEpQriVBNQzHzRcMfhpAnze4TCJBfTMzmGtOdTcWyOf4gYU
emKw/9GUDUTPGxR8Wj6EKigm4C68+GF33NmEvErYFHcKgj4QL9SdNeBIAS/tW8+s
0jV7CFLKw/7EApOUo/2VGiuzfBKYVCJ1jC1G2VsDu1AzmaZiRXbvh1xMNCzFrWTK
rU5iPgWLPY58nqewpxZHWt6eEUnafZa2v0A2td9tfPfBprilodcQSXa1Y9nY+0Ri
J17O+4K3rXVe4C64XpLt81c+qMQ5iIPu87DLmW6FmjdCMUAwZ1uIoh0JYCTiPqoZ
hchgzb9hMKhjP5D9W0sijdxBpv1/KKnNxkB6kr1jaa880nbpd57inKBNrglFbCzb
XkPgmqITFapq9CzVVQSR40uzCjMWaMRXpkwm1zjZe7lclDewTjGJjAiTX24P5f1w
PWKQJGRR3Lhw8fOYerUdYAlD6TKLRl87dMFxDdbMEbiijXxSVGBmo3GkSrTnApKk
7SG8mnH8Om4woH7kwqmftO5MDgW3dsSuQObs4u7IznrCDWjxqXSIfpBCla7b3WPI
krOlsUZ4+iM5iKA1BekieMkAGJlDjZz+8pQAPUV+2AUJRL17NV/VAAXdeG3SY95m
bvasphM5EZNZecspP2MUf4J3yfrXrVKVWcuL77QCdQ5dg5+YsNwBTB6Fkhp7MnQC
NZxvdtqj0JM7SFjEh5kepUfMIagWneylznfxB2i9CO7bEVH2cKo0mBtxcKnCviC5
03IGrYjU8eieRs/zfMMZAv6sniq6kbsXwSc7yj+wvUqRGmYlZFJQ3cKkt1L1AycM
RE4KDe8bENAvXjagHBKxkRAMYNwKDU0raFAo8V7o15kA3M0r4xLbgJYZshtCJM2q
Dd18GrSSH4HgV92O3qD76xn4siPCI4fREpXNikF+hs+6o/puL7sTVULmuXE8RTaO
QKe7zEi2JUx6DAoE3e6DCp5PFM6Q3OYe/Cpu68M0bxVTZGqy3p6cZDkxkncOqJfy
J8m3SMw2qnzVUBGK+jcsHzVNInXNH+V+uP+nOi0HHTyKcuff3DG8zDxXWxlTF3dK
zjs+sd60kau9aQh1TRivoL/3axJLCHQiGZHNz4EWvoeQZlqXReKlLFRfqfslLMgX
vGRdH2c8j15sdqDgFiCbHXiAdGJvgBDAfC6YXvAL8bqNrnse/DzPIlxNO9QvtaYQ
NKSZw7hMJLSkBGZLylU6SJeLlqme+Nz+f2sE7ZFw6igES3Fa0VGoEHkXpm/TAm5y
TrSZF1lVUuZzKp3+RAeyYgMLs2rTv+6WKJ7wg2DqfcVL8C+bbotpAxliZp0cCi9r
2pjyyAGwBu1B183gcCGeHYq1fB03xMF1/sAN34jucs3r79KopxpWLDtvk+72p/S1
9SIVxcvwv8xx1pgn+ifccXxk8N59xowtPhZJXMWIRdP1xtT2nNK54gTpBPk9Lxkt
skEDHPpjqgCN6tfIBTkHmix/W2TGi7IMw4zhHN5I8gvP2D0lKfdgmzea49rN5PQ4
mKhLDYlZHlILd2f9uyMWgZH3dBz4cbSxCjkqNoIzLmUouMe5ojCZJ++vwhzQ6kVa
xQU+CyiMsPNxPPZ9SnWKOBh9XXmJ4z1KfY6jr22iaHKzOCMf8FkvGSs6M1ma3NQP
pAgWzFYPo/jCElhKL+uFQiwWrOXprxMe5VcIKo6MOWnAqbqQ5+xZTgAIGamaRU5y
bP9wyFs4W5s/7DOujc7Kt1VY/q/SSqGYgT51NSiuSgq4gmQw4Pn0KOa5NYbvmOy7
noPzx8VpNdAdSsLxFBMrADmLciXgDN/5EPj0Hh/msreUdSgsZ1JLlk6k2OX6s8Iq
ngMUe2PWSNgtVFEsW+v/5jRi3N+fAUblCCscK0OOMW2P0ljh4lRJayNFtxxWmUz4
6dyg+wFsiYEbuuKE7zycNAlnt/BnB0Ro9ijmup0Z+vbnRDLXdyBi+oXRLNA7v6mT
ghQvkjY/llWdMpxys87S+4lW+L1hoPYVm4skl15dDTVPVb5Iojmu65aCcqNqvpVr
Hb4jf3inmiPjC0XQScLu3ZnMXPGEjF3zUDEklffO6kIjidNNqKQLErz+zQeMgrCn
bkOdo/5LRsPmDsCNduBmda2PRlE4fKd5U4G2EeCjyVILGsdyXsBDU7cvpA29Zghk
ckFCG7hfVVxpRG92ClIt/9QnAr5jpSfHfAMhLYDj4ph58JnrX6Sg4UgvKUn6zilx
BfDnaxmMEETrTFwodXjCjnAzUl1V1D5qdaYGybB6bMXMMA+H3qSE1mDTh95y9wql
RsTbZKJ9a3uKHGt0LhpYJREmAPy/5txQZW0etkokITwmUGaRcVg8KPmVU3Aa5FDC
52DFy9/cVgWiW4FOHwcvheH61XTLpkPEBVzygoKT/u+wsAsfgKkFW/RvV0o9DWr0
4eOMiwlRqLVazcSbATMLA4yyDU4UuhgFz8bSqxMTyjop95t35sDABvbEDYiZXJHh
gQsFxClLcwwvjK7uEqo5RZOCL7PBBucHBXZe2zJjnFoiFSXJEdB+JOZRI5U8b0o6
DANk300P4wdXjFLi8+Evo7XQOPMNXW+JKJEEIcMxlQctyiPgNqmF/rDYAiKtsv3P
f9I4DSafrTom/CHPFdzGIml1NQbRUzZ2gzqbiBInbd59L8S4i7WS/EPxA6Cj+2rp
shU/AAPI3I0+B6xq0S92/wY1xaTEzaieu3f60/tmKMUpnt+BRR6XaV6q8wwmqxMD
+FSqOUbslaBu6p1bnV2IzcwBl12mlTtJaNYjpj+N3Sf33vF/JZdrwqr7wH/9vrAS
rQ4OtloAVORJD55SRksIp9A1d9M8lsDw/BdsMLI6jnGVX7Aahes4ZP3xZlrLFyVn
eM3b7kJKauQlzFJY3EABZBZZNV822vt1++EajCqbWnkByyugMDOE2wneEcnDltG+
WM0H4MJSW5QymsJI1ShA/7Ywz7gYl9sI9JQBTgxapx51J54GKo4sf5Dy3QddBVBf
5b4oL1nBf1moxKIcW87f9ogQgB1hhj6TyFaQzc5+TV+Y3oN72JrdY+m6FpI6FimJ
ajwCUqEKaR9MC4tkmlPK9idbR9vfDgEFkcF6y4RO3gat6J9KV1KA4F/A2lFb00Sf
1vlkBIuBAa3yB1O3Z+DVNzRluNxamIV5VNWiTlUDA4JaO7imAjF89eku1X/8MQZm
tPSbRFkr7bVk1ACJ73unxP+bOfpyutplHFaWBjyrSNRXqORJZjLnYAMgOwRERyfw
O+D/mWNIJzrqepbvSCDmbHxFkpN2gOgz7AkpShpYFUeHE5pEh1h/bdIyfadRu9gv
pahKt/VgzgiJ0Vh4+CIyWJw70jsf/+pDXZSi/a8xVWxdeZbW2qOFY4KdbIbXaK+6
oOU41g7PAUBl2q8COpyMHkEqp+M8jKzEMRkybN78f0TMtn/QWjqrd1GTe5+kze9F
tyLziOMaZmOZ+PoABZg9BMkiGEh+qXfEFDIpMfMUVPx7tTDdNu3gIUjWLEbW2352
3JhHJryDkpRkpbXCRKgPhVyBJNqUSXqtX7YzQkncI9I1pM0hFhv2ii4HLYWtMXIU
/JG0YvFft4uLicNgM9nqxm+dTQ4EN2xWkvLYYA1grSu3n0v4dcPxy0RNoXEodWOU
1jVfXbLvWOL+c4IvFUuV9cjzpFVtczUHkS2xA+LIcatdr4gavxhKbNKtC5yrkf3U
0/mTP+IoXj76yfb+zRb4ZOcgcgWBYe/9sHNmx0gRN7jWHw1KWlpk+mVxpgCJUbhM
kScKGdU8iVjF38Q1YeTHe6Bt5KH0x4Zxb/h/89depheGNO7iFkzHDHR1lmFbAHy+
BWi84tHQEW+CmyzdWXIOgyEIy90gK0VtH5YmbItB5Zilw/Pl+mqSB8mJTpW4B9uq
FU7eIV2qYf0G+Hul4FbxxCVxH66AlfuhYhg9I5fbzdzeMWyvy34cff3tQFi/PM7w
aqa7IarZxhDXcPyBisQJJBMzUJPx4ZhPekCY0xIoGJwVq+bTQ3UCw8wPUHjrMBha
QPus8t0aVa0OhQTudzVaXMsZNICdwD0RXFzOeud4UCYaggYp95XvwZO/9AZYSPLq
dcVe3BpveWrfU13/a8/No+t7wXPLM9xpsC3gmlJsHRwTeNuylk/0S/oBwBFwl8I6
DMDlVSZ0o566ZgcI3XYZmQGwXvkIoFny46rKxySIbG9sZ2QZUch7DYefNbibvNEJ
k1qrRvPvdiBMIhUJtqjk61KTSUhMQK3rEcWC3mJ28zhlnMmBp4ujGewvtzZaOsAt
P/BdoM08dBY6eGFR9sA8xEgxkZEf4s0AynHnZ9q6zsQyHUpz510LvR5QljrBIgUX
AAiFPC3NZrGpC3sx63/pkwkfvce051b3b9H6KxxMybtVjB2/bvMig+c11Ff5k/IY
oWu4Ah/yUr5JBEIhwoM5Evgogvabtu/g3jcEGV++Q6/DRm2Ix5dnfBJgkZrhPC14
M8QJciuDokBbBZzobF9FwjNc0Kg4O10qm2SXAPeGdQnCXPt2PmUMUqZl/Vrv5ABM
AlS+AdpU5qkwjWyWLE/+iVucHffbUfkMZpF+7ZT2foa4N8Sjs8PNuDfzp/ITCTCH
bR/cG4NK++yHy/9nLedlUHQ7NfVZKRsF3WxpLptqPrWji1nMYKSOZLC9+4NPYzlc
xd7KWVL01bg7UHUSlngtwa1wvi7mywA4NUVRJiY/HX6g/DlY1dOp6qXiu8xzcW8b
VLmMNej5Cf/fnU/fRLQcquLPYqEQ0ak1NNFppBcQvbMlgzEZf0bt30W6B/6srX/D
KUUmMteUZ0gBTumo/jpDUmClmqmvyg+tn3sx2g04nqJihKyWj91Goid+VXn9tp42
rpVRPOf235kd2zaTsjMLcVZBmkX/6ZhKmbkSlrDq5crXUpc3SbYr+ihrfa4H0wIE
cYo8Gslus3szMFWmj1fLi/Zs+Da6+SoZhqA420FQ02ihGNyEVrPfVeWafsNaKT95
OErAn3wKdXyjk7zhWWXkOdlVa7vLGpzIuabuecCw0L+S1DyEtk6CZJ0j/YaTs+Hu
XP8+B4YAeWCrKQUm6L90H/wJ6hshy8+E+K+2IPm8+E/yZsrpuhY9PgbFAZZRDJDs
wLXaEXoM57KhaI0HTcUZCOJtxupfRF4vf/0jO15yd8whUQB7vha5Uow/LPaZJPEM
YrOcI7JmIdzXt+zvZkJDQjMBWefYJy87Ced43VKr/PGzq2iloGFjApeW7sFpUkN4
rdw4J8e0MBt5VbNO8kfByGhIg/lheZOgubpBHtJ4BsRcRslt82Ol2pCfO5G5hL2h
zgZXxuHI3YYwcjhJbzI9EgWeJDveXkKcLH1N4Fq/CCmrzEv5YVzj/kkuqyFeSTDu
4A8zyeDqirhoGcD8fLbVPFFtgImIVlHNYuMOxcBoCA9jArHJPE34cbQXKl96jL94
r8ym/Fu6L6nLNez2q+rcjlvTpTl4M8+GDjTKB0jwBIKHaCh5L7MAUg3+tr3gILvd
gj2zzyGAPEgorBf/leKnx1IiRBP6AO4HVDHyiDe9tPN9f9lj7qE+WAzyjZ3p3Rvh
X0S4ETN/Sh2SDQLzlkFsZGNMGzWv3W4iJ5ZssCNqBsGOIm1+uV5AjfUIOZ3TV1A5
S/uaESv1Vb7Cussofbknax1wWtCtm6+OoGcTy7UWrREqdORjFhx4XVYZ7bW+CjCU
vL8OMy811HYUfk6UmKy/wxq5PNytdt/rWkSQc/mF2NeKMVgl7wavVHwiCcJQyPSp
iULjA30KsWLtZntxeZBPX+3n8TvoTWWQF7UT27ni21KTeWnNrZkC7ohkPS+T1ROu
NPZJYnbeZx20Vc8LstPaMqng8L6sgV4yrnGGt7W5GB9ban3JpxEoug6g4uELmbFY
XxrVK4Mp8TTV5+mm6HKDRYQAv2nIe6afspNf20V87sFjMiDfYyz6x+UfY3hdQfs7
V4yHnjH+TZitgZPD+XJM2rxzWSKIa5AAeW5feVTmvpSQsCr4+rvAVY747tsWNNP0
FF5SBD1Xdl2MhP9U5/AJm/ioFKm9Xlvz7yFmpzZAZmTdE/CMO4XXFxUFHTtMFSyx
+SmoBoHIEhRFFvGHkJmgUdY/QLpur1J+ycFaGDERmL/k1MH9wnvFRLWu3xh8gME3
NYR1sG4cF/KNZJJGPEiy5UvCQeXai3G5eKZEuSDKXZVpyvfWZf2CxA23bQq1QSgu
iTZarVYTiG/F7f+AdJrNwu6uHH7ndbNgTdtivw9McCBkkM9kwyvx3dzJ3ahEFucp
Gwi4tLSpDgH0GvWnDzkPG4iA1k1bmV+FF/jUSBmiHR0KdQE4LQ10WZdFQSrR4HOc
vHx+wed8HZLzOTVrPt4xUC+dKXBWHxsrxvLk/2ESg7lJ9NhkB/8/FdpeQMYzoRds
5n1GKExSj27vGMc1GsCJfTq9k9zkqHuWQk3oTAoNolRsO5YhEz9w+E//QOzklUwt
QeJ+PG3IhBVSBXtzADFQ3D+eRV0Wa7jlIyxwwjETSh3rxukwG6X7Hvxy8LguGMRb
t+ol104gIob2mCIzjcj4SBBZ/z/K76/FOy7zxdE0/TWRbsKj6pnOw3rTEp5jr7KA
AYqgSwUJuXnohbX9OmkqJ7PzjZCs9+HzfuZWc57dAXkwL+9t2BwlxhIPsHp/qmRV
6MIZlscvwiuUcg5HqBxQHlUBWc+g+DtS5PEabaZa4xWFV4uTKWGmD8urvqzlaQHO
e1ioCNpsXGBXTob9p49EnFHNlicnwAgYJ27QqjLKtQnDNDnLqzhb82aoy+D10Sqv
5LCp0sjWyvDdTSBwxDSJN5wYlJ82OdSOLnfQ4U+3EEX0a37j+je+YssLEAHf9epD
0pSHLbsAJZdMU0bLA5NjhMr+EEN0l2GhvJ7AGElILAupY7jUFOcNTyLvpVsHrX3N
wQ3UkQUlji4PNcvQsf78+k7TS0gcLyrwh6OTfsbqxz5YadUWqt+AjF2OBlOmo28N
SJVtkBLipZ2K2SqYgMvR0/YgloSSqa1rjgBWO0clYEWyNu+QI5l6+MCMce6xcIN4
rKXlR0ZEMGO/avTUhbbblV9NQI6B8sH3kxBdALmBNlavhZNNa/Cwf0oHG2C73+Tq
ePglpMyG0qNgmEFG6kktMd9jTjAKksAYpFmnEsUPMJiEt+16VnW88ds/jyaB3J6d
iEn9YJQNvNrrYo+7WDBAW6Fl3Do8FLRcBOEfGG5omb8KeiKP7e8YKXAhwSAARTHs
HfiaehlXl5bmmutA6yu9omQzng1XxG8LMrCDD6JjobClR+mRBlSx4rvbpWKOdYoZ
dKvy510M9h26qPQw9chACYwuQq09s7H6s4wA+02pRMoC9vqoSDXERDIbYzbqLrps
V6n8NGGTXwA/WiLNb6ewRsCyYvklLT7ibNq4iJglfjpQyAolmLPmJG16CFrbf1v5
JWYsYO0VzSPpvaETCUqXMHgq20Cptmv+k4EoiIphZ9L1jAD4cQSTNOcsOs/tgFOo
5KLTj9RITrEJqfMqg25F4n00mefQpgBpURTUCIcYNmQapw3o4iM0Bmn0TNXtRDu+
/lxrVjykcKtoNbJDavP1C5/EZT9UGjnX+skHiBa5N552e6qABLdc3VUyAPP9SBEX
0I0nY+Mbea8WeSmpTJ8ButL1MY84iiJNoR3kwuQejc7qQobyGORpoV9+yNkH9Cvw
S2ZFziQY4Bd5LymwK+o2STAAPORTY5sN9zrsBKeHqfHXwXdjq2K55RZEsd8DBIoy
R+aGQnJipfT8bk/kigFoh3WRhATxqcJpczWSFFQ7Ckj7X21PdkKRrmcqC3/8/1la
p5Q+1eXwBAkSb0BZZjjdYuFkgsMiOXhk0OK1clEoKIcyQ1vwclj5mb2fzFDBQpOz
ePU184rrFaxW8Yjrft7/w2IkAicLoA/IZ2ixYenuZCVoRvZLCr+baCzQToE8f82y
6MMEIfIygF67fo4PaKEXFVGddxL6fBM9y4SlETDmhSNVfQnXSzK/+9MwLVJmEudW
Oad3hecjCF6dfJSM4gqXUkoHoBS+u5AR1MibsftdVBle56xCyHppRrXGGi1ayKy7
TI0Me6bq/jg9UHv7FVSHHu7kXVyLRm0tzypyEJFc1iKP+/Ldq3r9rkML0CoQI6mm
WBlXYr7OZbmqzvkRUROqzQXSiNl/XzBzG2GLyQXDeVz8n7i72kzHL2HJgKvoq2PK
rX5rjDj0ztEgBRYbsxVMfUeeEajG2zdXSkfGyEimMwcSzFsq8g/SVolzIU+MFln7
YytldQuqe5jgywyCvuFo2Kg1wYFY1nNbXThtS3+34xKlZu3GW3TzvQI0kQzE3Bay
Lv2N0rdjZXpkX8Tk5EXWVaursWhOeYd8L369jtvGiuB3YRHb8tJKi7VIgAQkTrY8
KiASXPkB3qDeE6QpTMOZMts2tFP6B2icp5VPr+FUnR4kbiHQXxJGfzcdlkevfrO5
BwwEz7BlhTrA0YoWIi/Q98DKeyk3YZ5RHv+HH4f31Bcb21casVsbbzfqnHuCA51h
4pOTnnbxPUcddnfpDm1GjCgiVdKELme2g1/If6i5c0FzYoAk0FdyLaGX3QW19uGy
jfSYa/RFPuTLVzS/+7PxiLj7Ihs/y5hDggWb4GgnAoWkCl2wsiMN6tgJCO3lwCYI
bu8HNHSZpCWcRQ1A7lYybU3NJm+X94B+1Ai/twQSP00HKe18dBtsycnFkmSniaxD
6IxIi6s3U52YJGGp49MWR7erDP5sMeNAlUvQ643X6AMnUUl5jEe+RASuPYs/9Rpp
RwTncFO5meqOAKd4JumoIgU9vV6B+Cg0S2ULZPjSR9OD6FxMs2aPPIFZn6S3PMUX
LYNhE4wP8Dczl2r2ewJOsksRFUtmyNO10UsYfxmOugpsfj/1L6XZHKNxuaGtuu6l
2yZtazF7eSG4jFWZZteA4Kbj5J4XV1+1kbNvugjjkd5BA2z5FtED4Ktf4t7xzJfG
LDqL+qGwXrFJp0SiN/1YFSPmjYXIV8SgcTuzXk+m227X+JwY55p1572fEKZ7sIax
TNRrA4s1cI/5krNx4CfuSYPCqB95syxPO0pIkjfOIOVZTmWjRxQr7xDi+6eibVQn
0UGuPAzLq83fAmlwK0jmJc+WQib8OKF5KxXsuRbNkRsfvZUlOaxJmGwjQWP4fHSn
0IlFQ4xS08yvYpecifKh1ZBepe/PMYq7/s1K8nRUyzPBbXnBuEnN1Mzx6PPSEebi
GEjdU5sgHaEjuVxBguXvXEnZwyvf9Cb1cyGne1nKqrBZMX7NLAyl8gOYr1Ah+tSK
ob6CYEzbiWs90ehK2DFPG2W6Eo+x3IdfVMDhdzK1ruWgIEjlNxZ97QB81x2zHhoV
Ks/VmDoeJ4KWuyjRS49UlszLd8uZpxjFae1/YR4v1WvqJyo7A6w7zUiTULlum8LA
pUE/IB3TAOE9RDVktlLsefJKwDcpxpX0eeyodb5ZJ6EIG/SvIj9JkEhW4a+d/5N0
4qPJ2oKm3ISISSZSCQU4tjOqNbaTZASIUQn73hcH68cM+x9bAOwaylHFm/JEYmeq
hoj6bf/6QB1btkBdedkPp5C6W77s85CFJqTSzuRoKwTELXl0IXUppPAj64MHvy8W
fzPUckSHS4eP+Ff5BaP9WLOQ9XynOLr8pm3UbMSlZd56QmGPutzJFCrYbHdP4e16
ic5sYy7KYdZv8PsDXhGevolswqMhos1QoItqt6q2p0Qm8sdXl0zX7zC8EFaLdArq
21Meujn62aEoS6xmODzaHtwMIZ7D4X6/bo7hEYIQR2pxJfZSOjycOxLzHvieqwwF
3a1xM7uE2lW2+omX4i7gHRDFD51tYH/UH9ZF/TucVIcRMiisOJJF2TxQgLo4kUtN
nJtY/W90C9NQOq8LOWzxXUtocqLGabWjBIG5TYSjj1yPXiKafFKCnmpkR24hNEU/
MzMbKGQYj7/CVI34tOldqgBmVtNrS6cIbUVnVgnfggGaStr3FOlo31mrWDR83+Pa
AQn2rnkHKmoUJqL8KZs6th4dg71cNhFMHc7eqfwuTamJNAh4x31mOvzOc+j66STI
ei/aM72DVbeQeSYp6fovZ/hLSNhcmYqLvCEa94nH0ik3dp9eOj2PyxPak1FJ4aRd
ASwqbf9lT+lPpth5ZA6mtpou1LozLVW7gW3reeGxPX3B2oz/TXbEGv2n+7xetPTg
m5JysiOR4UcPRAtrMZKsYOpqPNguX5QUdXKqMHYQQLdNjfrP0oDKr8dJfQTEul3v
tyeOIpBGkcZXeT5Pjf5JMdGvqzhSjt+J+WtQdMEsO5ZoERbqpD9iByWhZ98UUyl9
PlcBKcrurNfxCQqCVz1XsO2Vh4tNcaYt4ucE7Ryp5w5dtn6OleDjeD2mRx6GAPYS
7VZ6Q232GRuklxK182AEdzvoHR7/sApQdGftTPbekgDdeMqpBuKRaGNhXEqtcbtX
MsHJhrTJy7TfNTGgMq5gMTAjIzh0j7jMcKgOIWDDIEW4OYJl90kaEsxbVAgkiWwC
CaGWz8rGMP44mNReY9rQAShuzrk8eFwnxqPDH4HLnnGYG0zGMU4t8CEnUFGZU0Y9
jSgVaTPLXSZQSDdWgEB0u0Z0TiGozHGEhiRG9perI/PcT+A9TKRFfaMQLMlmAerk
ZDKofJKCssDnlVAAOqOdK7wsh+WM6il9PCfcI3ljo5m3ISYVvGfFbmwHUn0Q59u2
5aUH7doC2s/snJc9Y0ulgyGvbmS7d4bq4oOR6RUaqm6QIerXy+cLlQAuLJdrLhgO
cZpvQj5Uh5rX8PtZDVLmZjNTvbUg+FVQJrCpL/qvv/AsuOpSfoI7GT7DYG9f9UyO
YytMXoXnpHkWattOhvRmRaqocxhrCYWmP1g8HddwUEOtFUwzzRvLMwuzYUrhKR8t
3OvuVR+P7ck1zINFhzheJI/e6KaRh+DCl97pWGs+u+opCy6D3XCgnIyi6B3arL55
4feJIxjjTxPKX0g5OHoInxrZlcl8lROHB+vT668qbbyg+CeIUNemT5oKQP4B+spZ
pp7fbQobQ4JGv8EZPDac6Nw0lNPwUQ8Ejc0IHssZJvZ/sPSyQPOHwUHQD9TOyNBb
SRWdXVLx6qdBx187ss2fxE4xXLSLoMSAfV7YkbLLgYukLH+2uLeevGoFRzcC1O2n
sV0Tzj1v9KhAVh1Rdk8SMpc9tPJEK7owwDtf50RALzSrjjCXoEYjZ0wHWVNOW3tL
CYmMBspaMx16YvXPwbdlD5fI9e42d5miGVTyMKydAYt/b2mw7jjl9BCCV9mkSQCU
G4cD62lJAqRjLtvPL1YYZ/VWt585wDFklMvXIzkks/HOlmlodGzqaCg+/HmYBXWb
RbkePoc20PKCxsg6Ekf/u7hDJkTxfusLYrs1yV4fARTl8uK56eUCTkdVoSANNKc1
jPMIutxMnu61EdWMMkyU1JVP2OkIDPQ4BX+U+MPzV9oVHINPTdUQe6JZhgUNqz/W
/NjMfaDp3UhngsPaAOK+YwjidgXdY01zgRd/IkkDSqhOvYwRV3uUuz8jV0SA0t7v
hjZ93f9WDjzgfCyXYd2iwm0iBxih/3jRZxuRCaoTk/FTIYaA4l6GB1qvXEB85HAt
xXmmA/C830erogxFaG55NitCt1RYaQvCMhoMh76GhbdXOlVQwztSSIsPtgUNZXMb
6LmmIVf9SObME5XH7Mwz6LTcnVAEgCPcJzFHQdybv+dTtddxYrlgeo525er3gUjG
BJNMWnCC54uWz7y57vWWnPD2MG+A/e9Op+03jU+QekLEv+SrVpEXAgKb7SYx9el3
dLuxS3dKzgcaeeelryo6j7r7qnP7sZl3RrVXdCXldY5qVvA44jYlEFWkT7FMkttT
OcFFg32BvjKF697OPqLcy4rTRW5oxevtbo64lCPkiUVrF4y0mO/tU/X1C38nhyog
OKXWkrmGF8SRgiYyKPgtRvmg4XzuJdTl7hA3gjDLkcqbuxRbq7v8laQERf+SOInl
JsfiKoOTh+dujqwI/EoMQJjWPkWESymGVRoVUexP9c4gXKZAtLps2DnaidBLYO0s
3xyqnebl3NJJ72VRCCMFDHY3eyzBBfnTSrxlUdvBdghKN05WU0m0gUTCR2kKBv7n
98hiJNONjx3YWQTVno+414VQWSyhTtc3plc1AJ3EfpyK5eGu0TIq94VHmZtx9kSZ
FaMx292QEFKAj6Of9d/nzqIkrAcZG6kKnbT951YdHac94nTB1FFzFtP29341MbJn
IMren4a++qXFQ2hjOeA2i6Roi/BGqdiNPlGe7Nr/YUDixcSwyiYNqZWw4zFFPdWv
1yjXTj89INxE882Wo2CXMyC19lvgJB6kAT+YIvcrXW9xepEkVVuA0poSOJSWei6L
0yyWEd8SfW/ljaDwiNTLB+W0MDuuuBDLY81Obr269cLR6ck6clylthH24njFpyyP
xoV54DLXEcTuvpQoTHOJ9LehOWfWjSTDJUdDL1+MZwtaJ/d5pbcse+0s+QkToMUo
qnhh1c8iDUpzmRaXQL4ZdYkGsh4jEduEpVIEmI45LIR1ZNix/x4B3q6Lp+UuLGXO
5yEqTbYypieSk1y9U03s++XXkJHUc35xqPUlTVJFRUFlofQUeEoi8VoBLoveq3pB
/Tyh7DkA476fQAK/opM2DWzqqPQH7gdrPM03CPpMVz6nqBlTBvIzDddM8mTM5E3z
w4RY7I+ALIm2KHeB9Ra2Nn9LjBswylZEGoYK2+7iQ9Bl/KW28vr0WFICPUdCiYSo
daJfHcHAq/HZ9ht5RUFhUOVSkkdDWIF6nOGmxEH9aPwDVZcW/IvNe1e+UPkNEMdY
p8FtcUvEGbrGlturCjIgUurUXqBEiwLq8tLud4ieP/oePvQ3lyQANnYAyXEOgN10
01wU/pjn8Jsat1HDDwWkODAQ3wZSeOqYpYSbkEVY9iuXon2iiXBaqq2iWZwbZe3r
hE0xDlM9lOc44yF7aPpor9xF4ePKNV71F5SGIjlPd/4DqEYYKcrYmyYzggx28m2X
Qp+V2eJL1cnIkrNt5P3aqvBu03zspDWXfEHSLeIpQyKLF4tZ15RkTa7ZzpCxwFof
xhG7fQ8vK6AutMpnmhSE+32OnXdpqswVpc4Bg/9E0gCjYITN0aJoOj8ZFXkZ4FsF
7ZveySOvwHDF4KZbXIGktVJjk748aaygorNpcppNkH/JoRp524YWUk3mddQv/S0K
xf4tD58navkJRaU9Mei+g5V4YimRR/qoPkyP8WxYmhCd7JEdLALzVHiqm/GaLLkY
c8JUBrq+vEPxBovyElNgzOWjfodxalzISDfTbRqGq1pfwUG7WoTL2/ufGjkCd9Vf
mBOPw5CCRNNqZSeKh2DZiUBxu3KDmGHMjTF3uN8FLt4zeq38Vt0VfmO1YMm/ybu1
Y2kxd5pYo3ecvrwsyGY6qRlVY9/C/7cOGHMhAUdi60l/TNbKM5Ja5BEwv1qrIVp3
76bnu03zynUWcwx2i79icP9GDFMJzsJXZBExZpzcV0GQJsMsnq0tCGFwUw2O9p4O
BUgi06SuPbVDuap7aNTMVHc6dAQpRh+qG2TFBJV4jHFO/FFPsJv+xYIs4La8xmC5
UtvIA6DJ+FEbux9CcXgxAuElWgpk1MeOq4IY8sbqOjtcvyHdDz5k7+EQBwZjIK5K
GGFX8k+J6RIihsqvdSxl+7xIaK6AqW2vlx2TNemMTcv1I3EoOh7Xq1pYjhb0Jezg
pXvDLga0ZuS5aN4ZEUBAInEE0AK6LEGwwblL3HbC0VdOp82FDR8aobplXs8fCwk9
NECfhXwW1mYwgn41uHKgPZdVHmWVjl/wfPFFV1zWT4hnoiQNCEqEDuNujP3N5tJ0
idjK1PCBB8ooRCNHYDNsKpZCgHDnoaQ9v57Hay92bRLe905fmaccSNx4wb2QITaD
+5DCnOcVDWe5qXXKEBPVf65CAUlXCxj8RSpj0dI7FefanLdEaIrcJFRw6lVyLhtW
i+l31lHg3sWjX15yxHXRPOIOT2D9DvYo4iXMOzCxQKsET+Ji7lwSJK4w8hH3sCXJ
xPwqYabNqDs+YXANHXKIgoFEASjhpyAeepKZhEToPwYgMjvc86dOf4PFRDzNe0HL
wo98YYcTVGs4gzVQe7D6vx7qIpg0A8E3IjoyWaqs/WfViTTrGhfgEeisqFFRq7dl
KRMjW+H4tBDaBjHmVutd3ss3vK7KN8silW7VaAZrVHDAsNtB/MzKpRNVNtWjhAXD
jpR6yRIHlfgP3JDY8M6D7zqgoDj07A5H3FZB9sLHrsClO14agszvUYAo7c1lEONY
6ubPoK3UMMB9PvQRTbFBmsuUhQLH5oHhQH6FHiWjDRdZW2zGW2IbGGUoqiimLQk1
NKXooVgYI21SChuFtA+OmgcSOfIRu96zhoP4OvTe4gNMi2XFUfgD5uchoeR918dN
EtgFlCq+PU08VlNmPouKST/zFlJ9EtE0K5Ucyotb3B9A/HHrnWdffaXWy3UfJW80
wTUvWbeFtutSQTNwC96aeIjd3SRFFs1h2rE31ON04+QObZVvk+9NgVkYBrwZ717J
B1i1sGHZUHqCmBEGaIy7sMT8Chj2BP/lO6qFARSKJ4xw9EBUvIYKhs9PV2hfCgqi
uoF+O7rgEeZuts3IGTfx5EM+YXJn2bZ6cQUTpeTw8IGaQvjCZ3YwgxI3DPpQxxnL
zTl3sgLm+Qbsbs/soOACFF5m3u5EP/v7Ez8m5vS3M7s3noXjd2Wh3bOdtSifjaS2
2LKGgtxmdr2TVo73Bn72ZmUemW0pv1vfUYO1N11+OEF+mVq95RE8hwATkpZtZ3n1
dxmcTQDc2JA/VSxpKnihZZtOQLaHXK2NXsrO5LA2HRYR/1XW5OZ/kIFutfyIVSEn
clW6yFRHdEPNEnc9i9ocWCgMPYadgZg5+NjZcjHPl+VUkNbAO+d+ag6Mwihb+S08
lrz41wvKJOAryKMkv/8orIZ8WI0T8V6v9hdObncm+z+a64B2oMXTr2R5SrLwUEjB
pZoUrVFYMP0o9Lcr3tDhgsEdS008B36d0RM8pJfplX67+SsM0RYklrTSQ0dCUO2g
gu+wKPc9GSEv9dyFEkLp/griX5ctwNuVgf2aUoGdBFA2f8HbCFruVNj/Ej2c8eRv
XO/xXC8Rz78gpVM3G4wYuBTfEIEEnddIdbmIvNnsaYltfnZRIg+Vkt//6zzagphK
V6lj4qa1b8JRyRmrcChGHzJmFSC4n2zHqNhrVj0g+ZXazt1MteOFQNBmzDfNH/ce
H58YLaYmRIhVZHeMT7M7LHHiDzLtAyK6wSWQmkfeSYmUktanCM2lVZZlb1HPyJfx
WRu+s73WU2Px7vRA/9zNrn6C/V68G5bynN3LTxTFoZ+XiFLQuKZwBgDxFj7OiPOj
ESVO/a2M7RgW856YkDunL3xBvOFHl2s0GHcRrNOMLTsPe3FeOBvXr1jGiTb6NXss
LWNUqnvdt221sQqZhCfs/FYJ8Udb2eex+lYEsHahAMD6PphUkPFLcX2uWob43Hml
x4wmeunoeIz7VYGbbA5c9PuwjAsqjd8DC37AK2sfYiSOoyOHC1PUpXhpdDC7CxDl
tLt40xv656Ez/JTTQ7LRCsOsNcsMI/POSwmNWm1f5PusNtyICysBjo7HZQ0ts1q7
zaDB3nxhCWHw+bQM4a1n+1EByBhPfiEluwfyzmG+6nJQej0zsnEMERZD98InCftd
saO1ffO8SysAcPDJqsog+uOvoAA10hxeM7/GW6zDTr1R3/7d6ikqjlcLwZv+Fkop
LQ0HdYMJdflqmbqkPMl6WuPC8tNe68HW9SXU/youip+JhtMeJcCsQq4FhGc3J01m
faXOd0NPIPttQee738vM35wUkbENWH/r9FKIuUINuCI/FXPb9TwYmWyBe228xBcp
3mQobutV+H54YxdWqXJDUXoA+6vgDhndUhkwsjs6EWUka2Q9/eJ4lvjVMdLyVlPg
L3knHdN0TKANHHXDXOtv8hfjB2YH/+gzn5M28CvfxT6uvAVljyhppMiCDRl7yTHS
oHrF7LBLo1gYmJ2DoXferMMKWXdmFs/V+fl0W86LVIFZeDFC6JGfd9ZJFjn1kCPb
2M7sukcP5+dUNtOrPsXHVly0dec2b9Vzr83K30rmBBmMoAFN9ZNslhvy8IcfBaMV
jbYVkyD8DLwOnKVVVBY8n2RcNhr40wpg5tAXpz4njZwpqITuMIwQed75UgTKvlKu
9nm7pCfbDiayqair90neGpwdZcRl1CgY8uPB/LIPT7bX4IVT/HxaMIwJ8KifaEDo
crpJba8DClAUvNZoFX2UEKp5G9mdGmCirh0CqOpLirKyl3EEGLi5oCll+ybKRC5H
eGIa3ADDIjliKe8WfTCgFWw80LL3LzfQoYteTniTyIbQPWCDUkj8QJ6WYeMhJvRL
sGpF9wM1bIZGc5SGGaOLDhl45vpANujrquAN1urkXeNVKiMEUGKoQoci4re0dnvZ
127MKnrfrJAwlrZIuXC92AVq3QxNFm1/+3/lfzsP1cU2bFWjHT1x+cY+dHz22vLN
eQwaK0ZPKNfSFKuCJMkQ8+FLgQZ9qMbpzE96Y3Agbk2MKa/zCnvimq/nIGrya+yV
2/03b2X2IWT9vSXsx5qSJxmzm+AovkCU2SYyQf0xaBfCDCsJy5tzWHugH3EkAGyf
SYRXxywGq8qmjQma907wGtPqQTZ8NdNR/UMX7+rUNNufMxF7BXNEvXMvKOQilKeK
R6AaN3m0CsoEVUf/A+2ZPpDoGOAsO8ZJBDQ92Fw4whN1uKZDby57g3k3pWuo/KEL
1oCmIH/kGWy4pZmREZA+zrLL8bTmyNzCfRVSQZFObOIZhDSVGMRVXi4lCxh46l3x
UTDv2BYgUUf+k01LWKHWzxKXOA4huPPydVvR3YqWxxDDVp87lSNbAcXbAAGtLVSZ
3YljXlvwjGBO3BfNjkysEQov+f5WDrIYhN4pvikovu9295WPz5910E/BI4yArCok
xvOvXfaBdj+cGLz1QKiu2cOEpWnOsaeFEWLhcQp2mEP7SmLVA+OXUX0bMSNSsAHt
jjivrYDsYc+wom/Cco75v8Aclo2oB8M3SjAOOeeVJKa4G1kgjenuWLWPXxyXCQp2
fSlzjcluuSnTpGZGA8UfowXbadPnGLsoY4YV8a4Fq16zGPoUDyhRbj02SI+DzoWo
RxL15l5HMU4QtjK5fxBWH82yNlHtRPue/3/YU6b6K6IpsmMWif9bSMw0MJbCMpcH
GMfrhDC5T1dF6yUOMyP1V3iKIYH0E2Na2e7mwGjtWx8qgAZ+atZN8h5AHiVTLrdB
U9ZPjO3a9gX/J1uuPRSZJ2yamm2SDG2bc9s9CYZhFiR7QBPTR6cHYzIjW0qb+SiH
Z7UznMWJYt6YgTootQ2JwC4UIcvzIyiW+MLxGDbSDxMo4d97lhWxHDR4B4PgiSoi
hev9e5YVPs4Zj+j2E7bwiN9oMVPLOifn4ou0i+GptUGdbcqtWukVsCqLGc5+hS8D
SW/WvQTk1k3oLJphCiOcFcOQ2N5xC74/J9aChPjo9sYenpOROMuN/WTu4uE3/qmg
KNiAcgxkjepcBWesKVvWv8HBBXWmbkvPSt8UGWRMqWyw7XYrphFn7KsanwDB/Z4C
kOLjY8JyUQwA29HHRv1vvjKsfJz+o4kx64qo1s8WTuWitIwdAdeF8VT7rv55+Bbj
lEiH4uUwQo+0vlX2VxodJowPiZKhVnM1zag0mm8RB3CzPbhq0vkAoYb7oYSgJoT/
HkJYQMQpGymu/DKwRSPLVPcYGNjkoU513QksvZUtq4gGsmBkLAOSCHtwIg1Ql2Jd
4fJ6cVg+IMsAPJ1Z9I2SIgAfVoylU6DWVBKrsdqTtrz/DYoggERXgjdaZsoom+hG
HjcTRQNT18V+ZiNyN/82sBtM/elRc9jqTNQdTbgWK3hF92u3foHOin/F4GACjwQE
0UyHGaVvTnH5SD8c4N4imjq29jFzZboAYiS8vxmDdVC2WPMjNhfSwJ1E+DiXU0Uj
lQoQqbBn3CBgYD2GsF+4rH1OAnS/SGCTLxG0p6tc/qeI9b7mx5sDk5NhNs8r6Sta
ZAFVvZuoeVsf2vb1JV56Go+Q5eDWm90G16fME7cGaeNSpERcJ2VWtUmz5mmpM2lW
zAtmp9dnGIlzTJrOaB1V6uf1I2KrzxdEElfOCqTd9OWz6uDfjcNT6Nx6OGh3+yh+
eYNtrBEeAjFNMZvDAZXHGcfi5pZJqzvxXqimAwyWQ+UWGgxxhmAJ10vIkqrMyL+f
EcJ2kvcikG994fuNyWef0j2RitF72vaqwtJN6aZqi3Vw5t5gy8pUMDinC2Y9s1Sz
20XucXwTm0k48MFm/66aVqp0sKigTUmweRnj7RfTyFurybjtAli04sQu4MYvUGxQ
r1bwAbPI5IB2iIVaEF5JFw40wI42JqGf22VBvS7NV4MkvSjhNwiTDUYdixrjv2re
Rku6+j4u0ly26tUYAQ9jrZMls25Bjxzdbz2aKUjiZL6o/HiZeDOJ+RzCfc8UPBRT
UcvN9IOul6QD922189UaMxGgjVYWYM0nE8J52YwQcVEh9dg2TXmm2f+iVLmTwO94
AVFDOEAzVdfqgnhjpPvNOPl+J2qyDPRzY8WqsRdKpd9i1iJvMK6ssWbLvn2p0NYx
vohPc7iMqilLUhxNRC2I7PxLVs3Aq65DYQguBsDLcgylcIf86stt51O5EKAcndyt
TnS6cXBxUJSZHnDLkIZNempdzxf27l7pd8wGPJv7FT7yxGdIzEa+vlKRLttt9jQP
N5OQ6K7wqW2W7va8MbaPxKOHIDondtoUSSnhlsfYSfz56bse1TcVMxwIU2SjG5Fg
DA2+uJFRJlSMYnqtvx+cYphjhE335EKf3o0zdqmT3Y9p7+RypurFxTvfZsLpbX14
cyEaBFWTxfG3862mSyqLSfmd36Q0VRSUpXd1sumLU6kAU7wPH+gpxpwXf8eZTo2+
h/54IL9XeQtuzPAILoyWF6+T+vxAn9n788iMwXO4cLDHzSCd7PW+pNsJhviTErGW
VQpzwwY22D0XXZHONMlUyeCf6xlOXehClWw/yk2mMs5vfMyL1vRsPsWIIfFuFqXo
6RCfAPnEGhDs1XazFX11bNWW8Iv7SS32d8E81EMrAhTNatiXrmk+cLSrloPW8o0h
LIKKknvJLMoaAd/IyHcTIEsjqMnq+Mmu0TAGo6xZMYzdipC1L81YvW0agoVoke78
0e44cszwwMXIPwxtUQVSATpThZ6+BP+1spTZDSo2vC+Ef2ggc06qzJ5lcnEJ96Rt
G1RaBIkI46UD7jjRfSph9pdoDHGxDgU7ldz/MzCyxq2EXGTdUDlX+S/SJxI6DUY4
0l06GKv4thYPdnCIdQpeHr09tuM7VwJXoMkv64ob/M2oQgkWokNfBiwrKMG6yRYa
NsxYMAya986fhmm+6WL81sspwD2NkMZGzVvTCiGRbCAWYtD0ubEKQdwlMouAhysF
HxlFtfs5YCkEzuDSwoROO1nqh4rTQJ4OT944edVT7c1FXavquyE8DpQrVtFiujex
0LV4uBa0PvT451PS6NK+3mwDusS6LpUrZy9e/qh9Ldg0jExVBy+00Hd8XSmkMAoC
KjcmxGB3b6G/utoqJqL11Je7QPwmVt6NJVgVbIMAvS+mRk+lvwnWe33jYEp5/T1w
inyDJwEDbuo4tahvyYJhBQA/CqeakJpdeCXCj6iqVG6vcWzyQ2WIbmJqa+DEEN18
Fk/t+QVbKMhkwZ/u8+sq2LHG1+/VRBw+TMC4eAM9U7rJasO5nUNCij5I/nF2H+RO
JL3d3t9eDWL1pOEB/alainq5lrFVEtUgPIpjh6RRvfeZzDL5MjII2Dxer98QzA8B
CmuRJmVgkL4U+nt+JTcFw+9RxeKyNZuOvLh8zYELLaxjClh1nFD726IFsg1Wqtu/
6s0wL1cQN3src9/fD9db3g1Wja53Boidb/yF4zwMdODeb72nH7HCI86unpkJHAHW
MZypUD2VGVfbRn828SlJHJeVHvhXEImXe46g5sJenanz4wdnUTXauxz1fT5DrsZ5
XlzQzd2qXx9s1PEcYW/q1zwCraF8lMrHhT5PJ2o7UVoZWDu2PsgnD2nsMNVYB9qf
ft8XE9taoYuBQNfNcse3WNE6HtLUrae9hZloNJTHAUhGtwL4K96ZPOWvHTMoC7cs
wI9gY/3x5sRkjr8yEeOWTj7RlZEZc/Tu2a1DCIS0e152AQxapQI0oBs8T7krUzRk
5N/yV9ca4YYN/DVs0crGlc3HqrKLYAgtLZZ2JTNO7/PqotJDb60CfLtxrHVM62+z
bYDNtuzHh3FZU6xTWzWux5BM1ZHLbrOCMTtkD6u2wz269VxsUuAYOBwvZB1sVkNW
leYLIVWA3C/9a8uWVdHzxa/8rcI+mJh9StApOxPtqqY1/9+4I5ghwSiX42ItR8P0
TynOttl8LodH35UP34UGrUFpowmCAafPw0nXpIDPzCi5hhIh97nQTjX0PbMRDLbm
8DUrcHcSPFmTIZP9B5M3cBXz6NeJw9H4CtTAeY3FkEsgOhIrv51R5cKd8hdxylBA
J73EsXTTT4FdrnKbXHVihphHnpCPkNEoBe6mp2rvoe9mSB/zVhv+laSqBv2KvGht
Ok9ChQ0IMTklzHp5NH3E3SavWg+PKL/CtVPJkCPqz/vVETUgbuhAqePQNv6OIFEm
kU2GgczRZ5q2ek18+B/O24FyoMrM/AhZmxxE367dyEAziDrO8ziBQDQaNsmTfFIA
vKyjhhJqVV1j8mNXjzvRcBMRTVKh/PgvET2hBpn64D7MbYR4IZ7YE8TSQkj7qHVy
4aUiDfPSKFZ8oddTKPBx1nRKbz3664DfVDvFdoTUopELjXfN05u+LxKaTnJakc95
e5PQfXPSXIs0pi/zPp6vn+GlMExsYQNBxj9uAw6gAEAbCS1RYMnmB5vKg3P0aMEe
5zMAjXxKv4jyMk4NWkkW/enTVj7HsyYL5IZ2n5bq091t8ebn9T5KjEAYwtyFw6y1
Ovow7k/fi8mOs2Zj/Br0+Ydicp0gtgsLASWq0plkhWTrr7CLmSAdqpqYqg1JvkEf
Lh41wYGkwdbZCmNAepInI6Sc8YqKCNfsBX10xfYOPypqKEdnxe0ZfWVXAOJ49QPL
l7/1TxkNhrTCtXXMsf2PH0/BcM4Y69gc1cV2V2f25xa+j9m4w++RYxISGtR/a2nz
I+Huy1VRsGu2yrgIsXFTiptdUj/OMlR4VXA5MMWJG04RHOIe+4t+UjBLh7S4nX75
Gr2K9/8eg5p1W7VjxOYzIr4eEHHkCKZjKwffZNiocS6pQEfzpZLLhxxPpFBbRM7P
SoOegotGCY8FMrHnlQEAPdZEGSYg1gAaW/vx23CbN1NMopSRj8OU7PubxZsIiY4f
9bsQ0AnctwQ0aBANEzlknnQWE1zeDkkLrf1tPW/Gh45bgN7D42RsmKMbeYuR9g8h
tDN9oJjjVJhkcDElHwNqq+C5fbyixTKuSsVeUZcpUuKbJEa5i4RHYwG2VV0j6zF5
eNHjzByD6PD9VUqiWwXXIR2GXS3cXDgeRQLjGclP/Y/sO/S++nxSpJRAni51Cww5
yKNhxavYHSf5Q+ra9ckVbO8e1j9FbMahFgYP9PSwzp1KpGBymcGrExBW4RmcynYs
Sout0nIC33Q/VWq17+4afiRC3WpeBmcvvFh3z8Tj+ZiFTB57ODK2mgFSTmQRec7M
nvfNww/X5SG3nNtxz2bWDqoooEIMeP8YmtsD1Ew3eBr1DSH23HqljQrT7qqs9j7K
5Y6HZXENdHRUKQhASBnH3PoqZfkpyb6xA/y/o1Kr1FbgG2zXeMg5IhGMxm+b56Pn
m0zyM8iuMvvnLT9DJMzs8zAK2B6bBs0AIpEgGnnVDXUQ9208YpHkDNCEeN0/Shso
TN8HeivslvD9/49vTDV1ZvZt9WLPsBG2oNUhpfjZ9G1FTjoYNjVplmGj3d5TUqSP
RD3IeQkDXZCvNke+Rky1yQ+J78EWVXYjSh6aXL09cB/biDocewKuCQO8PJY47ro6
3ZXtxhkOr6lZ62Oix/fKOWXnboxZTx5VkuHnU6LzCKHc7i5NKg8u7XpoRJ2RZjOb
fHsX4oIlBQEUPoa8MrVF7hkJLMb/MlXhbYEZuAOrB1cFdS9iLS5MtSHDWpZ3MCt9
12p7whZAh6wFxI8kE0ylqWzeFaoZ8KaiLJINEeFYBdv/d7c7ZqJrUo+1nhI2tozq
XAZZMpJLITAnndQZILadoUn0uV7xnjIpnUkRujpoGCcrIgr3MeFFgKESPONCxurE
Nf/JQk6ZCpQIh3Ij6+VDDuWHnS4ZxiS6wqKjyma0kZ2UwFQXpUaNmTW89UVoZcWf
cF5V/qeDcZFFOjUmZ40UTDaLDQnwRiKzG1mZXKtVw3pyr18KUJD0l/9ZusWe+wCx
P0Fto1MOfOuLGcPtNRZrOlnzkSVynaY5FOtMhgL1t5AfmECqPUs+soAllrtsOCyV
bLC4h2Erc7taP4mc/GIqhe1fb/CkT9TRSQzVG2uoUddub39M0H8SugjvvqW3R1RJ
EW5M8v8wsTVW0qL/99aq86a+sLNs+hRqoRb3XzAtGzaI64CrSAfOurhUr+rGL2wG
gBcX9x9rbEHuZ2V1lW8zjzRMc0gwQVrawuJZixGitlM1fbaSnqjzjZhOlU6rzJBE
l9Be2cNx1aeawcJgx99hOxjY/5wTA8rSjNaAyr9dxDbQLC98rSy3lgRdOV75+rdi
Ae8ity1r0nLPAaj0gmMzDLxaL1z4gfc7TU8ApMS9Cv5h53LzwkO1DLCqG9oBok/C
RaUNfAbola16TkDMKr9g4qjP5bziTfthwVAds5VP9aFdSAMDWYPewqV45y2Y0dyd
RDzEl/CzLW9+LO+jo7qdF00oF31YofFwr44MkBRnm4HcYEGjMYj1FHDLy4z4++fM
cw1EZP0aphSzuGYitODQ2g8I3NG12L/K3TElUffr9vazdJBoy1Lw+pVYfHg3xl8E
h14mYNfubjooods3JCB31XvqaBxAzB1y7Vle3UjvEF0SfREq5K7+GJiwtIXQSy0v
dcMwcgf9tkxo/ZMqHsZ/EP2XXy1pVbcBUzcxcO9RmHdSbbxZJG0g7ik82rwujt72
GP/pE1Q3pfwbyanYOU9Pn7/4KYL+haaz90JlrFehZ5OhXkW1Flmkn3kkbx8KvJs0
BIFMmsks/uHe9FeodVjVN/Q3EMagtw/I72wZvI+Zu5TPQGRDopMTFLpA4oDpdv8J
qN4kMUKHQIHRXbILQ5Wi6TTZl8Uh3GqdOaOF2kHVK8UWpoQCkv+Qg7UnN2pHk67J
YhrfurZnGs/tuDJP1KIY+0HvBwNAVMOpaL/K9XakAwnmwa10n5fWwK89eX/VY/VA
AaPytMAd5ifEcf8A4mJHaZxlPtK0UctPdNJT0rIv3/uQaj8q4OlUKkMd6V8yAz7b
PWOYnhzjJNgC7jG4KPqOD6KcVmwMfRNbmfMfeqhveqGTmtpZFbw+FNFIxYCzCokT
BlLuYR5fUIeQ1/Z4WNlXmjssJRCTN3xPDyHO80hmwo3513/b3mselfhweipe0ieP
03TRB0kLmfMU5ktbvwSfcSMaKcUElAxr/SXmfP2DvXrbRsKqrp3SEgkMXE9PvOcd
pscstHFqO6I7nmONxD9ufiJputLh0KZy4hh+i/6RjYbRtP1gz7if15w+m2XN+9Cu
daYKlNZDo3eazD5tHlteR1xH/FYhzQUtT8oopYWvz93wWXdERU3fgXjq12/HhHg6
jpiOuKB8JWcOaEG1w5ERxwsqM4QPm+T3lanO4qdzf8lngeJvgAdmji4h4C8zFEw5
QbFJo9up+J/gXax3m1y/mTgQC8vSPDFmAK5g5w2gycQCe7gBrTLGJwknl9Pqs+m+
UmHLZnyR0E4jxE9ylulSr0jb2515KvZBnrm7i/ojlxMiz6r1tLO2rbV+U+HTP45e
l4mPVsfnJGK7qoK5b+dWrN/xcATdpyehyTWKHrMhGmfJwvDpLkB8FX0ryZMgB8Hb
crLlWQWmpi0rkyPr6IP+Zstq1zDvP70mr6irt7reWL/cLiLFlclJN5a3yfmDWx+c
WrdgYJduH+u8xF+TQ+ES8xgm5Tx2Q10ItX6oShaGa2hlz8LWw3eMcsfYO1aVgCA7
8ZpuYwtXn45GggvXkIxhyDKbPvluQVatdHmWwp+G28mTfVY+vvbKFMPRFhXR4ScH
hHrDbIn64pUO1AeEXFZHY9hzGUgCMzqg+QHPIHkaEmHe9EcwUEM9j8TIj6v30mGr
y6CbymOJpR8SqfKu6WWSevTzZDNUKGYw+XYG/O1Qk16MJh4OUOXwGSSfU22uoE9k
9dLJvhC98mYUHmV9F/G9D/9S7NNueqKat46IxIE6tEpCPTD/CoPC7zJ8x441vT3T
W5b8kdz1SofE6tPuimSVPj07EpHC7q3TWnYtd5Ccu+r1U7us2ziIKbVLaViIiz4P
B6zbL6zeWs9QmT1wQjdMWav6ysVrQBmuNAsGJqazefrndHNLdpr1AS4IMvJR24Nh
NGMxiCMJ2Du62KUxFo0N6eJXWgS5g6Pu/1efgBTjoRQg9QLaAHjn8J1coNcVQ4bD
bM66dHkfL2zY/eWBHnMegw8pNDT2n8qhvW5tqU0WGZLWe1o37AUJ5K2sTDveS4rt
KVGf2tJop0rE5Y6JIMzc8AB1uu3jqwBJU43NppjLCdaTGiGL1inBBW/dBbi5o7HL
5/d+aEGeYscEa1WEyF21JeQ7SotUOamYOg4H1K1fycenJIZB3Voi6Nbnwv7S+GMe
yszxyuTbDix5Zi31LpvHmW7o6UJT0otR5KZrbgdHCi8g9S3yNqjlcNcpx2RZZqLH
K1Cg+Ifa2I3mFPPZJWheT1BIJsOlhB2mqdJUypUGU1SbqOwjA0oa0iMCqTFlOMzW
q7PKqcnlNP7PL69k6GKp6QONMjbYX0fKtKgNlEO5fk/ivQaKcWLDHd2s5EPlNJzz
iBFB52cAM/wjm2FmA32j10C7UrMX5l16hQehINNdBJBRaUyfUPpyY7y9B65m70kk
2hvw2nevIX6D0NZiI8Xp8DlxZtf+6iChXnHF0Qwm23R14xHr4/OZf88LHlKZNZPP
IIofyhZszmiPpkp6rYkx2zwLGyiIMTFF84O/EUFpUHKwMLaCY+G8cPy3mxPM0qc2
cnuUwRAV0gRWQ+5EI+e7YidKPIVsnxI3//W5G1htRu7VqNeah5osMR2/QbAhpime
Hv6Q5tUqzXmWq+ty+kf2uz4pd3uvQLmGF0RkY5jNxhlBK206GMFzxieYXU8YRl+0
cdo2BYr3iuGsu+XxySWC5F+BQQtNpxAAV9gtUUNKsiMN5lsUlvMViDpSemnG8wZ3
SIT+pJ44W9Dt0cMZFtIBSyQCQ9zg/ppt7qAkbByZgtGBrxGSGjO7EHc6hgRHRtf+
4gCSgkB1gzZSLfDlGhrBpbLPrDTuZZHNsKo6qf7cCa9dxMz1B6mJDt8EwKk8IjWu
vFL2Or65IEoui/20oMbdPNBanDATyw4qNhDnUDst++s2/WUWl1hNVGPVuNiznfmg
Sw2UEYz9JzRR/o7Mw/5BGi/QhS5yRH47rsvd8ayjx4yHTVMUcx8KmHiniXnJo6g3
lv4C2V6r8zDf1zFKumCZYwmVWcmjIpkeCGa3tARV5r6LSmNPmPfikjApg3pPGQ9y
1YKD2A64yF3/X2EnsRFdpMbzUp/+KNlaumaBnpM+k+X+gkGkKCvN9yrDeNHxNwsA
aFs6OSGiDjnwJPBjLAeyV5VMONnV6S4Ni3ll/NGzyV31rWx/QvFNjoqLL8PQKn8b
xfYXOoHtgEs6IZy77PE7a9tgr77Qfxf6uI6OqIYS3tPMpQEp4pUqgxQcDWfSm/IG
0Hb4DMk+hlk4AexVP+ASWV6HWhAgNbM3PIHmZm09eCumm/bd9iBFVsmXr9Il+1O4
N1eaboXE7GZdlgl73NtHfNeZplS4CapRxK2vOpv2UTjmRRGbf8DWLiwT0X3jtC+p
Z1cLpl186OOZ6SLPTrJ9Z5W03P2To2TquUp1d6daOMRGLzNg475nwlMz3fEvZu+O
VWMcWvpyHpd4iBhdJU0dankrwLC10FFXnZugZpafBRqDJnD47a3XEDai1xQmXk48
LLyuqThCZhi7KkGgfrFHYQt1QQo+vcN4OTKrq9Mzb/WMdokM9hQCvpMxE8Yr090o
CNg63/tzgPqFDeyv8JD/ignG8b3QrisFrTqwWAwcBfAKyNEM+nOsS6OwNbcH74Kg
+f/DuAMvTT9QmAdbKkmBtc93n/OHQXokp7dtEF6jFhUcMGULt3k6o0olGsykUNLg
5p2xKpj+YwLFcu7bxotVYuQezowh9nRrtI/ihpawWPwsz9THodCeWUx5Zg58tZ4P
Y5GsEZkaDqq+SDnVnmpiqN2WEiuRv6++xrLUvgoBzPOJCliIqWqgQUkMRPgzTQtQ
5Cqus2kkMjAL4teji0kzfkFGNWn7APKz7kMKYe4fSBmTF2ew9tnI6HCKRwxb99P3
0DFLD4rXzOVjPE6O3RLvvwenIys89fqYTaemHDWYMAn+V8sfVWjrzewmMHn7HCqH
z8gKdkpHF4ySLQGiPmk+NtEbW6QPKcC+qdLdkDRYKbbPGvalHL4b2VWcH/ZsAoig
kxqxzAMIYpCqvSos6zcjOqBWsh2RzEACmn9T9HkLzRfjZdc4mmjlsridg8PSAvfC
Sy+Htqtn0koDR2G7gDTcm9UpN3voYt3ehm4X4LojfDqj0ArDivp1xEUIXoE+rcLZ
Re1f0Ok2nllDgb5wevgsZAFb8nge1xBnUt3RrgfpjHQAl1gewzrTfW78pD4kLECk
km49PMDGwf7prRSiNeFNWynTT7pziz57L29o4ATL2p0QezT3fxxPiam5ACtqP4vR
caLZmYJ6H6R91CLHIbSaN81po27/GNJ/duPNHswSRKvWZeysiyx/drSC4EpDNtEc
Iw6G9BKoHJtXpauF7NWbBrdOMx1jEFQZ78Oo9eVq7KbuHnLht/Iy8t9tDPf6DQze
JQtyarqlr66VLpO1b7CfqEev9tzwwGbHZPXoGIy+QP42opZQyXEjC0qS/NI0WukX
VXYHnlHdsRucfCtQ8TrJU/Ckgl7eQvm+DspzaSFnznb+zIaS6CIHk9vwLvK0JXzn
x1LdFz56gqsumr/zP15uYocH03GYbuhxl6Mg01Hg19bJrd7kBv+DrqL6nd60IGFc
itXW0innrqhc6wJvKR7taaYt/uu6T4KJfXlblNaQ5MqhfluloZjIclFvubF8lWLD
0k240mXq1662AxI82P/3bcharRBIeMB/TQ5hX6lR3tgImje27+NNJU5n66S1jEie
JIloKgpfsVw9EUYf7fHxftr4FojCzSDMcTgzpGiq2480a7rwqn3SS69czHRfcYfI
OdH8Cp5Somn5AFdajP2RMAxG+eqM0h8Hg93JDaQUeVxchCBc4QGy8v1fv5HzSe2E
rDK9eSx9lp3QLcMwWlWuRs9hvS95T4cI7ZFam8sUUOkfAnsG+6VEuMGH7Ig2/3mi
GYj/WgBkfXRodk8IQ5jPF5ZvNr9i9MrtrxG2KOrx8wZWqTsq6r6EGfe8sHhvWInG
4RUXanSrZnAdV3ED7SF7bL49eep5LBsfYP3tVL7zJsp8dfeofD3669ORXGDvciFn
/V1Q3IZAJBwOhbzy0j4CcPGUOh/mYejmAE1PRaquMfGKZff14xDrLGllvUmPiO8a
G1MkzuYJXl0ANo8nSDkBmgDjiGIrC8tCIxyFJH+Jl1BG3U7ah8qC8thAQlkMWzhp
+sbDtC/3VN7XFoHbxe55UDmS8pG3DU9hZpODEAzuXapGfA9mCZhF5WadYvdPDPGu
pBMdwTscK+KS5bIyGF5jg70zXEA+lCCwbPsFMsVyDZDyUFKsWRf+xwkzbRTN9/XX
labHnEki3ghQ0FT9oppMyYpLsP/G1Ea/bS9YylB87/WfC+xLfycGbwAIbrdJFfKs
q1kLYUY3pZTCvkZSR+bodhHWzS4H1x0E1eVTIMfhmoU/vEKu/Sqm1pTgsUZMF1Cz
giOlcBw6XG5pbaJVKrRXEumzjSvG/riZerGVogUsm5gm1VgrHUjBNg8sLDq+GFf6
Nf04JKpRX+WIp99OGrZVgQOgJkfH2/OzICOYlca4wQPcQm/y1/2zoSijeNTHOLI0
gbdwT6ZjcXV/wN6a+8PFi3WN6M7YfIdEDWaKEZxyZsYrDf7SoLf5nlkXwMZtt9V8
Jj9O314P+T9hzfPx4gHKh883wLXOq5anCsiTq/cTHdeiLdB8dv/LPUwtkuePvXJ+
6JC+xsXcYgqV8MyjA5ohVxXJcPHwt48O4Ix23oofproCf4V3LdjsMlFAZJiGNj2p
u73i4idX7m/EzP//iq267/bYAPXGNu/RB2/0/moTEVop0JtC8vHVaoSSsB/oBdnL
V1/cTtz49zv7MjUtMWl5TUdVMGZ15ctW+hU9U9mZvirBZ++ytWl9adZ0d4EK+dRD
zY8qfGv0bbLnA0Kg84udf2prwciluiqih8J53OqyhEk6+FKnlsE5oOx6nMJ9A0GH
Im5PlogfAro9clqOxG/cOPiPNRmHGi1vPPjuqN+QmG7cQiDDMd11QKGBot0jMxLr
pxD9t0Re0wG06U/LXqK3XNIjFT6aq6pu8cDmfUwF1hfxAqyEp2rDp6hBH6Q4MzVi
TQhwZh+XNSJ81XMfk9k4v1wW5euyv7Cb8HWyh2jhwnIal1hL0Yu3KqCp/A4qKIyg
rwWwvb6sR0hWbvMfBb9fugBcvsRw1j5wQID6DcXXJhHIfastRV9WefVvNWCpoF2k
mhFP+/KpMwm+TqQEeMNB720vYzKt7DqD9R3BBZ081hMBUGZe3HZdJquVxvOTlj+h
poYdzF1TFs5BfuoyB1MsFwCGcFsL6Z9x4vPZZTKjUT5wj96K2oLuTWVV6Mebi1Rw
hcdX4RQe7FCz0104u0MGSiy5hle5MVCtJdDZVeqJWOiq4PNOR0oQ/2ZVtqYPFP3z
UOTFMeCxqWnbhktFwqdrTyBE8vGN17eRtKO5nGZ9H+a4804GSU6aDUX9ZxL37+YX
mZqSWIrcb9k8RICCbFjOj/rEuJ8hWHDDitbsYZToz8UzxL5MmBvgVqI/tpKXDMMP
LX2mBP6m/bQyTid4IHD4GIHOZxvsQ3iMW8qeZiR+OBUxgMMSC5jCvXlzeGft3QQH
MrDM7/EAo2P+2NpRmMvbwygym1YGgLoUBOEcR8eIQceY5rmaKoA3K6GmBf1bwpe4
DPSnkLWHKpKlBrMU3wdGb8jLlk/qB10sDMZ9SMsq0ImcMEJGgOhKH1j9fcGWd5GX
wIWdMgenKFxc0nmZhEwzviNdcjRss4oC2yBRflSfGONApru3BKTU2hRdJdR/C7cY
C4qvPhDKGAgKBKqWTwChzYfSOyLUTQds3at3OLSePRnhrF4pGvC71wutzO3uAs05
8Rb+eMUY9jebSyLNobnuIrCrRvwd4ZLXv+NKP9FbV6wg5Ycal+9kfAOdskbpCw/e
8QbP81M3sdRqEYtnTtm3GxP3cYsXFFUocqmjBEJo/KU70FLLCwj5elYdGvzmhvek
oGsDMK9VwWeil25C7wNzwobQTa0naAlhuIaiHjJNP/TpUzIRd4w8nzOi4/9FGzpM
jeua/qEsaCsH73/iBcfqFvAuIpW15QAflHMlBOXs+Gtd6o+C0KPrsUGdU2eNWIzn
lC1NIfBQfIx/M0F/ziTxuVsh3SXvBOFgwXwLppWMUE8cPMAFZDXmtrch6u3oxnBb
OBy54/f2oDFogt/RKsUindxy5WTZ0lp3SfbAnSE8kQQY1ib9ixUef7XSEtG2GN99
yGVMt5VtwVfvqYudLfYWznj8oZtgWLbg2RqYaxOaSbpxZ8ZvPet27gCfJc9mPTI4
oDgtfVUhAzEKMQ0hb9KIoUytWeTGOzvXIfNgWA04xOHs1fPHB1qKNkvS5N5LtGDs
N8uvG38YLM4I4g8QT9DM+ALlotSNLfgcLFwC806i7H2HzuFq2TZ0KM4I+CJN3P2L
NAAloSEX5L2KmvtDmZAQiwnoIQPPnOCzJKmSBn7W5ZsBde24J3Qpc0YXY/zfyUzN
51RP9p8De96J222PJmAlDtXaT1IBodBBGsqtdcxvPls1kUJC8iyoU37LsQAPsbjp
SZ8pkEEPS9Eab34vjHOfk6kZRcdXCqtQFWa1aObi1Hg9tWk2oAZ5km0IbTCmM20v
DVU3Usxe9S9nTpNcxko/6TK9ZgVFgGbf1YBTdC90tLRTKfCx1KUzbRhSIVEFaCFx
9Zo5mOxKmT71mEXp29CnSViJ5ZqGT1gw3oWY/eGv/eFyZ7p5adWjUlrpkej+S+Ck
qMTHrtMhi8SuZn6OnISepJQJVyjTkKCtZsnRNCDiGIrZkjxKAyTUKri6iE3im6vL
W1XTk0iFe1mbDUnyKqj+MKdYD3ZGBhMXUD5zdk6a3ha8XX3EHIVqf3v7o44FIS6x
Fqu5F4y1Z32zSRywzaceIZXH/k0o59on9Me8B0LNmXQG6sBG0N9ay42uvr0Lduqj
mEPO388rX/ffMNLTnlM8cmEFWWjl9YIwNuNarQxvxAzAd13L2ah/FcDsesPkq7nF
AUQLQXmL4RyG23OPoXsZp10OHksF9yIyatp9UHOKvTPt8Hhaxd3YRlcia3g6EjmL
CU6sRdfgsDgXAkzsifsAjl9wBfCFOoMVZjRf5lbl5uuUHyeMd5fLkjUDs2ajHUhH
mvjCAIf1i6/dts+WJpg2lFDpAEW7ZQ2Oqddg9OtCohr7z5v9QK+ag1oYajyx86bW
2ecaQFToz48IQR+L9Jv7zPoAESEMolAUijGBVOwvPeIOyIGXhWlMaiouoWfP0V6p
uCGzmG7HghPHbBcXgECyt4C9CYllb2aBm1j6LRwDwqNaFzUEA9uhpxch7Y3Qvssz
E9dI6qUa2n6HeJVRkGZSo9pEyg52+TRZl52eIpKUP81p2HUlse+E6/qU9cKepnqn
s5RWZDSGwsz+IcX9GaI8C409SbQBytKAvn3APGylog2eYBq4YlUkDXH3J/q7XN1d
lplEdG9d6wYvU17DBS/IPpVe8cwFXCtZUqQ4xVzh/GBJiWP5TxuV8tSUvvJfntqd
rgPxGnUPbzXXV8qMvlCKpwBqRxLuxJpiCtu7sXZiIFr61RQ0kMLfg4nZakJjJx20
fjfoD71mmPRZDYwOhfguhqj2hTHEc/poE4UxRRZts/eWjRNWCu4iLWDJfWyNsMHV
8dxgNOMYoK83NBCp+4Tx9BlGEeJnPEKS/eMqhoCWoUWKtpsL3fnvciZtRQQofh2Z
t3EXjYOHgsc9sf9uM3MTBgM/1mKAMVpzj3JFTVSclKk8XFf7UY+JCsYy2DZEPVWL
LPnLrcggTRj1KarfZDWBcbIOc7lzuIKsciCSe4WMopQxL5crNU94ftSXT4yNbQkg
TBIWgwrxm5wFheDFficJTLqGoo5DEdIML6QKxv1I2z+F33iprynLOMJ9cdS9LDBO
OlIx/m64GqvEmVgWZ5+s04h2xEO1mv4LLpNdT+fUNqdbYGMAOVLACSvQlvS3FD4J
7EmPudzkuoV8c5K+xOftRfUx7mJxwtelaIH5FH8PIgxwXZzjmEF8WsdMJ8uqaSZw
nD72Hxu6iA+RkFgHu7X754vEdORrNMRNlaFk9BcNO2D6GNrIWRsn9TQmE+Sdw7me
x8rOr+AD9w/uAoHsQay/clEoac1Eac8zXktkp467g49vPEu8BzlTBafldXY9B6xV
qvooWTSb+XfbwzB/NBN5KS4mk5pZp3FY9fbV50k6jn0Jr//JiqpIXch7Uopop1my
YOxcSFlqmko1YkPg89yLryuSxQE06wc23hofWxhiKwBOOdtNVc3FqX8nNDSG0pJZ
gzgHUxSkloYqSb//cFgKvDxz6oQoDlxeXmnm0aDIBUSrVI6Uxis13cobZ46z6eZS
eAuX8/jtSo1F76I0pWxJW6rxYx4TGzFV5dM3L4i2SOU1MlybzNItGGIk8UC0a7nR
bnkpqzMoPWdLSZXRAzaPQtu0kBECYWx8WClXg0L8QzKjiKuns+K6j/foJ42yEZc6
qti4saTvWfcPF1D39zQvjXL9z3vfYlqrrnVNYWP0/31S3LoW5UOe405Ly4jOXssb
Mj38CRdfJo9q3LZ3ZLTEj4gPjLexcTGKK7a/5LjJwFXv9NLjyof6YHwh3EhGx8u6
2mYLJ1kv6+4dE2Ol5GTDPTgcvm+C1aqi0/2iOBvg1m9jsH46jZoOIObJ0FgM6Lsn
Jv3uEdmB7tfhgnwYtrXg4axZyyi/br2x+oX7pW3ywiGDiX2MylNfHdtjSomV9XjT
KIL4P5SXqlWJoYwC0rLLQOhUT2REFV5bMbXnG9q2JwO0h+gkwR41TBXjIUNytKHs
Q+65OjqfnHL0bF1wowFVbUlT0ME6rg4qTBfWLpyvQrFxz+te+HR/P2tjMhY2a5cs
Dq8l6IizVzLAqBk1RvCG/xkzDZgk1iYvqz3HFO8BvhObqnJz6MpH0bLsBBkeMTfD
kUiA4KzGQ3wnHSSMRnva252mRATq844Wthi1Soo/M761wLHC5HICm5Uy7Ka2x6NF
lGuSlVLWNfY2eU6YM1I4FtFlEbvzBtn8pOZZW094g28foJR0qCGxbAkBVEZJQJJu
O+lSPtnTq6PAAvxdeo8tMOQ92hWrbhGQhZwPH2ilp2FALm8uWqeE/fjioxikMtcs
/Unoz542RpstTVKCzIkzcOIfJ0OQwAyyfZ49ygynOSSS9XSlDtyMR5n14li7PILI
Vd/7+MS6YxKg6+Jn8MiuMqvCr5JHNXT4giXoOcLGMiPefvB8zhXMy7MDglqFX0AL
yvI94J2fBntkhj0mmjgQX0Gn4pHLY38+y+5ZELANgpL/r9AeInpwR+EnOfa4M4Ys
BcwLPcI7iHGFmrsXEfYANkV6aGb1esS8bF40XtmPqnE+Al4Tqd4RMh3dEBmfwVyC
oLyatJaoP+H5ckr+h9r9k/TdZUPSeiv0QmIoN+fvELg7PExae6FPjemRsjfc0/V3
xVXlj4J5Ze6XdwFRizPiPgcUTDNIFKvyE/RdqHaFMigjGTg6yqMixSICDRZ+bT88
/jDZ79i0vlEovyNhXXLFF1+TXKD5zHjf5kl7ppQNGIpBPT3quV311z/d+oVkSc9u
PxyS+MDuYD5ipv7rFpfy99sRNbCZxvcNiD14icNuqPMiSMp9uQDcDdqA5dmMnyiq
MmyKmuwwV34uCl5C9CQ9W7vfiE5cURlvk5XbFdIEV9SM/biEc5kCCBdYTiQREOyc
MnUcKfrRVA6z1nKjer1Sb8v6Pw3/w+Dbx6sbBhqWGoy8DAka7y1NjVtQwSfrqo9R
As7hk95STyymY4YZodGPXMBXVeo4MHx9pV+Idmj/U/A26lgDiAf/q15d+lbMhK03
EioozTElwg5cmh7FMm6QY7B3YsDYi1vtgNEfX2gbifrU3/B8QkiaTm1QrcyX7wSM
W1MciAM/v9RtfcUzD8YbpFUVEh22fFjobThL+EZz9w3zuSlCDNRFshqSuUT/kMFX
lbw76bSJJzw/lH1d4/3gT1jdIyHOYoWuR+9zz6bI4DfOm9XB1aIg9LHeTkZBygcR
00kNSH+CajMbmPqP+EShFVRPeCwawbB0fs8OmGj/JS6Poaed2uBognC5VHIgRnxW
Gq6pCe3uqWZpgCsHYM3QKyDTRCbQ5BgOKTKOWIaGT6USfwZXtYMlTceW+unf7p8C
RKgAGVgnD/hRE78Q/mlVkXEIeV1QHnrvOVD9zuNQIqub8niM6DeHfrJA8Qbp1BgM
PWsEVSRHI4f8b/PinAWNEEdUQffCx1LA/hheQyiNfYMUDLMZLtiKTktxR6gGn1Ec
vvcLYMnbRfMwg3dqvTDRoS2xlsLDWNdLwCjU17vdWKaFduNTi2hiqOtR6FvFwl8m
TeWQ5BlVU3iQc72MJs65ZSyE6WdGA9dGeisfgywegKqKUAXvJ1ajiIgX4utPuyeU
KmLrWN3q572ukNac9AwF1T7r3QBgCBidvwqRTL3MPoieDJB2EkfTAm1HORlsXOBf
S1w+MB8F8MjH0HkfOwQnu/Jo2Ab+p6UV0eXkVijO6qHu4DDpZG42OTl5cgwndYcC
0rFUTq4lETtY8FG2TilSye3/Ly/WZRizAsVB5Y3h8Q3E4y7ARe/2E63slBQOFmz6
95FTXSGY9HPCWqSIJRbDAbwNIW/1fJPryFVwmjgtBL16SIZtYiqaLEDLm47szCH9
tUPkRTuSeP5Vz1gw9Mmp1yLSh19zyyh5uL5HsSIUPX3SY1mohKZcQ2t2LZlj3vGx
Bd3Bwuw6JAQhrNA+3q+/SuyU5znlUBg+LxoPRdA4NKr1AOHo0PECwbOftRD9v5tA
L6pOqY0k95nTLpkT8wiD+30WnoDdrS1MSmZJX3GuGBqWbJhckpODQVeBPjRk9TmS
XDIPWcSKtf4J0e3nxpws1cjBs9MV3PGhu8Yxf2ySLvdnAHY9lReKKgWDv5CzwkWk
wMgT+FMzoKnMOYQhQe2Q+ZSwOod1HnKLIm2AbLaUH+h0e+5iiOQEWLwDXn6LuaXc
ctiZ/PAk0EFJkJg+pefcNnBB5lVcW4slBrpcXPJC+abTNsOpomtaYEjdSyVQYoyF
9pilSH+QVnR4qQtTB0axM54BvHN0UErnnSQ3G4NtSz0h/kV2uAXzFbi6sc77ykty
CdUUj5IJT1TKwlbKlR+dGFUuzeQjjyhiBU3HWR6fj91fgauLeoP7V/cxYxvkaxFV
H4FuaLZ8gyGhKmxuWD1/8k0A6v82rHYrlSHkjI9H8Q1X6VFQXFJJCgmeL3Mxihrt
weZfqhbXxQlRU8MXMNusg8c/lSHWJRQG3DpCiXwpihd6xvkFG7bKf6Spqc4IRHbo
20UpDwhvYLTWSDL88vlPakMy7XGRX8BO1A8sxQAOOFLOrzf85vwzSZYFe2I3n4kD
T/dWY4qtd9PWbe8UI3S6akcyq9pQuCZX73y9RDhqsxn4987n9KJWH6knCeB/RGnO
bOSq/t/pppvNeZ76GLIEHpFHJ3dJD2zsQRpI0CqM2W85WVYzO7TRAtaMFnP6lohM
WsYHEp9I5j+SCGOcXWHxZPtwqg5njpjiVD3+ERbM5sk/4V1CC+Ob54eXQRpXSUXV
2LCg3aZ2Wl4l0mOV26ye+0O9Elv/rSjZBpmQO06XpRCrYkWI2RE+tvx+ihzBfrAi
3c3dFA4uQ02OKE4AVfZc4f+soIToAC++M/N9zV89LjhD+dVDhAHNDm540OZmgkzH
5KaepzueXIvwzQXSYPn7RNDqMkQLhvZpqOhpzVhFNccAZ8ssKxrT4EaOCisKAxO5
LhXSxI1MShomKr3sQmk3lXoAsVCbKuXqClTgGXAJJktoZRElAGPqqpZoC9dsdQLh
MpQlU9nAaUL9h8Hy5RyLw7Pn2FOBDuV/NSpnI/y1Pw8mfJczgAnbfPlPW4V8Gbj0
n4XRNZ6cYxHpR/eVRplLgAQVu+SXTaF3Iwy7+ql/kBCxezg7LKe85Ve4UlTh4UzF
zAhQD3aJl0Yo7p/+nTphL9JeewvqO8QKH0R8dFqmpyaF5Qb0XgXMAoCr5ZoVTigh
vfBT+uCNbvi22LA6tpk+TFUNBJLHduyDt65KQQQqw1PPWCI+24kCITlykVQsVQ1Y
4pXdRokmxWJe0Od1a/KPCR5NdZy4YtQqJrZa9UHU35JP5UUa1//ZGq3rbJxJAZh7
m55WC8linp9CMIS+yLIckcHL8KQhKVHs09gAM9ZkWgTPFpf87IrOx4py82GN8eHV
pldZ+oMWRKn+zgHhGZPN2icX7uenbTTvQwQSnd8p4RMo6NwejHRAYDZK/PPU2jT0
Y9p7YBpXcVzS4DQg6Xe5fZfGsi9xvIn0EwmsGJyZlazWkPuCw4B2GmFBiuuwiWD7
qFj+Zx4pkEV1SN1xbZbM5WvNAQDNZS0Yz3k5T1bzhjxv0TYYk8VnHyos359HZEYN
Kfffc54dkpHVwAoxHMumAMFiytMSagvp1AoAO2/OThtrkZ78hPJc1Ui4KVk7thGf
ZzIdHpUfqC87GRzXn93DL1l7132/O+7zeLyBV71EJS3ItXaFSVJ5CoTWsnjhYw+L
f+c2UmLDFxewcWxeBNdjYrJMn+4ZfAMg8Y6fh3+RGWYasKaqzpSXjm+u3sQdtjrC
5FaBQ6Gh0OWh+/fU5ceWIm8eQF6j/+5xAPDpswrwfilKfL3RePKTs6qwoU8YO/1D
coqAZx6Peaf2UPU2SdlzlOZz4yZxUWLol5GaLf104ncO3nmsiEXu8lzzDVV3kjmg
VD2OjHw+yTYRN4O0OJyTI8J6//Cgq18Kq8EaXrcU+iuChCrsTp1s21yTO9otoEQT
G+W/qpshA2E/as9DcYynodpB1w2YAMIfzkG9R/it1LfjMbN+aqetoOOyY3wqk2Ue
WjktHfirQGAJdLcAHgmas+XEyz2G3vBPmi1MViiujy6YD2MJZJGFkN3uYIaaCYqa
EDmpa99A0pUDH9xJ1jytSVGxro+MZCCcyOa7E56RKiEh4Z5eyv5lzDyBJjjDyBKR
4vOigp25MojBDm1gmNQstbnUuYWOWGMJicTSRzcoGonM2ScwcbGhwpaH+gFWh6dm
YFRB1M1qQYiqzlZElquiihHSenYgBY531o8C4B5kSH1QWHQreyQwRGRnmPu5qrCV
EfNSKEuaaePGzTL4KuUSeiqtepAILJVKe+2K8roWxDR8UHCUhVWGz6W97p29VBsQ
yyr+3K8J796S0urJZYVJdmguJfuPpUB1nj9nKykh/87Bd2Inuc4Tkou0junBwj/q
o/0AyOOcLdNpMYSPoWSAy+qeH6SDK5ozKIsuowSg418347ZYcFsKMel9yXA3Vbt8
hYxoFkQ1OCalCeZ/eOJylFoq4vLArlp/KXjgPaGMOkARB5A9ipJ66vTECHiqKf0S
yMXWEwqRBXQJz1nDmpsFbYdAJ6lMBnKoZiAbaOvUNnvb+YTbHmxYyvP8tx6lz6A4
TdGKS3hPukfxge0Fz78cXWF+D0I+FxvJyoGrcnNyWS5W8Fbpxu+0n1IENn6S2J5n
s2om/PCC9b+i9MGwUJc/DWDkZLUmiQ65Yo8/YUizt3ClbUXjwUfJVQSCdJshmOre
yvezEpfmvi0rV1nRUwtG3Jri6q3yF1en/J4dxTB3WOTKxNntzjIyiMHsVTMu+LxT
rrl9ZhMK80bJTt5hbLIB6pXlYAuHfMJ9odJ8WPmOMIAYevsZ2maiwhz3pUszEPKQ
kMLwVE3VGeEvrCCh0a8WPWBC4yLD6uJApvUgadGvb6tcYvAEV2fFasLvxz5HECs7
9E0VB4pIm0jg/J2FN8PXvJsmHUbWhph4ZK5r2UMqEX85LY3a9/TtYaKge4IkQqCe
GFrR3PV76dPNcEPN8/+fn9r3VaBGinkcni3QClXRd0U9z7UuWwhwAn1Ahj7LkoM+
NGJFl3NaVT9OKd8VamMjI1SOf2zRz2MIjL3/BxBIHK53pMhehFrGvR1o0CjyEBpI
FeOC9cdpp5HgIlQhODYy+34NB6y43TqesGrNmdqjGNkG4w6hMZHNrLduWqlsJPaX
GmLn0NQL47yfF4ZTSEIT/wi8uaMc59jfWNvkEqs50jQG+Ut9fsTG+zPC+k6Au4Zy
2FG0uaNb/F8ugX1NL1nnOcy1UMxoR3w0Ynd8D3I0z3dlJjqcXMTkSgmOGo4nFGJY
YgJFqdV5edgZIPHuXWV3e7pwUtUHgaXFFvduCUUR9A+F0fQ4BXruYEEgVsYc8lvU
tDggUwOjht4STqBBHo4TMEe1yci7t5N++XIBqavILvxgB6q8uaPO42v2QHx/vBRE
fmR4ep/UAi4S6GivdHgVo06OKbq2I2UWyuL/RuVee3150qn2SoYaP6Y0yQ02yEix
job4wGyl9nKuvC6o9daxcnwqJ6q4qJvyqVYQPyk6VslvkV9KKedhOVMo5ZPSwlKR
l2vpCuUICzX03SM6uBQ34uGV+pdYkSXZxG1Jou9HeQp6jA16r22l/DDOLMoOZFF1
npHX/30D/fC/aakOXlnO2IJBzOfczy2gRbwYrRaAxoayecviP5ZMh44VZSE5OytM
qmWpatPbl4D9wD5BSYSXsdKPVaUqHvXYcrJNwheHmLjPn0HW/tK69A6uPgyXRYaK
CqLJ2GjNOuz66n4hi+Z/8/5LHl+8ZuuPIDh6SXdo5mBBuNyz8E1M2q9j3S5yY5ko
iq9WX4u6u45hUVrV/k1cTKxHR3/Ako/dtm7wo/msYt8YovbmrPoV3gYj3Htve+/s
+6bFNgiAnBXl/uKwKuojzOS83dwqL2SvyISJm9+ZItIyCj7r+FMpUxyX1C0Ud/cK
GzfaAE4oP5ROXpFPfsmgEX4tehDn3VERUfieC+Up0l+k56fnEs7iqoX1p7tqgEz0
hCYv2KoY1PPs2uPLZ0OskMvrILTLXYHwX54HPbWpmzvmjZdHpfw0UpLAQDlsxh3O
RXdCQiumJS6UUlSG4VDz0ZU9vfMb/MGGcX7Iw0uL+FLZw4BegX7N1mCANuzacG8U
bHk3UO0GGKiJx1k9bBmmh3cYf3jXgBCAEsXNfyj+iyfynWB/Mz5ANN5Lh3U1QwoS
JppMGRiIMVBqih88deKe5194X7aKBp8oZLeqaHtwj+MfnsF2CJ62q58M8TpQ/Ub5
yXEL51aXR73noRHt+jzJqH3XsGDMfgE8T5VnwlIh/QLBpG9VdpoJbUrhYsP1W9AO
ZVb+FA5+Yyi8fB8Sb+7STYn5pg1smWfT8Uz0NPBbtnbDzdv3DPojzWCe6YcaQsCV
pKkcRwPVgebpFSUPuEgp+QM+qk5NfEkCn1MLuMZNlFtmGUa5Lck3m6PweTMZzZdH
dMuECZYBBoGFZJb+tCg0++She5e4HG9udL4DKEBKwHJQdsHaQezbsmF0zoOTYbar
xdGuo6dY8gpzylcnFDU6mkxsK3P3jGivzUBJo+TOhBYSbW64vAvHRNoahpVHXBrN
dJahhXy79CnceDArQigo9c7QbTndVkaQ9b9+fG2O+lKClcSlU94d0YQuWdgUg6kR
XsjQ+mhb9jhYiAS8mVnSDFEI1ESLKueA28BpV64XNJ16v8TI5Q4qX4Y8TCE+TuhC
nigNCNYfEFm+kdxGS6W/KBH2CVnYpH50jT9K5eKphgrAvNKHtc0ErT/1O5NVz3ie
2WYvBiyiG3XPy7FNYzi3B4wdfnDrjaD75ddBVRhXJLBRdQAt3GoKxTK6Hj0NHMjW
5l/PS4ZvXGSLEX4AspdZfXZFlJQqYZR3NhqINqdsaCBmaK9X21CEF3XXztHsuu/I
J67WeIyXS01B3B9SE+28DNwdBwIIRKd5TA9uauDufJbVoq7mthoZC82Vaw1XWIex
EG6CbIrQITASKE0sWWmrLIk/PsbsxfFTGOh+mhKQ5UHgW5pzREC/FhB2tvjU7YKv
hNJq5N4PbikfDbrINkkLsNTudQRIAri0JAVIDzIckwwJqdZBCXq6BuGQA3JXVIEQ
IOlt0SmdfFFcWLXc+GJ4YgWRDe4FxTfMYvvBNmLT2zRZllyZ3npgHFy9iVRUuRoC
llEZuETXB9t0IDkFGY3IF5M6eYgLGuxS3axEloe67opJWfenMHLrBo6/AK3mOa9P
3n3scgY4CbRlh5sbDB6xmI0rH5m7xUT3RpJ/+abVhmsQ/YaezQ/CYGZyQQ7tW7ZN
qOrll9M3QWH2SufSuOCfUvynb5O4nh7cMosg3NHIlX3HxWxImQ3v8/M2T1hvdMv+
dty4S8bSD6fIJfY0Q+wWA72oZgo3WkvjK+FTpixajG5xcLmi+kwsPwOOshLzxa+C
ppp8hXZXlsZn/7hErv3AiEWnNgCayIBnJZM2FoO/CSZ/g8n1jEqR3RT6vjm+qEms
qvYSQgiPK8VmsSUWNErosdSYRM9a//AGYdwLSWShe3TYzQFKLR5iSqUM3WeFc5Qk
mOG/Ic6iqJMZRup2BjJHLGmsz3LGRwU5yaBJQEYNUvkzHWQ2Pf5FiYvZP0l3GiQj
T96RpQoAUqWCp0cgWXAUSNLqJi3REQNO9a2puSLshTajFlEz6XuH30jc3pq/qzUk
6Tb0tlMIB2xQE9pZVyEmL0t1M3NvoOmmi64Vzd8VUtBlQBbXWF02VlE0Qh3p1kBW
31RhsqDK1/cDm3mJAGGx+5GeFDif+K9SbetkmkDjJiAywuN+kYMT3EX8v4JcdDnn
ccis1aJlicHkoCR8Xnv5hnYTj09sUvwYL+9wGzFBOMmyajIng0dT5ptK62NrbX5R
oojnJCI2kHVOztk34GpjgFdidEtX8wLZ6b3UwuCvWyHcKyJr+sUVhQyvdQplFpsk
JvIFmIl7u1K6jJhmDGpuFwyArlsWvs9uAzQVJMGCWHCgwQ8m6lM9X5CzpeqpAQiT
39otbZqhInkeS4nhWWIIoP1Obco2y3ApVHQFSdGfUK6Z25LGSZkxD3QhJXJw/aqc
aOWO4XL9nJNOX0VjDDUgiJf8EnsC0AzX/r0mBSI9VtTyVcwoJ4Sq8hJMtR+Cg6Gp
nLBhMkf6CIMBzgb/Ukgd8KlcC3xuS4lKhIm5oEK6qS8SBctVSg3JELELrx7kTWKX
RhkiYD199Ox7a/N37q7iFEn2Xv2F2KFycL5/NLcueuWwE6xIcAWephB9lzNuPzXs
tWk3oqJqlXZJT4kf1QwrM65ymby2/K4vxWR2Yf2oRaFL4A/ub+2S25UW3i4Da7lL
ckp/PlaOGy7OzKesErza1yiA9RP1Ap2tHEVjJ0FlDaezqrtlSYh0sJvsijL+Bvr1
1v/nZPVZJW9MYG9rxXCpQuTRVBPwC3aFgb4yapXLz7xViAb4w5mLDayNLr3YTR/A
3uvcZoBTiuY+KlZX/fjxDelSL1UW4w0nm9kLC75Ws9znqKeG8TNm12HyegX68L1b
EHIx8tI1YPqYOIpRemOe/nAWBYqaiBDMD5chf61Oq/86Y1r1QdUSBrIeTtyCw0OE
fok5Gy/NxuHAiYjC99rBMvMcB1Nr16R5r9v9qF3Me8UGplnmTwqGbOBvn4B8CRbv
1gVHzeRjFw3QFE2/haOr10kwie/n1vWsQUIGJkIk1yqIOlNT6dqFukpwOzzdqZTk
rWCw+3wRRNSrIwelI9xUvFdUIWYmz3CHP1Nua41pXEKMDFYFr+5jQ+WWPqfoj1aw
haDRUJrPD6cNVxzSIps1alsgE9idQ7ZrSF3Uhv2HGU8IdP7cUSIRZay3i02ldUM8
qt6zDaonc1jM5bgM9Y6eqmSO7qDLOh3RR3UahuWBRR67KMgF0KUNuyyZwGh+qR+y
lOiQXIBGdGjK9KFHDstkYmRnhJMf+MEAczcRBRJJqXAIX2RJwBMEME1xrLGH8fSp
OkVZueaYkXHCCMRoofJlu5+TYVQSG+MPPxUTxTikgkcDhj1dcf+fCDkHihmCUe90
WqpArqy1nWs4gHjdbJFdyPgd7wEBrNLsMzD/HpblwQnac3+U32Hn+q4KQdi9EsAw
6RVmzRU4QhS1XmYv4CvIxzfpApWqpkP8ZMEOl0iGRefpunChIVotLqZuvmBYBBEb
t+nsAIYOL9KVegTL5xHb4JWHUGhb9vdMRvFnz783nznrunSxDScf31l+bPGxTIai
BQL8t+ci13JLR4O/3BlwECj9TBTVaamhmCTBy/566I8HYv1gjDaiK0XKdf7zkZFC
S0D+TYSO3nd/uUH/jl/yTjGej1wYiuAkf+4ulUoZxjv7GRwT6auFCTu6G9TvK9o4
GWt+IZJjTLva47wbezw3bFrNB0Vobuub3qz6WiQEEJDrDvcHzgQKldV+b/0HkBx7
SdHgrdlt/q1kXXGh+qTieHXXJIzlCQVS1sGtJIgolOADVTlIw6ebeUnQeGiCZ2iQ
V3VLsFwM4GveNPJXDRxRqKeB9VJ6gBxFWNGw/ayIEjjShgdjaywHbGSFgiMMOcMr
84sYir11lFAgf430Xjf6hLS/3/0FPD18T13wELVzA2yl//13g1T02sOn/0uPUuD1
8ZreiD57WpiE+iZ8Ybwh/G+2TcKcOWGi4hHVp+O+88lt2OuoDK2WnIb+HezA7eWr
BP557wy2/uDSnpITpthaRAmm/46/duIJgZKUG6pP737m/fRgP9NjK7+hCZx/925I
DWJYbROy/Dqmdq6FeZ4sWK3yufOIqRrAiFJ9OqS+YUB494ZMdVho/QtBobxuD04O
Ft0kuxjo6U9MtcTnmFqc9+sKF6/92QHcKnTS8z8pUENwOKoJ47EoiFSuP0A91Qoo
BKsSKHyE+HOegEZigX8IxcOFVbu0QXeR2tAepKwKaMP6wqqHYfCeH/KAqsyqwr+4
eCF9jUIw8SRv6TDofOqnTkCdFOykp3dJcEH8slB/RoucC66yXVTx6bUFRxns2qGk
b58vunRvz5oApPYx7eLrddKtM8YBDNLgNhAtWe0BQWZjxyhXvXdByEaKOns9QCpU
zNdI8y7y63ejevf22if6fwp27zwkGB2l3YR86J5D6tIJ2+kW02LX2G837rwGymCP
WdPK1rvArzuX/M6L+H5aHv8l7zLxVnvSIX5irDhrgiGYgL56mkoqxpelQqT0iBF/
5CW/0llc0EOdTNWj9390ccetDULEJP2DZtcbTCeg+HT5tp66olnrsPFAe4e5csmF
CwWEQQw6CxYuHPflrndMoMfDZIQckTH12K6dd9FSj7haJw2dAV5SmaUGk3uzH2Qt
mTlyhKWpyWZKaI38pFQC7WQhOXN/qzJP+su83TQlk5y5fT+EQqZRaszyvJUEq72w
Slu7FCkQ44cEfC7HfFKy629Oj7rC6ncgr0J9e0hgAUD94CY/FDHcHCssDZOXiGPY
gDAfEGMmjtjw/Rnzky1lXibMNO0eA75THnaspDIS9s0FqT2E7hq9OtTzqcX3PCJx
lXvc91JqDFB9MY05qCxAkn/aQOOiG26JuabJ/9+tJNNRq2B9pNX8RlStI2L2IB5w
CRtZZ7H6/dT2llcwl4xW+I1VssY5z/mLicoh/vRc0oSAvneERPGRmzOyBmwNQA+b
nloFTdZEWUcx65jQI+Lci2hIOMtC/tQFEXtBS3DLV1NNib41TFB6qcDcFswFSIkc
zHAICm+uuKuZyIp1U+Uwby8vNZRGsHB5SEmoK+G1qNyQ7YecqOD8LQW8+ZOon+DG
bSrRc5/02GmHMhQG0zik5rqch0AMlgKde49Y5DR7BRZXvIH6Qp0YpHw14szq/PXG
5LScUOCeOmmVyCPlgetybch7toZ5lRhYoWxA2ImLny8JMYyTA1abAIiZq3PSLSlY
6x/9U6+LBLpHcxqY6C9TLRCElcsah0NzKcpIBKTYOryLJ+xk0b9/V704fLIh6ARZ
nPfk17ojRP5t7ZcHFk1vznj568n2ls2SNF67ikiwxLfoORCLNmNTwQJfI2nuH7AM
Nd90WWnlYCFdEOVS2Y+4RSINA4IsjaKeNTtxFPd5cR0oqaUs04Bec2khikA56KJU
xaD6R6JuIZetq0LXJO4jrA+8iVbABc340r467uMJ42eWhaM8gF3kGFaZslhLUD2m
y0kz20V/lbc4hO1tJN91UUL9LhPiHXlmihsvjJXKHpS6OWu13faN7PpEGeU5sLNM
nHy3jxOv6532e7gvIr//W6pr/ACXI7GOwvfn7eMG/dR2NanoG/RB/yKRAHpJf1Zi
Q0FSfV3Q8sgjsNZJZnc0Lrpa0lce0vwT8T2n/4Tpb6vLjNhGV9OpWra+JrJZ9w3p
/9z86wNGPCJVad6quFUYcFD9TA9PKTOXk7L/2aio/xpl36ONRtjuzu7iZEoPjONA
RBvYdZSEWcEVz5C+VxSYr0r505pXtQkbhLZ9xOSSuA9iP9PS8m13if10CvsrXVHJ
RnoE4lqficSs8ZGAuIF9ltCYIHKfcx2r46aOlZDRED0Z+0Vc8WCHQVrJ/cfS7NFD
6f+OXLjIQezwYQVK/2wxnS+10RgiH/4QJp0qrmDafPJtuyzWdw2dxXPS8OI3L78L
Zxbwe2OUaEz5kLOq92+RxjPnFDnFUeP2K5EDft5yD94hKplfSnEYf4I9E+OuONtO
zDxbLcMx2UDeqfNkdpxvwEBUZMFu5ZcofApiQGoZyTy6PIJiu0M+8hwHMkKKatEw
KZyzEt9MqNOO/3LEYnTGf4cbZuSEGQxtlDn5682uExTeNW8ayhemPlTk3ypqQu0t
C+1rYZm37z9MoP5o/EWsBKKaf+Yr1c9TChgGk6aA1z/7Fd6x6ZYyp8noji+8UTaS
Ab763zOtZT6ZYDwWOL7HttnlFjDZukUQhHmFbGz7r9rxy0noI1vm961ueQNa6ITL
YeCrOdPKC/Hdg8KEPSEWwovMIbAVud3CVmjgQMC1I443hB5erS9899ydjatYF0s4
TPLl6KOUaUpQVotOruK231vp6NjJ2fpfQwI2WbgZHxRmcKY0YZrA1xsmtEYnxvKz
umBNwzzU+PT1a/GLAh/Cfoi+/uSNSRtpLxuzZtmVl5UrsRsAPvLFovSRXQ7Sj4dH
q8UR+k4aqrn2T9ZLf4XNqScJkSSVUyIJjuYJBCKAb/WvVd+5iRPVHwePnoGk+2sY
hGqLkugrd8acfGYFzGEN0Xdw5daD32ysMgzNX9tz9juutozgJjc4ssLPMt6p+ZXx
Gias+eJ8zaSNS/A9v47lY2WT/t1VKSFQKcLfeIJ1dqW8vTYY5sUmajShmsYBkbmG
BztdW84RPEDKk7yjdDceHoAk57enamWTQBDOjo139WZ0xaWRB0b2SOGprHw9kICz
QjMBUSUfXub8ioEl3OG5aYTGuUK4r9F2ZAWcjula6JUOPhlPVz0jJ3UWPk4j4zhj
vK0BG5LSdT7IkEBVF3gtcV41HbTBhv9n0ah3tfoJeG9sD6x6dICwGP0YjgMSWluw
FDL8UeX/2sYCkr+7yei0VnINNM9DULaNiaZcW5iMiYeo2LDlFXHOgsvat65Lt+F9
smx94JhRJnC6+aw+/MAYEG9LozrIq2Nc++I/nSPvQnCvQ8EUaFN/pjVVUf4BQYBM
HlK4+JHVZU2o0kY9GXh6XXFaZP2SDcl2NicbQmJ+zu9XnAQJOTnfn4cVF6JRTdfe
KuRRtAfy2DTu5GcZHr4e5kP1KsBPP3FSoB9LrW8arFpSa2nGGzhmTiKR7Md9cXMX
LbnNpjB/Ltde5WYKTATFl3TqSgEc9qxEY/ADdfMeFSx8Q3Q1hHswRyeGK60kAVEt
4u/r+DoqgNicELsQXVmnennlbTu8Nya9nGLOeSWcfJ7plM7QIOFl8ZvTngOv9FDj
btb839+ovK950C3gynPIcNUEycU/NhGqPrkC93zVPdDNKGqFK4dpy0Ru4f63txT1
1F7dHDfqDvEvP2mNprXfyxC4lVbnTZtRG2gKDEEAlsIoPhej/Jx87/S2BrNitD5L
FRLZoZCEhamvQCsa0xddt/AVDkiFqIsw8Ae1H6AixjUgedIYIpdlCF5BdfGdurSi
CVOuvj7T3sP+1O/qUaF+sKasFtYqA23q5Q9VGcpwBg+RKz2lGO/+TwJ5xKE955Uy
uWQjxPjFUnyhCTQ1GJPmvop59b4PJMOKcO9XN8sLLJ4FoHCagu1uAafXyNMXiO10
PmUax9Vu7vr6T5XeCHotSs6S5CpI9fIywypSj17eMM76hE9TGwmzklitSu6NeNhU
HfMT4ucBEoLSrVyjjSQah/eWnruon0FK+Yw9urtdyF18UCHulJ08fcIXJguS+kLt
OA2XmmfCRbtfTKc/kdMMTdwMJdXTK/EE6S/j15R5Rk3HdjhrSWZ8eBOD8oR1KueD
U5MC19nlsBvrSqXy8XXleDwGukKxyD0pUH4uSZq5zoE6KWYJ3srbzbEokdgNxwQd
0TWb5ZCZfCXrbZz6lB/r5ITzpjw+puXuJymXUFt+brgTJKPUZai5SmCTi9XNnIRS
BkT9fahLN93CDix7u2RAS80Bgktm5MBNelyh3hnzlXoZDwCPP4AzQS9KeCKhrXoP
GkkMGnYUjgj/QjgUjmXP+Qg+s20QVPVmPgTZVbo9tm+SgyW9E5QPmyrzWqp7750I
unwIzl8PD1IOzZ8WwwfmJ3pJBQcnqebB3nzjDthzrw7Q0GalVkgBjKL4V1U58+Mg
NsNKUgbaj2jA45nN2Ckptonk3gYyi0/rSjyqSDwrYV27Dn0Cjq9Ob8esi1zXU+lw
Z0hlSolqsPZciu9QqalWuh5PbXm5bupc/jiVIImNI5Pwg6dwARQCPptuK38dbe4y
FBX7p/SjUcRJNubW9xu9X2Nv9CeCUuiSbLXSpK0uq6rADWRQR7rNyQrdlxJ++m6P
qV1KJl7F+xs+Npc52S7sSet5SG4fh2nWT4nAPs8GksX+eJfwAmIBnS3GutZWFmH3
16S9y1jxC1J3HCaP1Ws29s3nqYaApK4Qz8D/gTshkibTNiQ93ZEgofdXVDPCkqAg
geYpxFpkiMFooAe/16nY5IK8H4UHCgKeVtq1gYKXQBNLnHofmjcYGr/YSzDn08hK
e/ghd7HQ8wAxrxm32exvFUhRg+32FXCUqLZqWstVXbRf0WgVRSWGAmKHdwDZJxnC
7yfs0bwwgHTXt6abnF1+m5KXe2LACXO6qqfqQvK3/LQquH9HtifjC4MD/DGuwNJ3
dIYoO8s90EiKQuaWmoJ8lUFL7BPE0MaTBkQTca26rDYzcUz3PLx2tjRKPAzJxtkM
FzxbgLwF7L4kctqE8EI8bA1fcOxcQPQ3loXBdSqfbZDqSmNcDCcA/f72Ox6+fhiK
zLyIB4AcOixqVcVkNeM0u2VoYEXLKwWNfvBlPuCWSCUoLRJ0MuYH7z5aHt5iUQeI
q/28LHMF3gPRwqJnvmmGywI08m9i7cvYPDjGTqiF6eLSZ5keuEwZOh4F6Q9OzYdm
5+RLutsIkBJH8MbkXuSnBJwJSSHuKI+2tkHoDEwGpJMSSyPndKiABvRTFn0EnrQI
uTfG1O5pVdFr6rbhw91tU4a5wgcBhCTQmOSejWMPQfC9QB4ufbAmL81zziUN344a
4j/24St9CEVP8GOSJdFd7P9IYQWfVG+5aprChrlmNr0xaL0xpIxVV3tZVu02mioE
AFWZ3aBJV/0iGS7TOM1z/Nm+ru/ay1SRpRmwB598h+3+qRpmske676fESIlHnBSu
j63d1QAEcOqvbuCaw143Fb9cIYI0ajw2sM9NLrIbKf+KnkGZqG99G447Z+StdznE
vt3AkMMybSM+5qvGFE5bTrS3oCdfqkJbJ8h3U1r9BX3yb9RgtrdtbdA8eYN4RNID
8fenovL8B1Ooww62ifZbzxsh2PYG2Vf/i9QNmTlCHfmu6lW7+VybEhRln3VHy6XL
1OJ+E0yvLuvKdCG+NOaXMaNbxEzVB2O2emDwDmyUSFGd6vbLufmqF+HHPZLa9Xj9
etUh54YzfX8TGiH9ZKpYCrBMl+3sGCS2tQc60gqHVlPOxF//apuemRQzosB5a/8b
iOcoNtHzGvVLLXSLmsSS71zUo7TDNOnI6F9sAPZfqbXVRbM9XP3vBYiZFdwRaEUC
T0W+dzfP50KSjVXzFLKjMUu+WyGzqjGsEfqpEez0PBHTh92cz5Kuk+fRdHEloCQP
dd9J4z1wXPhszIawjqadm2hRhPZBGzWeBwF7OWDvBgqspreKc94UkhhO+pumgp0R
2M0cr4DYQjV4I5YYB1qAmRbyi4AIG+o+unWRKo6A1mpli5H0vGWRKgp+laGDDYM6
ngiDMqhTaNMq7EArKA/kEywBb5yz4g7RnUsfz3SKOzHgkG0CgDLJkKq8tD82aYVg
FoHj/iRkWgbVHAiDMGbzXsfFNAFitf6IQtqaC6nGotA8IbbFwA0rkYqFP8Vme2n5
XV4TqaSdGccL7gv1U0ycnfIHW/5Qtk5OEuDkSZR9ObdbjQ8Wu6oYnfvtG+Zzqz6o
Z2N4QHc2gk925lJQhBDxPFt4vTIOP6XjwsxgumbnU9+3umIwOOjuqfJG5e+tHKFB
LDIx40m/mHNjAlE3UTgQM+fyeYbT2RICYk2PKfNk42ByvC9dWUYnVWDPKOVQYoW7
TF3zTCZ1pI6ay8SV7qVUdRQqE6HH8SlUnIkDmhghamPOdMm0DWOUEVYRncjUBR3u
NGFa7lcuRxNMzI7L4VnbH553Akd1w1EThDMbpMRHo26jpaL+danbhGVkLrdZIamX
fz6f/1qWvRGCwDfSq2N8afnOCS+PyiGFgVbpV21Z9L/Cp+tHKRvebQQzVOI+ltIe
qNGZIWg7+oJdnFg7bErGhMNutqujZavte61qcOTfk7dsguH4KJhT7hqSyDWxw5bu
4W73qSQAaUaiG8VVtHszJYof8CMKBOC7ypoP8hUDGmW7T2NsYJrFXE1y1DaEp3QP
8oBUnqLZCj+c11kdr3FqAq3PLmaT1Kd8MS4WLlJSrfLi9yeikL/1MpmL4m/jZiz8
9MZmUQk/2ub4AJT5QuHge8I/hLvgkzzp7EpDsn8tflo10LJu90dCDxQ64g2PdWm/
J2aMnSh57DvY0fV4h1El5cyB7PPsRKGTGxmhGDMWhAWtDMcAiX/k5zZ3pHdTt8Ac
/tCOZDPcDlVnL3nIMLDzjOixbg/VdDszwSvRwdCBWgdCjNQeFnr3AXAMtjfFq9Wb
yKkPLWoibIPxbaz9/3kCPu6h784okcaxLCMYpd9sp813UQtM585FuaWOUzB/M/4p
UWlEmkaXioewFgLK+dODKdmCZYX1y8e/7RP2qXXRZwYGPKt3sbJ5y+ZPCYws57Y6
29JRRSBiAIghvcc0/wfTU9NtBfsmSltOOVXoO3+ES/8e8VYaoF7s26AGp+2Zbm2m
w8eouDyFawkEDb9IcWn/YecRInlCngkrq9aSgtgmTJoiey1SOsXPKSIZjOOX5EVp
qs3n3D9g4FSZnvlYMo00upSdLYYlXN1Y++UeZTcRXCLCdYg4Sl+Jj1rQGE6HQT2o
70QSjn2jXPxG8Db6LOiPR3GRfRKXp7Je+tlWgk4UmzhpPPKaZ04ZfGcJtBXkh/sV
30St57ZvD8HDpd6Bk0TqrfN/2zV7d2bUKiAtIH2rCi04wK5FxgdlewsGBIid5Ym/
depT6PfialwhzVszKMGrqUBySHzWD1Qxg4fmottdHlb7+WyTKRAzlihFmUQMKney
raNSY39DEObi7bVgbWOgXKTbJN7mn06jPd1zCfQOF5B1eyGstSjvGRpI+kZtlzZM
bRHyKTyfkcZRCHG9ERIBk7CFM0gkk+NDbNvn/WoGFq/Vs6Ga8sDFtttpfreJoCDm
Qrkl8cRoNI67TovI03FcO7p+DJU0agxR/CB77wM0ThvWYpDje0Txb2wkpJ84pOTT
GV3nyUQyFZHCWU3hqGB7MDSzz2J/E5g8QV4pQqTfnR825xqf8xkea7GmJcWZ+yGw
ej3SYzi8nV/gvzo8QcrQhg9NlYCsKN0ycdC+Zp/TMurqwqrsoixyXF25E4HP2g0U
fphc/Bu2c3I81GMbhvEXxXnU9BcxRiqUaWkMmsRzuI4ban7Ha58BzmQ86ed7eG+5
EWVunEyfSC3S62WIiYpRnBuofvDQSzgPsgWMyqkKy34snB+HtER2bH4Kc2/d9O30
wNj2Tpr31/NCtvauvrlAOX/MNSkA9rszPZSrrXy8eCEwfRB7DyhJ87zoEFHJ5THR
67ZuIOpk/C3EeOOJ/LvqOBXsoKMAiF/rfuW/opUl+Qb4iWoOOk3aQhJIkOktFwi5
cM4Yejf2q+G+TY99z8Cql+/RYqAthibygmNVfCfbo3El9Vl6/ikjhmwvSeedokAI
IsaG3mdNrOxWxqGGUsgUhF0O5AoMVdblA3N4uqEdrrDYr75QAhI0jO+Jga24GcgE
MlRvvsE1+GJx/zU7SqnhE1CqAvjedsDwzh0mp61ki6mDU4choU21QJnxov/Cd1ar
hLbYXcOeVg0W56NhZtSYyHSBKCTw9Xilf5tNuo6UGho3LiqR3+8LlWN06fewBJsc
5PZWzs48RR4emvo3ClS4wONFoT+M/T/KHjd67qWjhoXXnBJd9hBAta46zVaBnKxB
pOTfzfDAnJRjdlRUP0ZOZC5fY+Zu7yUebzbhUYBrB7NIOTAevO1szdhDHc61eqnP
o4OPPpSxfvlcaNa+zCpVmm9CtfPIG4O5Ak8REFd2k8ADaSvAu57fQrn3ZWs8HcKq
13SaYk2G28i0353/kG9eXa00Ev/cqH/hnVcOT4qgVIPW/HWXT9it90aJZkJ03/fu
Ez+hXtArbKyd/ZXkUSv36rY2oYd4JBql6AzLgyU9ewHH/oASyqV9YLuQx0+Qv6BL
roB/sGYDG5zN5kx6GTjwssVId1FNv6qVwd6iuXKc/SwwXHYOR56n1io8gwXJX4p5
yR3QwhX1s8InvkopXTiwu1UrpygOxO4W4g8IChwyUB2oGosbDmtRIIS/XTtokZjy
XYRet3Rz9tpFY5/MtVd4TQLsIaiABC8AKXkxrDJauNO+JLq3SbEGNZVGlzZ0jhXO
hD+kajdFRnIQbIwAp6aC2sU56OMDA7wCDGhWB5GHXBP2KPknHi3qlxiIo39HdK/R
rSfDFoFjQWebkJHRPXjo8YjBiCpp9G5EFBwulIZpvGK60AWCn7LAjEnArWzcin1o
Oh6wiE0TIuSkhFRyqGjaut7QvntktUbOP45s+reQLUmxMZcED3FK8uFoQSvy+v37
F15lBebUG+D2nSKMPkJyWF+Ssx1KSwrZCLIoAteXCDZBTEB35iz+1L8D/ayz4JA9
/rfBpbmuyVbfY9CDvrKUfv8Qu+4FtEMlaPz9+hq0QSWFp5JfYYrZOOF2D2HNzyAU
fZ8B1qPM+7eAvt5L/EERGkT9isYOmL6gvydrZh0/2O0ByvLVnHmDpZgxYL66VNkQ
54nRIJbQG0ks3sAp+J2O/Jrt7MNKzYyaYxsp7GAMFiec4rF+d+aX+jvBo3pjl1UI
XIlcdKXvNd6Du5iE7d/GJ3kKttQdz24o9FdugflS+102oKSmCIXdSVwKpm2CrdmG
85MN4HattPkA9cCdcsO70kq5oIpl/SnPMWUcMsN28BjpxyBu3ILUv9xiwjRmYfcc
bJTMfEisRQYfeY9gOvH3Bj9JkhPyaNXhjXlZrRISwkwFHJ2ICfurU1X9+Z8o2u6C
77QhNM9sY4iMUNqmWdbgvRj+49Y643wyqbkVJNky3kCEv6SEI9DrXoR3xzIYodhN
576cOgWIQk/jv9zV+sb04cSaoNVfI9P+cQSY0lQgd8WslJgdqF4saLdVxzgY81Zj
KVvRaXr6ix4Xxg7XsomYCJcvpxBnj3Ho33HQexTk85RQwgjZ/0xfOR6DnmeRdymN
JhaRB2dy3na23adgmppagIychNktrhhIyCcXu7aT3IX32l62MYj6wjahFtGCKX4+
wmRMVwjSFKei2C/spLMV1P2fZNeLKwdDLqU74ixQYFgcxe/aprppxQQqC1RJceYm
NyKSWdVchUtPAdcS/TrXmi609oo8VcQKAtD01sgyvzQkpcuYL2jAvs2ZDu7C3PQC
izIR85Fj5hyh3BGLxnJP9iFy3aRLfB9VYsNdDdXXLh9UNJH1pYoDI43NNuEVgR7s
gU+TmDNyoaF8SnrogkvqL6Bn4yYHLCXRV/Fo5UNcMOgauOjqRDDdOCJqBBlaZpKN
+iMnY+YlME+/BBFfrT5p5Q2HyV+JqUmHu3faMIpJkeKMiKTsI3Z5tua0MR5rsNA2
cxbDUCnx1BU1596pO1/W1omlFAt1FHq63l4C0xq4RYlU5uGWX7AtN6kxXCE1O7n2
tzp760mKXN1hLnXIaTzKHwkT2oS3XoIWzIOBQuNz7/cEk4qM2ioApOUJgVq8ZF2A
qu+UtNqUaDmJMGU4zLvI9wy3oMuM4c5I2VWVgadHaN4mC8GUhhDV1JPB16LY17MP
2aYOhP5Tq/7Q3U797Ss6p9Q8TxPP903cBLY94+WMwu486ty/q36bEhRMykQsmFfR
R30U71ljbB2lXs5dRnuFHxfupNYF/8c5J3gkT9Ta0e33VEho6sIz4h8beP/FgG9C
XbTvJFfk22aVZ01owBZujpZlGsi+M2eUAqMc3fwqnTB5ZLYO3zDe+ON8+X2wzZmf
M2clCoW+pSYWtKJhebWzfPH3nuGE1uTci6ObQGEbK/W9I6vtzUZKOH2Rb9wUYlbO
DCrdf83baJBeAIgEMbnxaXw5vJs/OHXlfEv2Uw+nhgPSzQsfw1HSMr+w5Kss+PAM
CPtLx/GU7j6dBZ3jI/l6fdt5OyVOlH5Rk6sZyn25gbp9rhCgmHp06gU5eiJZsaFq
sIbdZEJLae9Gl3i0Um8MbM5kY26djmjKpyHBBV9ZcW5S/nMbsZqsANp193eesDZ8
LN++EuOi0mQYd3P3omgTfnzRw6O5+UvvLr9giqDMRPpCXkgqFLZp57l9tFeZ35k9
NCvArx2w/h/JAO01eScLLN314Pa1I9NChUqs3qGA/nzVe2tEnm9fK3s1V2ROFxwe
5wnjP5XSWt/TIcoYuN65Or75RfpvTdsHDchjMhQDG5SpUAk6cdrvjl3R4fbadg3l
LTDMnBmRljQwo8Nn96Q/ptAmsew7P+2aZdVbOCB7xx6F1m4nUlDwXMNBjHx/hxU+
SALxjAWvRjMXf3qhJ0Vo9hkEaCqZ4/F8p5TwiqziteiuMxmVGiRf4yUtE1K21eu3
gVIN+1Pd8kM+sbVmQ8qVyKioFbkUT93EMD+mbE5qMlY64v87We/+kEGuGmlWlZdG
MAyo5lURe800vzT1tsr3tr0u8HntH/HUP7pQE/vi4jO2opKq2a1K1l6e6+VQsTji
ZGdCp8Y74QtmkJwbrH9BgUBxH7YZKsFZZOP2OFFi23DVprHeHXmijpSUXwLTyvJh
sfKqXawvgoUK1dFX/2TKW2il0NUQvNSID9FjNzgfqT5GrJv4HLijCk0GPDURqtrQ
greotlwSwQugIgg3ei1SOzHrRSww8T5v1L7cUSrXKnABCktQdl4AsH/4tEMCcmyr
VUf4rrVG+RML0B45Jll4vzSl/XIVtvc6n3LYD3q5amSFSscjONLHSFZ8tSOI8X7x
mQDm5SGVSRySIxjAcBAEcswkUc/O803p8tUox2Gxzla+zCIYOJ94TyldqE9oslHS
JYaq3HidllnA1p9TXoKaKdSEB96Xs2+VU+yHMkWeSA3JE0SPr2c3npJOKhkg3GKO
govMvWXUAs5vKK8xzYF6WZmFXy10yi7L/OwRyfFpY8XP3LipkB5/M8h+TU5JrjrS
3Dym4Ed3EQsXH+bmwZ2NdwueQUx3O8lSygHgBdiAw3Sgy04T+bJ9PzCGkk7AyZb2
12wASul7+nLcjrRDUlZ8ZBSu7miBwscnZtaQcspwAG8zsgE/up2LsS9E3XS3BlMb
YMy6jKntf/VodkoiCV8w4fa2iNrTZijpIkpf5D7uvq2xbXrkjk2ZppfEwp27j1RL
p9uaOpbtrRpFiz0snkKTqSNWj8W4KYCxmRV3fiCGyW6qmAp5HaCR7dJMkAEjzMpp
CaNcm08ndha6tCo3zx9Honsja/SakPhpSvqn/zd6pQo9BGjpDdr3uGF7F3v18gTN
t8DPHmZFyBF3/Ubph3veAH7jMUCp3LydRN6kaf7OccPdwY54/GqGSV6QJa+wBT2B
TufbqFhqr6w/rHmW7JxR8rNDYmA7f9IVCuY9yJaIR67wGT8fFGJMLs9hMJHIWDJz
vJtY8I6096lBpwO1OIsDBNIILKWnpSg0anFjkxf4CecgbUNBfxmiphd3N2QbWrOD
9071m5tSE5g8fvFAUVhTTE/PCfMEWT1wpZh6MOBXLNMNLXmkIsbO94Z0pQYgMdA+
eeKbN1RO5n7y64dVr+RHPEC/toWsnzZb6POUAaRVcKSg0hKbxGYycksEhBfiEBt9
f4EdI1IyyQeyj7fHMxKX2sZk92kKwLE3VYybMZVXbTJBbT2LeWquerX4LdHrqf4I
lVaJRMY1cQ2E3A9cuRh8S9mu2PHK1MDJ+i9Yl82joiyDsc6c/1YXFX6ljNCtOJh7
PzPhrejaa4jhfYUq0bn6T6IDP3L0tyS0LRY1ql0k+t1YCjJFeuoyxbroXpf4bE2v
6nZAPqGzpIMmzv6kA6D2oS5ZKcAS2GmRKYb4sWavG2WjGkaamZ9n4zhbRdt63meq
YGSwdyxggdwhegWXvz111LMMCRcPB1KbXcY0IFVRW4HGa1wB0pMyWA4BU2U1azRj
bvh8xY/V8wK3WZzsc0ncFvA//3SoGCr2IU1tLlxq/+xOY2pYTpU6NMZL+eJIkj7S
fB1EYfghrAhIK/JvVcf5nxF5mjO6PVNlB6UjC4JAVA3iIJuEI+HUp1NRlx3i+cLz
AtBWdvouwZb3wOJgsjmrPGV7Yx077UuWujm/ayQcJgqWLhhEBYtloRzlpoxc5FM9
/ybZItyqSMDc1hEatBRceCvf+e3fNpvVoWFmaLSUAIm2Ebb/Pr3LH5dEykaEmRA2
tWUzYJpq7QgmOMZXyF50/xdNTQPlXgJFGbBnYz4ADZXo8XHfiWGHBHmHmIB9FU6O
ZpVuj8xhQsDLdUPOB6xUynAsSA03cYooee3Ca4D1cKHM18xirW+pw+7WjA3zGsS5
/MVri5eSTE3rGzdJI+RUKnh2NZ9ga3eALAzzBmj4tQQogVCIyT9RMZReC9kvcOy9
mwM8NkoGKUfID4XOJrdRhVwGgjP0VtkE8DJZp9AUoHI97lFj0iRU8cKlcldxB2bB
kXxDjGEn8JuUGmIbUDJmLD2peEJVVW7yAP89hzPlybrztZ8xzcKW9QZFzmXylG7e
gtjtLUb/157Hb65gebP7wo207VqtrOqyQ3Y6MZbftjOEX17iloKHGAyuKjsefJfx
UXGfoNkNEtEXFL+il0zNKeiWSzLA1NGVzwzRz5TOX5sAlsGGfhiEgCv9e2muW69N
6Sveq8Vk0mvCZi+D73tygm9svzWsNBIzsYpii9tMVgxEiAfVKxmtiDBr85SyvtOr
2vvs3ubAxXYQI9TFnCKmZ1wlMx1cjcnEDQnDtSh2h9rb45eWu8pUSquZyZhLV92x
TiLZArOIb1q5ibx4OuLZUZK17rDhmjvlpoZFAtZXm5cI/HL2y3p9fgiqAu6IAVSt
q2FB7iAjWbns76cwLQnbJBBQnQ/r4kF4touZ5wzdwSkLlfi5haSZ4z8xYmTpCRpu
BhjFKecKlCz8tacEGdlY9a9qsyNyT2wfJGb2YhX6j39DmyxI76xbHIBIqPQfQXDa
oM845UupQXQR2siNMAlWCb+JaWQBI5dHBWYrJkaXCYUDLKSFTMX1ItvoEM2ZkiNw
58mH1EKoQh7U6JBiIisXEKnlJnsFh+bIexVkr+zjBoJEJrwtNAefXyWBNRXVg0tn
TbTFvZTurLDb/JmMjidmEt17Tz4HS20Jn1AIVgqQaLygmey0PGH8QQ2w0D++GjN0
wbhkFrucLRgp+tT+QvoQE/Jbn7cRHmn3JMXRESyP/bhLuB2PJsxhWpN76hBHmV+4
26YpIlx1M5zeGVfXvoZK208gqi5KAs0zDk6qrIV3vpLUNUfAfI+XIxJtG2XCOeZ6
3f549XVyNxAx676Fjz+6NXoaACTU1kqGkYicy8qShrwM78m6iRueQn1QNwh2SfRk
N6TXSoHoDSUeVk73//Lk9lHj9PYpAa3Z2ISEySMCezUERp7tyeAMoj0NizwY/xKI
y6BYDv8XNtPgviIL5CGx+VMJ0offMiZIwM+u6tTaLroGzbwIahS11v8z3VVEntqo
vZJKb3FUcSnRCK8Y6IPqdY7zgnxpZZvtYcLn3qB3GllJDCvIUrTn8F1rE7muQ73Y
bIfyg6tQGw2BxH7bafYwAgQZo/5Yrg/E1OCD1AdI2wqIjfw9h47/D2NRNUpJZTa+
QSg3ykg9B3aNZVdpr8A/NuAjTuuf18T4uUNLsfZpG06BUiC2eV2WNXKZMrM0oiAw
jIXgW+fLNwW1tY5xJa9sAGV95u4M5C4pNj0zV3nZ3GJO+yVoRqDTdgHCrYdzb3LS
1Lo9EJeixqMUvIUd8x3M6nUPAFt7kuwBkFr60ib29hzrdLlX27cOJTQQS8j/rjPj
WK2LPRzU25ZFpHnJqSUPszz4bnYk+htZt6MbS1IjXmdOG4/sf68Wi1dN9qf2GsdZ
wI5aboAuddjDBYo4/Fck6nBeIU52K2NHv7pLHaUXc3Wnaz7FuzRQyiH9NOAB31HM
vWC5OBouvmeC2xBEqaJxacjyxoMJoolskidUu7UJyxSEB/RH4QTlzQSxtc/PkEDt
yYwbfA3IoHiMxOYiILFTFydacd++DIfDvq7zt7sahy8U8nql4yaAOVuuZWZ/bU1T
b840GP1KKLoJKP8ofPrMB15wx+lTzs18VXBaLTbPh7h0i89Y28qA1fbdZCfIIQMY
qC4QedFDUYElaaaEy3dRuZtSWeRCEyz+PbkPiOhngGykT0MLkYgGq1lY0w+VwTiT
eVoSKttumdiLiq3/4qk9uM1vWrwwkMVi54T+JiOt8iloOEDQ/hWumexdcuHAB4z6
z3ma0z0ju9X23lADHtE8a0Rm3fkUKFkOz192qUWQChJJBYmOkk94e5RNH/8W2mgs
WfXBeMPj9B2AM4lDnqbmjWCHmc3tJoxnMcc84Q+03/37WQp3d3nDDBJKHmzwdGPT
16o9zVUX3U2qwsSOY13IkfkX8tM6Wfa1HVpqaEvEI1SJJ44/5fM/47QFNYc+FKFZ
XnEqlTwZkdn1tnXiQv3BXSe2eop4X9FpDVX1tR+ZvHX8UMQHNYX1Vd1GM7d0uCgZ
T2Urk7eP0Otx4uTX7I/Ardje7u/OGZyxjLZWs5ScT8fFpyIW7kSpB8WBS6wiOpyA
jLCCR/KzFr6J0A2qC8GoSOgyWCQzC747ldfb1VmIyohgJbSCoP7Mvfa2P5a6e/xk
THgQJoGRr9oPkrpF0eXOpl8Z/fLfMYssF5Vjpk61lLmLsQ+eUzCJfT9sgMU22ivH
Z7gv3uMP6EUWduv8RSSQFJVpvpXaftQAosjiojRwEilDYiS2CbwskugEFkXJByLR
VHx3NMGCChUmZzffzo3XUJqNBAX3LkTR8fL7bfc92ua8yLD2xYzyBthKcLPUwAUt
NTIrUxacgafKD5GVH4YnZMtqY/EoxIed27xkG76E5m8nutKIzfPczN9tz3T6R7s2
IAreEVI2AS67h1jQ2TlmIngsmRxotnIHldsU8jyCqQ7v3AQfDCSKRiXM402Ji9LD
QEc02/SnhQDX8lK82lL/j4iYazR5BPo7g8clFNSfZhGSObQqZBYHJH4d00b3Jjw2
NhbORTHmvEXolgpzo4lzJN38vvxwyjwxRwh/RzTF5Vw6hCO8II11MbY7uI9K5Z8r
EomckclXu6vCfQZR/m+HAcRQhrVEbb0wX+dE31p+nbT7ZVmCve2zwCULy6ahTDpc
wb7AMvrIvSb6QR/Ov+7zOImjReiv0Rc3UtKr4yz9RGKqeqOKx+NA2hGv5mXIs0ep
ynB8tffF0/d7SMqgI8MKirb26FuuEgHZxECD8fNiaywVUriZ2K9PNGQu1jzNAVjE
bASenakB6p9ctn1U2TI12ki4V+zm9o9n3fdfzxHOi5NnsOnV04ux8EHgRP4Qd/Gk
2e4t8eTA9YfJ1VEnk1OqKHno+5BsoL+dU6isQ4D/Fa1RDCyRHur4c6tBFA3l3YUc
V97pEo96JjufMwVtwsn8RlVLRqKHNgdt6Bk7UjrGDQEytrxEA+E0DFzJcqt+qY7Y
3X89BK5Bgqh5ZbUl3nh2usTEm5MoI6e4Rh6wO6lNBmwzVtR2JZ5tSwA6tODm8usJ
FsDihvBkrGz2T9HC7kguh7wrV/l3eV5kz+JIwijkWl9dtlRo0kODCXxG+H2FAiTI
wCW6MHaWC7Ndi4lt7UKclsEjMNgk4FJB6XxvXjgvONvG68Qi6qo8MGjtKOq7nSH4
Kb6TA8cVRLamyZ4xaHDXCWDMDURthdjhc4P8rbLL8rgsGn1/gmbLPV6APJAsL2HM
WsKoTTj0zchQGxYZMSkR7j/BEdPXA1o1RGgCmhIAYKUNvIghGvXKnhxAtEze2k+t
NO1Wgizbytq/deVsWvT8nkrk5bGVgpEwXOyWCXQtpZMNGaKw7ByBhlqBI0Fqd9nF
pofW4UbGd9OEXx58rGgTT8bjzOB+I4T4K3zI3MAZvVc9zroMIOXNMDgwdo/21gWV
GpCvXvvEKiaVVodpgJom+A/WB+lCjA+3nNRUujuwgTVCR0R/peIa94jqfImtMShg
NhvyynfrVAvfq6jU6R8whZeeasbQn1XfPon1Ss4c0DJ94K4fWhD2KnxhvYTePrft
KO+N0EqgW9TpnNjgJdiffEFZKIyj3FaVBGLY+hj7aEnspYAZEDnV28I2i3zKcEoa
1a23+P2EvkGrCZRVkT8QQRhfA97G1ue/gZWYeBCbnbu6Dk5UmYwvhnvhgxMM9fyw
cMliqOl9XGARZdycQkmhIKfYDcg5swUFJ5TsAjRJzy+gGDwsxvUBXH3aDU2GDES6
YzoKlcKLKcmE3E0Fxb9RNn2hGAfg/FHrVMtoaSTF1FT7znrRRX28vwS0nEyjfFNy
AeN54X9KoWRSiQPj29obTZE+Womzvpat/VuTN75xmqAXjck2AZb6vl23wvq1FGhQ
WxsmRGwKj/29j0gaW7DUNpNgwR9cvQyRr84/CpfrsYJETTo/bh8eMSbVqppCT25b
QBCEwokgfimW047v3DkQ0pdeqjf3WKrjt3uqvL7tqLMP0sEwknocKLiO/1cU7wU+
Q6bopR8ucXMAQXlSfSSfk1XC8yMMPW+ebb1gDjC8PBUy0ve5sdsnzj/Mua4grG1u
j/J9zUlLF1PticW2hd48aDQIs+d/Y5gPLSCTKzL5+PulFAhXJeFi+j1AuzgUBEJC
exkpxnZK9u9a0LF20Cw0KSILrZMToJughg1hLRLW1MS+u9n2hQOx8Zrg4FkX7ITW
jm8au5eUjcYWpRNWRX5iuTBHY3b/l/4sNrRwileqJLkqVFuapnj3J82H7Pir0cxo
BWw8e/+m4aLpuqIFH9gycHNPyF2QmYkOnHJuSWhVv690G+AtWBDztT+g6fqoYURC
MWdaue+Fm6L4CQYRQpHLCN7Ax7jpmFUP43+G3gs7//jujojKWu9O1FosUks9ubWD
oWdqVB9InQGresOCVFDTtOrbaDJr3phRbyoiLx1S47dVS+y6RLwdXsK9Xl2NZp5I
H8DQFKD4cHu+KhM1B3uTrIG54GZDf9k7WIZhweuwTUGq9KGmop9HYGEqUYkr1TaF
RjlIhfpqKyyG8HmArrNDEFJ9srzOROGmvIEVX0+5pPwsXSouB1nmNOcl+qGPMamz
qxS+YSnrZqEEyTuRD6Rr+wqNJOZ758NbNK8HZn6uEkwFmsKBIo6A9a9DHY+yf+MZ
y8YXfD/T+FyC2mN9IbnVPHwt87upVTf+RWnWqp3Z373m5bQSXLKVSICkzu9FunvD
SQPNV23qKSVn3Sc4k16/SG6yQ3GvcUpUwXftfT3qOJ8d6Cl/yt05KZJAg6HeoI1M
0vk0YWNNqJuCUHaO9GvwCLL5Xo9S2dHIQPLCFnIT+Q4anJxVVSvQU4+SUXXCjPjj
jx7/4Q3BIJlQ4vsPoZazFyLXKyBNW35N7J291zRjys0ywCYb5nvZSGcRwYPKWZnO
7QGH9/ZdmgnO8nnNT+mW7iLFrngTiW46h6PLHyKZ6CqLDhpwHs/wWtdTjaPUu+Hi
3nvUv6sY0Oc2K52wW/kGab4IyAf0FPyC5zudAn8EvvnLBq3V27fd35khO8n3BhOb
gCkMPTSohsnBA5+8iDbxo/2l+yPBjVPdA7zQ6lqxEVwhvkCu8z+cFCQpa9Wf20Wa
0inCW6CzzqHTEzf79Mt3+CbtxnM+5nMWuLMilZfYA5MInf6fH3s4io8u9nGMbKwY
bsbvFoA4ptTVqfYeafjpHOBR/cD4/Z3sWdhfiphuVPIG9tVB7RnhNpzW/2vKxgKf
VMBSOHnK2ivI6jBcAoMwQlafKKat+/fCXv0zmbjWJ35GQ40f3V3JFxK4FDVFcru/
VTsfHtpjvLBpXGObXn6NEchM1WDCSWCGIanC0xij2nEnzz+hOYVtO4a48M+K21LM
6rwwtLQqH9kftgwmzxUmZFRBix/A5dy0gEjddjxVSdWk1F0nksjpxQP1vf4BHu+9
zxIOipSS5zcfee+7qZSdQ00CjIkdlWM5h27jQW/2tn8kgDPRL33zCIk4Zt7vH9zn
NLATZYWoyFo4SKEmmY4UmoTCRy6PCf3UNt8WHc/kBWd1wC172UrFnS6oF71mXIYr
uQW4o7bEkxIaU2fFkSUzx5Dsohmgx6f5Qy61MytrXXmG9OxHl99aWxZm2de0dZ2h
azmsSKhLej25avWoD97qQeQq/bbT/hfA4LBPTGlZQB08DGCrPy2K3t6eNAnR4aHY
P0lwIDWlKeKNauWYUR4l9MXL79eSDuSy+kLCv3Cp/POQF/cCOJys5PpnZPNCF7WV
Hw7eoVKeefMGjzmoNpH38iC7a5DKi4tRfGhcIe174Gr1dwnohFfMTKdeubGJP42Q
RpOoZ0yzBBBrhqgCsdb3gAixAzhgY7ks6+CwqY2E0KHZqHT0jWFJliqx7oYMgDwY
jS6CnUcTZYngbcX9lfWgcn5DqFbs69A8U6SJZm0lb4KGGLmzWQkqR/lGzdYyQY15
RhfbnrPyRH6gO8tW+tlvMcU41UPUsYAO2t6hmCpdX1Zrq9BI0pCYfo7Qe4ZRLMVb
90RSc48xCf5tuD7twVC91/u+qexjh3lwJAR/0lySEu1QalH03WOiAX7piVDpkfSp
xnzqhgMKKGkQpv9OeU2/zMHx3/ImX3KMNA5nrxjaHjwxIqLdw5lfTmhsGf8cRI/Q
yBna7zeGdgpP5WJJ3NwjL9b0w4+2ROjU5wc41r6VXvzImMhiJNHAzAC1KbHJfATS
MRj1Ci0ecZGW+CWmEwoQve7dWb+pzgyXsmu8JJ4fX7FZE8p46vNGYkVP09+Jjq/8
sQq5GRq7eqN7MuKdt5ScBLh5eqHsBql3Dd0MRoWUkeuDqn6UuivQrAHPpk411bng
QRNbdM6ov37uLYhxPva0fNDUASd6UWLer2ZSq+mJjqYdh0C/JmCy7q5F27M6NK2i
LHNXnMs7v9EPq5yUCVV7ulSQ62JFwZTQt2AH2MK7c1lHVrVrCQLkQUm8eqYTeKvm
1DLDpYhUEeZQBMpHpswoo8PTWgH01kkWuO3XyCbA8oaAJLMfwqcxFJBoxAJ92lvg
+w2XwAgT4+3kytyuyp89go7ZdOglHMuWt1cqHZ9g23cJAwU9qWrwhVvE06Q6DN5O
LsTz6Ol2KRBdYVsDz5k+jRVt3Nv04wrEY+ziZsoeLf6uErl5d+ouIiBfcRJWtqYP
01FQbcAUGSf4FvpCRKDPYIvpOF/YhvGH9Sl4ire+YkMmJ4duaGS5Z7g4O4TTsh3k
a+yhz+vw4Pjq90WXhmJTyctAjgA5y6WychEj0ELdU2gHH+RlqXW1m7pYC2x03epa
Hjpl5KLPmd7hIhq4yYXKNu4DxA399GqhgVorRYNnSgTt3e8EBFKDVtZG1TwxKDxq
mfBiMUxngdjBskGgSFZHG5ICQVTTCp75OspMEyK7a+0baGLWh585kVDimzDBZGzg
C91owRas8Spre0ta7PNs2omi29/OgsHaiv4U4Nefl51PtWMJDUim+/glp7E2I/9t
qsRF0I52Gxrl3rDoIRblsKbMX49xy849yoWxwPXyqJTN2EJkmZYSf1tbEmElSVGB
fGDWfWKj92S4gkwNf15CjW76twGwVvVdLINB6E3ifry5eeRCpVl+kOC4Lmtc4huu
dT0qTLTY+GCeKv4Y7uLefclc2EJbL0x5qD5hHeqH3MhBMWBA8N1AlRjBw+kBQmZU
dIjgrKS/kikTkpEt5O70eKXWQlrUN2sZAlQElmQVuVZX4JGkI7IHpvAeuCy3mo0x
Wffq4kgLG43SlnpSIE0hdbsmoDvnVEhy7kQptV8GkqmhgiDCkxdjOh9/VOwYg9KP
Y+U5macCVc470CcuqUiQKxFbbFoKv/WKs3lBXbB8fei9kwEwa6zBbDm5l0RFSpTq
/iAxd8Qk6yeLbOQVuW/AhwgGIa17GkzadcmOpEGjAiaYWmd5cEFLjmeIZ+4kkksa
RM5vkS8RtJ/9xtX/eVqFTWo8MgvLQzAgSl4IB7JxQq7r2rCNSSbaYJHNKPko0BnI
AvO8YE9MeZw66qUMwMR5Ezlgd9rYzN4UaeTAy4bqvvX/6i99TzUf5wK4zf+i+dbM
z4diC0h7i9K9RtRB/fZfiRnUVYCxjzedAOroaZyATjOvmywJYiiJuDHzsSvP1CA4
iyHeIYvB0vSgxJ744Ef1+94RDkyq40vMFT3k3bCV6xsDxQz9ySkt8FDunTkBjShi
ejRoMfufnDCrSQiI/DUvPSZ8nBMgLAtWSusJOBrwfI23AsSZxQWT/QfW1FIOR8lR
DROU6x351JFqabxEvdMNhKOX7oqh+QPF0YmuvVvePZqxWSR67sEq7QtN8CmVxqvw
fM16hWCtPg3dBvYCo+LSN8V8ZMauXATWloV3GsVU72sFq7FWJ9qg4b5wpCtlvnuq
byAg0zTX/6VRWRifZlKAZebm3vQqREgcUz1FwmhFvBuENnrCFJb/I6IuihIzbH43
4rMDL9rObU56uI/XTrBxKg0JLlT4LuZD2G2O7Ju/HWKPTXwCEVAiXF+ZF1kjaoZ0
kM5LbLhrn922M1fgrZDfKmE3y3QWfTlXkEATCZWOZb2rxy0XBZ71uvri0HaNra1d
fAcFl4nPo6y1LXWYbJ9EzbBNgbbsYCnKnrYsNQ+RTcnL2laWP7IM3DXFyDpLGF1x
pSs0Po+twtroExZMpy3YfKIpmtaulSjUG58bQMXM8tMq2Hfd4a9Cod9zq48AKH7X
xK0OeCADVFumK5coWe6YHDZ18wuCfiWkW8jKKyxysSIz78cCWZAxk5/oCQBcBET2
fdPafQuKjUNh00wllBS1EGIIeEe6kiNYcov4kry9A6TgfkJR1qWU1l19QFtZLUSk
ox1h0L4DbdtrnIdVKDdOLzJbXSAH1KAx0Xkj285KnJc9V3/V9K5NkHI77TWKVg7j
c620Ns3+9azlAKbCj4DXNYXTUj+/Yw8rL41KE9N1oNz2qXXpi9TbhnTInxPihtrq
ehdjsd1BMFfrMDJhwW49BnbI1SbS//7SF9/yT79KQmulTLf9VDH+KwTA+hCpJS9C
wRURiW2HgAbHxnCYmThYgK4y7RsvfXioWvifayoxzhmhSvn7ONSs9WZ79a5c8Muz
JS/5JGlSUtlvmeAKWlWcmGMXyo1DB2Dwd2/BIjJLaCQpRE8DQKXOy9L+KQ6+DR5B
6ViebBlYsM3OBqtjTNogV7j+ZwIdBWA6Ksb1VmfDT6tvwXyJnRgPWxA0+4nw2q/e
Ysg2gJMzABF7dze2sxLOFD7MmjtnyubIbvTDXPftPIADgaK13QwswSJnwlyfrgNk
GxHjW604RdV2ioHl+hEv3teIJjtL4hRoMFETYYbkTxKNmuvFFYejPgB4Htdojlhl
6WGqSAX8OsR/apDCn7d8Uqm8tfBAWhTVcqf5Nw2s96mhZxDWUHiyLgrasmOhvDad
rWgQYROl49IRM7wJ5bLK3aF6t059KqlaSRuMjG9orhpY0lOgOsaormcITk0a6Zj2
07LqscRGaguGM7YKDxj5jhlsx5twRnzJrOjSlNUnrsJj0ue0ILdR2t495T6PG+Dn
rPXcua9MdxYvl3M632mVQXpJCMmkuQMuile14AZt7PwmLo5sVWnsZInqCBsaF+iQ
tbw9EXdiejajAVxxp6i7MYteIqCYWfuiAPJfQS0EZP6LTRZEmdRfv/MVfDXt6K3y
F0FoiD6/OzGJ55TAACRTVW6QLGsRGLjQZUjThZpuWnpx2YaPUpC9PvDlShqv+VlP
2MiK68udkke0gX+YeQ7XOFTxYFIBACE6f1MZYgPimH7O+tn3R8zUxp3Ea15dODf2
24wB57noziWAkGzx03aPsDAPYkr1FEKsW86Pc4UO876pRMDw0WbOiLqn8gVJU9aE
xl/Hg7Q9EJhkQP3Emsxgt0osSvsQdfL6mjg3EogBwpOPHKGFtXLyI9FA21K05hAy
5wNNE0G8eO/iIkGtON9ZzqLkD9j6p1N4/m4Vgv2cuLVhGfCiDk3i0hd97yRxzGF3
f42Q0EWLxSMPVrF+nNRGqGZ7541mlbyza5uj5EdEbpiM5rqPV4QKVqRbf51ornDi
Dmc6fus6VZFbIm2Us3QeuWMzjpSriuAGZVIr6jsjz6UWuOv15btkL5Hq2lmvyFjz
iszH90uHilPUOgmfV737Ryr2CFQOQwIQ5ypzAtyKjyNQ/E4mZ5LlhE9as0khKWtV
uyJLX0ndGyZA05j+5j+Dixq3DANtm5hh3EvaBokWAMEfZnaEKE1lu2zCmUv3PDWu
m34FXqIUCA1WYuuoE0+QaqCgO4RoLDGZggiuldm45xgBVPOyoc+VPMUNuTXtpft0
RR+J3ngbopHz24NRNdb8uxIWCggn8qEZ83bay/LSa38PRu79DJK/rHfrFfe1ghH2
6hprWQRW1uWW1ShrKCNygi3grbS/OysSqO54ypf09o9rZnE1E3KENbyrUImNPTy9
gYWplsHKiGyfxdW9vsND5YtpGb6fvZLtwe6vNLD7wWLeTfzH9O0NA0MwUHpXsKo2
caygSWWca7RIQIIuMq2cXsl0sD9TXEI3JVucz2t2tuhRXIO1G43A5/ZKTAPPDNRA
QQFrxvm+vcMJgZBaWITqMxYZS4acm9i6A5ZFR66HoU0ZzgtnV/OFoC8ediKx11lo
wHg+6diZLoWEKRh6xyCcCnsHDmTSCJYQzA/+eCgxjSA6Ewb8O3OFv497xMzu4zVm
HZUc49U3xgoQhizauetoWMX379q+qIKV6hxKFQfKozoSIT9RvM8rAInZRcy567Ox
2SPtaMK9S6JBQ+rFr2YkD0LVf6e6N9kTRO4dIu8WTUjyWancCJ5IAZsJFafMzreS
DKxlLWufjKxIp4bWzGSfK7zX8ix3BgAdV0OEhyAkAIFKFKI2h+rUqYRZ/EkZ+PGE
vGNplYwhXUlFCmjTLtESZ6dOF1qLxQ3CQpkPW0qBUdMNvRpSkKoTRoNzFqq45kBW
+D+LVL/Q6+OlAGRGL2VI+UyISEKq4AjS7us9/sJmaZZI8ENie1Oer6iBRA9h4JU2
9KfORgwsgsGxlVWWk8AM+opOEkN6lzEsu/Exbq5o4rw4dnGPMZVmiXPGcv3TQQMq
GnBFeZvaZMjytOskUvRsAcwcHvqmXNGz7UQaZg+KE/b+NaNkQdL6ohpbcWHh6ePS
UMIuqF0QNBeQjiGOlS+aAgHfKdOE0aBeC989G6npGOtyapxl/isE7Aq5GL5l7Ln6
XWbHewWi804e7oj+wcBbwgm9o48zAIr09MZf6apBIv7GGJ1DYNafOXktlA2BLLYu
InP5/Tlh4isy9DNqYm7KxW0uSDsW/FzSAtnE8F1WCE5mZvGqnXEuuCk97hTz2yRL
5md6s7WpGx3wcwXzJBWOqJRNdkJRNcyUE0zbvdfiAIfC/s2oY/SsRvAhZlunUs7h
XxbRNDBOQtWqR83UdBhAo1Kcn1wpw8LN3a/TMEzXzFg/nP2uN3tW72ubjeBPi7PD
dCSsKn3x5Eb/ZFpeGU5Reea+1oyWR73KWWKDUL+SV9r01UN8xQDKethy98cTczF0
IK6sTQf7SdjAjilHm/sBTbDTaHK8GmxvqwNLz8TMqMKp5Y3hPWk3pzyqACdicYwW
Jo7ThSOi3J7NC4HwsjQCaxzL/0AlwDRMewOxUhJaZCtD8odaQ75xKJZcQYF5kb+s
Xi9GbPynmTE+BJMwIXJSKtCixSTzJrW4nA536EBZ8q40M/ufOEPiA6qwdpF3WAL4
q1IVzGMQD9w8qJzMO94ZC37vJ+1LbtjBeDoDNmKSlDofrepRl7NjbcnHlvQK3kkV
TpN2+Ds4V0tsyIzJoXpZMSCC/lEkRDksUARs6VSZvYCVxrXcT0JJBPwfsFZOroTL
mvgEB4fLIO14epnolJREclZ5BE8cvLN1H1rJR0xZJLW0BCgsMHQ6auKdJLY4dQdf
AGujZu4ME37Nk10SvA3gp6QwC+vfHHKeb0RQZScAuh/CmlhksgYo2wvK63nK5kmO
hcbKICuuHt6SobYH1bz27A7nqPgcLnIuRTEXi8/SXD/5x4B5X1V1FX5fvVFw5byF
JWV7SHZVpnUYxownKH9sXQ59+rhOEN3GpI5ofHlBhbggohDn3+MHa7cWTyp2BLen
sCuWcorrESl03fNMLlZyHINrZM4X6cfLOmPuD8JQX9DHqLHVdQG570hhjT+iYCka
DLEq5ETGv6eKmSW30gRCTr/Iomt+2BttQ/ZcMnkhvfcL3cCQQDjimSuoGG7fGP2c
wKbKvc0ZqdDzrcTvf8DbKWx93KcIPN9uwIZd+a3u11lxgLF0YQqhGMDCEpgAMfNF
RmqJxxcdWkPsubEQiJ195LFBsnaAqsW8GhXWBF+SXjJMVjL+dOBwN+1+YC7MGUg2
ctYtXoSv92ZjgLHwXWmfGVnXlj7O0aDtVaqteRK9Xoc+qxKzEutW0MLwVQQ/bdRp
eaZJ1Lp4rwsW8LPUCMgrRX2zTeIPRGDnMBdRGTdKJ5Js1DaskhLn929s8xiyFO/u
rCN5cKBdJQjXBKhUGd47zqdIMXMT3JnWQOZyKgagZkKXBE88cuVe/E0/aLL9AQ2H
UDOv31Lq3gw2i2mqJstTs+WjxocWm0rW86AdZJYFdohdq3rQr4t635DyaVujsVyy
fQYE9Far4WtWzyeBFjQttuIT2sxSiIC879bPZ49FHykEe86FZkpVRgJsDdLFsChp
LucTPZq63LpH4nU8RtLNyX5XnsJc1YhMbrf6VKZcIHXyLG9FODQiAUz1niuESHPu
ytt6nMY8UQyzcDUdjFEydwWL3CMbvCBopI6blmRlAGiXLAYG4VKumqwD+GDq2kJj
P3r3c1sKq2/vSyL8BYfrreVj5drbcMmXl6F0Oojr2BzcGjUF4eqBKpZ+1s6B6LIi
gRm5fh2ayroVl0WG6D9GXydfeY2a+OyEltE4IDTs21os2bpk5fG1z2IGgAErhazl
HZtUEvEy98IyAMzhrV+lAwW8EreyEZUoNwnGfPE0n7Be8XDARMXeEYnhJrWz14LM
QZwtaI8etW1uRBAW/FnGApYQaNffGS//2CFhKaFKsTt77bn3Ops6DoVTYvb4Q2kz
PYKc3RdYc8nzIMyk5U/5bhMUeolCS0W0IQCaRUH3VRXAinaUi+JN5jRSrkny2cEz
0UUf6JtfsbX257JLyp/8z9tWZofEX6YsvN7zG4DQbqngsazulJkFlwIX+9TByA1f
h3DlFVz1R1cfxa2TYFaYIwJPsDG4eTEoQ5pSU9u2amZNB8tkuNelKeYJAVP0J6E7
w/5k6zBPkNW+nV8gor30JzMW2YsuHANeSUhPLVmlpshWN3neHEYbfztkQNFWTELr
hTGAC9OK6K5YLCt8c9Bi5gp9Zqg7miF+qWY2bDXRBHAmMCyzHyx2aPzDV005McWM
8uIplWpsiM0GMyiYas75Z+KpIW8wgHY5x/OB1jnUgC0td81pPTfCnrnJHyKS0DtE
QsInTOrFmrixcvSwREPokegHOrB+ohJMefkZokrCadUb/9V+xeweZ/6swqz/+DV0
eUPnkLoMPWW+aacg/3/SuklXJ4iVtq43TH41Hqtji76ucl3SFzUGXZYw2Ln9adFA
8sBVyYjRjX+Mgv3yjLQIErUW9HHMCUmpiWHo5Ze6qPXKSlKKFL/h322AQp/gaHyX
zuLSmMWKJZc5yzmZPadTfpZZEqNJQtXDEYlakKjRZTFB29xtuJ889j6wd4rZsRem
FCFx7Jp2lvXaU4FNo2A3NGW7qRnYnefmOtYRMAtu8+tL6R+eSuauxpMHRwlT/A8z
MpgVtvgQ1nKMkOi6YkWrMRT3B89lXBHjLHNKSqsHRJJrpL0/xAlpasCtr4EfKn7s
Hr6LQqMaqs9YF4sVx6kRbQBNQF8mvUHZG/xuO6y0fnRWk+ytBpIO2kTnvJM10bZB
BF2G8aYjmpcLqsVSM3T7rpfUq95McRDp3TM52HflDrlmuH8E+ZbOkboP6HfSm7qu
z0NqEJLSPX3X6dk3rZCfdEVidovM4G//CjTVmKb7UiCnk/HnQSP7/1DvJGtkNMP1
j00fbX7HRoKWvK3dtV1q/pHUCELeihqFe8BjBQH3nnR0i4kUqvsm617ewLF+jK4D
0t9QGDWc4R1jZg5GtdsLUfbnROeAFraA04pnVw0U+MyVyqti8Nrv9zjYyjr8XjVI
AMEmugiHs0/OPLcTcG7OdkgdPYF7phAw/SibcZ6wtnR4nnjaOR/+zC909DwCaYRE
26Qa4zZ6p0pQknwvObv1LODlkaAOsiKWCwwBUUvKGgYYDPaXD3Ry97Q8DrivV8Jn
EjcnLfP6/qkSknPSip2XV/2tgIH8kbQKH+Ot7NOf+2vRFKhBx6ZyRZVyVnaF1D2D
mHohNQEZarVP9qDED1Zi8F6zyHxaXtPJtfF1r+pSf1I+xmTZzQ51d+XNDTQ5ef2R
mjUM7ua/DQIFSct9wfmKEsDCTYOyHlphPMZuLhZxZLGqFscOLD3hsDUtBdCuWMrM
eBMcfM05DPL5Ptcq+3ifZo5OGGVsfKayTwbJpN4zYFuouHY+CAa6MCvhMCb+MkFg
kN3AU4tdCQ+Y9sFKKCMs7YNtSCnxVE/GVgStDUTMubAVrXQvckBLhknyF1RCBvLB
tV3OdAut0MEhzjdGgfV9iDfGIHwAb2HyJqcb1CBdLgduIv787DKAmS/bwB7Tt6/7
UrfGH4zTRiWFGj5AFpYVojvh+5/svgHOKrS0Q7yoWaQSs6ugSLSw9Wn610w8E9Vl
OfmIzihQbezYWmaf/PBVkV5jzt0dpaSJYKXw1O+GlzdRRvnEmqFoOqNbb2wAzNQx
4QBguT81vkBvbwR5C8zDsg8bOewLyRZXg8BkkXsCodPP0xrbF53HRefpfsl2NAK1
sB9JWGFLxGziV2FbvRy9O67tTm1GmToYKhnWY83fSinzYRammqp/IAgYpryeZ+/X
77NCuCdFUOEQHGpWgLQhfiCUU2qkZfS2LaZXznC0NB+3fE0GJRiAAwPtxilAvL//
LWcEwSyl0A4ScXoBCdXl6ddNmXt1oI1XsHv53+vo2Jt/x8KExfILJuUyl8Bdba2u
Wj7jq0wrDVNymWutXwS74CgUlljUZn1QFA2aObcXMIoqdzmqdYx76pMXfmA6ZVlo
8m2lKiGPYgnWLZ7PEOiSNagNs1CBqhmlTovnDBbrulQe80rkgAWWFj3EmxifIyu1
hdYih60rDTdc1wOnJyQXJOq+t5NEau/kp6I/PyD35KRYjU888kblqpzNx2/cHqz1
64HWXIu7kwscBkg0IRaLZ2eXx7ALKtPTY9jMOdGMyqE4uqCEd0bDuRQ+fD+z7ys3
eJ0lObVWJS8EIxjie1Z2+r+jDDug5DuzO1TEFS2KndOvIg5rujS/JNuwWGmnGS7K
N0JdLwcpH7EDKoh/nuulBfCaJSX+xdEWnKT2pz4463uSkbGpDewWiEwpKy5mI1CO
q+hfoPmYg/23GV2bZYiW9bcvDsIcSlzQzF2INT/sRd7Ly+EP9+aMN/hH+blE8v/5
iZXAASrgJ6TQ+MK4FC+H8x3bWLX6h7/UrDkwclaNlSv+aa078Mb/Z6C1Ir3tslWm
vMu7qxwID8uJPAbT1LjWERGomhlWksNtFIMCf6/wRaCvA7wq/hL7IpEpSEmjTOOL
Wd6YhEZvVrzrCgEEQQ5YweYY9Pz/9PUx6KdPi7l91ASDyV1rfONN8Ftt0y+TvWaU
r9tqwu4ZnI8qBdXcXtXxQgKjme1QeMwfsTWdVsyB6RJl7k6UgUcLD3bWlZvHf2rf
m/dTRJJK2y4YG+uVDxvlb73WvOs/oYOnIgyvrbZDze7db9NVjCGqtwPRduPLxrMW
M5ttsLRXJW+LsAmg5ewdVktSEO3t5QiNoumRwjkfIgbnGHgcfBXCWR7XoBgU4gXq
se1Th3eU7X3AOcoJ77dI0fKMspg2Sn6duKODc5+BusZwZEYE2V9F6VNW5qn1T1aa
fJ+JOdy1gCmqs3delbyeouINy0oK/gmdX8wKOhuzlHGTPPsVl0GxwZOkSxpDihXR
0PeuCo0agQFmVGaDtxTh/2P1GAF4iwTIPmRE6C7/6FQ5+519N3sByyQc+rOEkoJU
uoFqVa4WFY8TcDiG/AlZpqQjsieTfr0QejCfT0CtdU9mMy3a7E3SW/erj7uzYlqt
Ff1sP82TTYqzznBBeQI+wPSrBL10TqiSJtHfLoQJcpLPWkuLyeMGGwVkoMADU1wb
++uXRIOEWYMwNh8kUfFmH9yZM+poruyjfWfK6PyMoDE7IuMXRnGXPHjAvWtqyx1L
KAzFB5mw2SOm5EqNhEHfmrjYm2P++9vRVleSIbwWsB4guj/fr0A9pnIFGUmGzof3
IbTDEq0h5/ms0YWOSXhtniuR9hWuGnpIuSnCk1XmMOSxGewDo6JdXYF/kLCmdpXd
R/1KEXgj5TFsS/u0fsS32QP8vu7/6iG2MgiN/pP5sFvXrM/dOIOreTaCeHHTWKin
K07YKPXuT4ahbdraaT3IHroihRD3K4FyThyUKCqfcf68otr0MkWSKVdty+4Gf4im
noN9a4mnndIN+gtGWHIVrpkfcOc1MNWVPke39XldrxN8lqEhoA7XQrSrM/vi/8b4
dNLL/FE7jQrybK2ux52S9cUWisuxG+DIgqdIfBXDsJ30HDJkJS3Gpcsjo0VhxUdt
kbRtX0YgEevrfEXfJh7Taih3jec1TS0LkkbSNPTMwgEAbwtq7FU5yDxrGdYEjB3B
qXSUajJqeaFMFE8hXzq7WF8YPBm0jzl6y2HsSvVjfVCOYUn62E8eQJEMKBFpvCWW
6pLke4kAm0ZiDxN16W+OA78nIcy6+2vkvaE8scnBSZReH9jdCTJANa+61VyKM0mo
TEyl9bsqAuXsRD1f2bLRJ8aUS4BtNTr4oijIkIm4mqDZFW5YwHUL5CEsLft5i9C8
ZTzNlC6JqQQCIe9AlkA3wVE0ZEACkNE7yfUZgtLzR12fKR8jsxsk2zth/j4w0RPz
SknP5Pu9aivWtMVwr79xGjqfTHUoLcOH2ag2tZOKWIzNiSSk9ntoOpwHyXEc6nva
TDrBF565VRwoVsKbKPFK4foB7g0sJEKLQkzAcrlU9r1ciEZeQvjxUvXvXLNAYC4u
EdzrhF9B24HK+vMov39kYtriAns4JGE916TzazM5KFJFSjR4GrrYdCT22+o/SIZ3
Rg1j38967ixZUIAfcxx4veAe1rZr85FsKesi5DAcDEnirDdULfj6rClpNOGK1KEf
qtJpayhnRfw1k1S5j3Bog+MjcDKkYyNG7Uw865CDYVEolk+H6sytWIXs6fwojDWN
NqJzpgBQgekrehBwHygTsMDYv82U0WButVKEV1LH5ZIuGU00/VboU3954nSieT+a
39dIOyE3R6S0xOoWgE2fikP7tg7zyq9CPqHEVXwwWxMRFIfcMdr/5NsakNzXdDeQ
+IcQadhdFDHmS6S2dgVjAYlWeIREWhowBX3W+or3P5pK3tK61j/j6q1T5IVMcR9U
ahTmbh+i7hzSQOUwv3rLxaPWC/BDXySJQC85VbvUf/Srdqwd2HtSmhg790/Oz+kd
J5HR0rjzWS22qCNAf7Q3SbVDu820eBNOMb9h2G7p5RPUn+JVUQEdszazHb8pwyU1
KzhLvw0oJVku0hpVyk5xKV1vA/Ef1p/Ehbl3M3Mk0H0pa+GJl7rth/AeapEWASYa
AfuONt6BydtuPOw2kBCqstcyiPpuKmdfn3rwrqftHbEyToWGGAaE5FWUuYbHwV/f
kdr85zCp+hrw1N1jr86A9mIv1fFdEyA1pr21JS7DgoZB1av1NxZoI8hAYNJ+2sEr
7spNubZ0OPjOdMneFDE6ATtnfYV6q9n4DEUe6OG3fnqGOvPh1dXQOiaHUvlnoC1k
4FEhOdpFfHfCBUMwgKH5It4x/6Jcip1Puuuee1pdKP8II92dh2dMOrZgXYoui7og
TPZ6cuS5EWa+y1698CPL0o60Z/5+v45iOgB+XxEU4Tnx8tSslA2aswxpjfadkpyf
Z+2T03K9sYVyB9fyDVjGremRz8XWeTqyBEGDsg1pwqeHKYn64qWsWrsB4J6jo00z
tO21X+dOUB/hEbNztG8XVzyIQDNX+xDEN2tUjidPF7Q8zmqGka9Ubu2yEtvq3N2T
LxtaJsy4ycQjzH2QepTq4F8NTaBqy5dS+Dry37q4gUu1ut1xy9JtKw3MExrj048j
rUkY8yhIHWD3JsOuGz0SGCvhlfVhwbiCkFWVbYFfkS4GExqcjIwELHhDVigBX0hi
iXQRrvW8DHKycMcHWR8X21J3H98Q0GbzCdNVLojO4JVeYDiFVc1v6zLN5Bdf9imj
UVzOUJ551FAtjnedd4AlPPMLnoyn88mTQQM+jOkxhltKoYiw1eYbuFe0LJ+cr7av
DuekKI9MWOmQhoUKshBK120NBnUbZgVBCros2ujz4BjotHaOjzsn9+x0AVdOL0q/
LQxmv9y8YDFAGKxz++DJFuHL0BgCGHtwuKa8NQw6nws+TYy5r7sGYwrqFR3uDj6S
vh0w1XJYgQSlkicPALBouK4iJZGZbGhetDI4ftZBuxd4/7QXnolXd9+ggcFog2IN
Wnw2hMe7EJIZe6Td0rgOBd6ZOuS+qmTNnre0mHu+0U2DJdknYivTdOk2sGhybnx1
X960sPcCHzxRW5X1cEczMX854/uOsI2gljv2UT8xc+Qz23fTu/xLBwVXG6CCaYGC
xugRZX5kQxwPqt5bZz16W2ykFUZNlDcqDcts/u5jnGD2NPQXy6m6Cd3wVkK9Unjr
EQDMymbohoun9gTb/KJ36/AcOfFLQmgjNZpi4LJWafZhal8Qt/kd9dRxOmT3KnI2
QjwZ+N7qKyiSaJYR6o7xsUzbZwzq6gVK4buWsF+q2IjZp2WA9vBJ4HMgDKXcXf8q
nVGDhj35G2XXPnlEWiFHrYHb0upOjoqFtggIKSugYr6Yngg6A7xB5qDH/t6Hlj3s
SgEi92pIFaygAm4DrquLeA8GsxM7NLyne1dGzvcyzWHM285uN9ydFzkHTVr3SGqu
nItaLA7oyrcP0LnQa+xSEgb0tedj2z0g41h8qycq/Un51N3nz22skZuXS6Hwaa/z
65W1qmjpCMCoVeF/LHV2YFc5UNV27sjhodP0zdLZ2HVGozkOZNgKeWT0iiXU+zh2
jeuRAFXpon4Z/5DUkiJSQaDEOqbauKaqAgZUU+DjkYDpnZRhEcnqpYZoZ2DjCrlm
zomlQyU82cELuy3yI6gvXM3WRG3qtB2MZjdchBEJxqurjJ1VAclwl4qMx9ISndgy
dNAd5QVhf5YGhNev5ku80Uq7RZGRczloXZR16hNHZaZ8pPEOt+W1EYSKucBj2LiR
deStweL/ypuKr/jgaE/L4IeCp+uqpqU0WrPYDCiur590rJyc6L+dptFJomRdnPN6
8IbI8zE57VHFHUfau6PrUY1Xiye77eim3uqLfWdFby/ulj39EPQiQAePlZf3kF+a
i+Z+t7XJNjG+G8gj8LZObRO8fJAudvkSajrmpODkuLsGm9/qh+7Wywckb+8R/shn
vZ7KifhAkPN6EY/uWnq8mdJ4wvrdOLNDD5SYVMYV4P9LOP3FfWv8FqwpeALBsKu9
bQrt7oJKSVqUR3Ko32JZ1e9Rs0+S/vZSTMaeONzOx9L2LGONQFczx7PyX1uC3m3n
vcXLapEJ2e94JedCWLXPi1vTREU8XML9i+iGq9iHXWiRCCC73cgw7+3JIL/jizLx
I2oTSlZt/stzIoHo0BITY3hg51IArLdhec49ffPOLGNEWPFe9DCF41dQOj+YRC2y
/pUyDy/5u/J37q64enxx0QCdlzeDd/fxPJSiU0JlLjjdifAcmwZ+KTdbYptPddP2
Msrb3nOicWwEIo8N6KlfG/ROIX/DAKavZH3tOFVDThi/P6Ql99veljBVtecKdcPP
gs76W4/OH0pv744x8tvCjajBoZQEVCWQe0SLYTiqvvHE9zEbFOYbXeYyhDh44kUo
16oyDLVDYcMUChDq3ksS2XSzKc3fEmFsBZXEnOU1mcQQ5tljDJK969O1ZiH8o54Y
q7M938pugYukelCQwtBcByFZcX12/Swcji9+GsLUziI+XUmK/w6Gh91TM487IGIp
Kb5jjkuvjRpuvRhaEw/paR+L8tBArmoo6ZIzsDvsie4QahCdu5q0v5hJS8GBKubv
o1Gj8S9fcwUuuB8bTcUO2HqEqV2V6h7GdusCdIrVZusC9uv3P8J3H7HcO+JP2Ut5
ceVuLkH8ts2JU9oHra1uSGi0hY4FHrqoZXZowrvsaQC0RB63mha6Wh7MkX9UI7gb
BgNP66WECFO7BQfxO5wAtbRNxJ3eqHwgLMBlX9CwRYYto7ML2pJWD9/bKd7tG2L1
5FYO5tN2NxNvyD5V53civIlti2ZvOLeyhm5UI/PXBWd+buhmnApalLsCj2cVsOSi
pYkLC9xeuvKr2xaMm/71wFEbeGgbHbczgZ97bcDQIyrmn4sB8unPZFRbyr6zhLCo
ZkYTkhyG+9t4iobiVGI8mYCUd0Mc6387aObVxWKhcVhvdzk+yiwoDaa6Id7U8Ict
J+wZ2jdcn3ABHrfWf+czJouISMXPgvfbffqAx47Xq/Pnpii+Gk08kmyFJS5oAExl
SaKzDseymSnFej7R0ntL/MGcQpiogULl0o504sPX9UE1Q2YrBNDGwayWrenvi+ak
ZTndleDXUls9kwhtMPKZGePEf3z6aX9tanDB9Am5tbrfRvh2jR7sbVmD/aHRYSng
o9ZG8X/mR7YelapuI89bs++pdMHILj3yZO2Oyx1o/x/sW6l8odyTglzSp2jJLoTG
BqDm+4iCP2+4nUM13alp9rNTKjvCJWbZ24fknVOsPYiJS+PLRMPHrxXOAEiMzjG8
Kva2zzXTTZfeqBcoLu53TzxZMfNJ5Ng0i8goiyIwCY6aNsnzUaaklTAqsazO4J9l
jdnbar0J5y1qS95cKyWlu+OwxTBxzSd5v6XGg7COX00wTIf0b4vQ/KeOby5SZZBP
aKlc/NSarcKQD2RsLyzUz3ybZmzqFxA3AYUro0URs0kf+sBLNTeunSUoETOa9F94
ZBkqKIlctcizSKuqTMzSgiDVsm9qYSwJs8b2DDRE6FLZZmMdKGsTqNmswYWN/d5M
L6EcIhhCr3pRzPyPYm2JCl3+2Flhmjqur/A3UsVLpbQ1ZrEvi2jh3w4tNgb7zYSB
2CGWdpFijegwa9PXpmIp7tOjt27ZK+HBrnUPe4ZMM4gqg7RLeCt8iY/QB0dePhrx
/nLLOhPKhP++wzehWAAwSQaBuE6ziySsu5y9q5Pdgwa/gOq8aS5euzuuGt0VuQUd
MB0ymaknjsi2Yl6j2kyiJSpSjKHByITF2zRjvqGffvtKlBIbq3YHROkZQLt5nuCa
ycTTKDamvH2sZV7xtfelFJ/n5BBcfIASNCTAJR6XJL9VGHPC3aeOOId9mRMEcg0I
fDTbBstY+6ViW02Exg3d2zbvb05d6xxfJ4PjIY8D7Er26Lv47/RoWyGnKsqrUp+v
KLbVR0qAHy6zuCNMEyubKTGW2eNaLSTrVS+K07ViKVAtLNiHp7Yp2SzpquH0ucn+
FRujgrQs0v+EUyVOCs5uXvMESlXIC4ILUpKdfYa4vP03xNRMAA1noVjkE/kACpKf
K5YdzwzPTphtbLzseYP9JqH6ymhscY2BE/Zv7IXBg9Oyp5HtqnNB4ocRKYH1XGkd
So5wrjmEeAHtWH2rAofWH6sQ6U+TXOovfKYZ4yc9n4iRdHGARju/ReTZAhzigAHS
bDoTuzJBJnyfEaZpToGLj9Vlx3j+Z8YRoAes9cucRkMiGAMLgt9qyF45OjT3Gnh7
4MbQnL4phUd4FoSnh8336CncGlJ2sjD+h8FsPFneBPJ5ty4Tnzy552EHfLRK2Lol
oxP9bfZtvuBRqcoy+TDWpYAy6Ol7NAo7G8C6PAdwZRTJGqLZMos/ughAump6T9Fx
d2UyiivwK/iRM5TlBh+Nh68xfeq6x2NjZtRBxw3PjKKIhmgOTt7Qxjjg7rRoDQ3t
vwDz0L1I3ZabtmvIqEvbm9UzLjI7zvuZ6kf3BWshka/+JPgoFPE/QmVA48KJVkV2
EGyC9C/Qoh25uu4tStzSG2Wn4GcRCj182TpL6j/QCCfetNzE39ds5fLtkuqa6+9r
jRkprkc1i6EhqQ1AUs0QiBwy0ypPnW8imod1CuXOvhAy1y2SLyEszI1O3CeVvXTJ
W0wGEm6X1bOglXK2uwdsT5l4Bj/zZ8o1muRZ6+fEY4oevb/vD9YBYYegVaJ3CSBG
4Cz/7RGQ5TNc/jTkqFyLjCMJ32hisB7o89Pf0Y4OcpbIyFV6s0gDJgPakJWE/BS/
v3ec6WtI6fLrf+JYGOSkxtXgRq7MXFeFFW66KneV2yrhMxNRIK099f4d8rBp3zk7
gl370AlxM5K+cQ5QuJ/BIavYFv5PVKvLk+Q6ftk3WN0F/GdgpVM884xjWtB+QqPx
yX4PNBuliJz9fBDkxtx76BNsfe+iXwJsEIIrCIGH/9yMomesjDVpj24c08nhLPh+
pd+mE2IIIGKbULHpTQcRDc9cXMzYO715dT53klftoniz7K4OfDv58xHaOAGlXvTz
xrltQoW3kZxUuwzYAP7XSWVhvl3fWye/V8G+hgemPAeacDT+us+IetQMc84XoUM9
jlJuvvNfL0FTrztFnmXP60mb4G8lzrOZksbS7aW9TSMMshfIkRjOuUa1/s/2Tzdn
gX8zku2UEG7N3EZSF4/KWOMiVd+w4y5B7Y/fayaj4FwU+B/pEGxjS27FonRV+J/N
GiZ939jqF8NHYvQAySlOPjChUaDWg2OBbEtMESteczZFhIXFeODKy9zkFtR7JCKo
17OMp4C7jjNGe6DOcA0tf6Ua8WH0TMVnS13c6zL1HsKWgmXFPAwlNpnf4zp3JlUD
ajPldIVGsV64b84FtY7cYYz9eW0oSsToiKdu16z1hX7KRaY42t2hWwEoOtitfsVE
sjlgybc2mmH4WU3HkL2KanK04LkPXPZshBJCDe6O8kx6JaVDh7P4YeGbdxqxdKFC
Sp5cpYIxUjt83vs/d0bEFL8KSolN0AgUtMift4PjoapYV0pjnmMGN8ZQJJ6LZOEB
avOXZtwL0+p1JuBcXCv/rIUamBpHAg04BjOOzrKMJhDOIA6b5bz9qRz3U+nNtMZp
HOQ8impdKhYqkl37f8kCpecHqpQMEy9SpVbaiB3O4LATt5Z8bslncVgUxLSehJFE
1jOwNjcSj5dff0TJJlMSOw/E01QBmphiyFi6sMuyKN0mr//c0RVYNIWEbpZwgaJt
5SHHLRLRtn4rBo2Gl3+AdeGzo2CLTJZw2zma8tCrX6wzZ4Yx2WW+yaddTAoBbvi1
IpcIq83skYHfUREoBGjIJbJQJuG93e8tj1YE0CSQ3hjt57updz/W5vl+lVOHA7E8
J6WzDKqknxJah8hEaV1Z75qUlb5Q88XnRQZtHMyIVNZjA8mIiJQIWESTQceyEdB+
T4qhgDhj1BqEQwr5we+Mr9KLn5YkLhbiXDY/lWzz7SOkTWKnfaI2ghKJ7iW0G4JY
tx1kV/tBKMZGcY0aOuU1gbUlB73KN5au1e8HbHTtIm3rN5VCOmxwppzhvY4L3G+k
ATA7GnLx6o01XpRStZ2HLdtzkhmTn2l2uMqF7eUb9hEhW3M0/m/qffrF0A3rGcdr
0tYcrjMZrzWAnqd6BdahYWZ497Hb5RflihfFmlskgx0nJugZM3VJ/n79GWIOKA+q
wOcM1vY8QltVEnquy97BS8ekZO4xADrg2kiJrwD5zhUwuQxBjq1spdXcFyTcy+h8
8nGxY5kQ+0DVfyScpYv5Qc0cFJBZ9xyrM3VJVdsQxTWbUOOMr6KW3Mdoh7sbNy2i
X0lD+udqXJqnpZcel8h76ruOCQdWw9PB0Ql+kLFC7FMHFtFxxGLrahnNjC+4qbM8
0RyXsb3ciT0mO2s4iDRYAeZTfvfqLvT8A6RrmsffRLOHwTnV2c1oiQm+bjX9JTCI
ge1aB5HomcAVEj400NVPgb9DuQJullfpIVsyBUxproqvEMeWBYIjfj3lhdgoyneF
9DfAC5GKbQbQ7SUq+w4F28MzVqbMtBBuLyWe+28yufILA6V0dQ02k0FhAEwvGt4r
MW+8k8xqputnPCzoBidbJNTac3a8aeunIu6wvXePnaBtCdzuO1sD/6MPsyOTQh+i
iC943LHHZ4KND2dLrASs0No/62EM+Xh/1V0+qml/w/LP9VqJJadew6EjX30zgwWH
/YRmKblwbbTbQrEURdLY2oD3thZjy6cpkof+7o2XmOERtB83PGkZK5Vf4RO9WRej
+4rjSbVmNrDBLIuMYiT5u0yycLUOvL8cpgAVl/J0xYSIwk/YXI4D6+AM7bT2kVC1
VEboTaeIcc4giAF7nmfjFVlCfSeth9rhWFxSOjhn5cotEO9Jk0C8TbSBZICTcsIK
4iTcaI6IGkRo/+AXjRn8Q/hJmMJSDGVDvZsKv3f0PQqe0+/GORc+PqJUKWrBon4b
ATDvdHhXCsWiCd3dOOUCJzF7OCUBVxfws81R8Yxe6hUCJscV/LlNpXB8WLfjyE8G
8uqwR0PmA9B1BrIyxhP+13fVB+YaxgR/3jb5k8r4WGm/XCLhJafsHnCi2VlkGTJy
xkWPYFULzrfAPk9ijCnoLLP8wAzL1JKVEl0rC6iHZzKR9nLTgzifvvHv3+f7KQLB
/0VguZPF2wUSmL4YN9TYPjDnaPm0IhGstzMfWdVj8K+A3xmPPGa6YZO2ESGPFVa7
6W8h0+z3rB1j7VFIX6vzXpBKj/lNmYvb/B5XfXolHhkQnYFXE42PGOB51LNV/Sw5
sQTZUwBPpMoLMKeVogvfAE7KeLqz8zqJ7Tafa7A9BdtkBZZtF0t/SromcwV0U4vQ
y5chsIMM+cyyNPO4UTrbD6eg19+6jNsHPAjWEGyR4T+DGRpJ2pGt15e0OzqT/YvS
Y7ovNyrTc3wtp5d7j3OeAhby+g5MSkdpIi3xCSmeWquMDO6hE6DLGtLxJMaDOcSD
uIVjPaiLNJGxnVpyhech65RcS8Nfn9FxjBeLuhpLExrdoXqdVzBp+z+j9xtp+Jlt
K9ZNu+goQnqrZ0W3W4YxA7utmcfVHs+uIR2bDWxuDS0pvp+3aB/kHIEEZA5/66m/
4amoZ9wbvocEfSLyysOlk3aRKQtPIjID/C9iWAaIiokYYvhZaR+c2DEURtZNWnuI
FWBL/riDX5q6h8aFqfPAhpRuthTNB2hy+bjM+PHka0xL3tbzwecOggScLPC3m+NC
f4AYPNFXKFW02ez1zPyZieWzKoHzxpB/9ruu3iTsban1L33qN985VxqFDwFN1D+O
1Pg/lPboqr55su0PWZS71bg5hlq1mdTIBw7mHzK5GMGooqJ+aW7X7PdTkeWMExUx
jpAVKNJb5bXrSRvEjxZr2ptomesZUk93Jw1acAnYy92gJds5vgjXJ957zeWh0TxZ
p9zoXnuySlC3EBK4duHrbF04FC+gN/taXxhtsSR7Q9fXFUumd7SnV4fMnAFyiWoq
Qjoj6mJNaJi5Kat0K10OdAWBErk7XWDF/VZeXeBlsAaNKLCzhcUMwyrCht82vWOK
APIsioNY/qyGj3hArjpZtJVONgNfvjyd/vFjfHX5t5WSpNYlkrygPOE5PNz7ltq4
km67ygmqS7Q+e/BYEmrkCVhszNCOZ+mKxeQPmwm7SbyqbFjtOYki5ykkV9Fx/19t
eIVrsCT3u63AbTInzzLhMvjf/Sz1utu1TZKzV8ZAcTDpygnlflmxBQXGGh4TmiCA
UFFqErzCmVhpnZ8c0x8zhI1MzGZbDGA50b4pu9Nyf9q1b8MuCLwZvaRLRlQU2ip+
NHbwJMgx+jIBdjHsF9f/UckNki2wWtxpYVit7PjsdKtTCieGhM4TikwUOONja9+6
L+LR7Ymo22jDywMOyhT2H9yxikil4BeSColI3jB2f4QMMwg6aldKQkYTVhdoFiTg
3Pnij2oVcvUWbBLVfID+dFotnYMe2P8aFUPApJHXOuGaKp3wusy/zRaLfILyKT2I
M/qje0L3rDS6NPnP6V36SI8VcGprriqbAY55MAfA2AYJoWZ7FbRE2nmwqOAhDVhw
LWgprC4paNS5xGEwhDDSgQeGjz972SO+awTpqt1c6BZEUXeTK5YeoNgJbGx+qLSo
UwG3GGzxxEJGlT3TIBSeEPmYeu23iOXBitjqgrw1XWBpCKb70wiVqF1ai4tcIW+i
aJfj+jvXy5oQLf/naHUkLZN1LlUj/b+w/eMp5aitK4w5iHqGJaRBPrkTQTDq+j13
Qg+VngLYENVihYCRACsDSDTNMXicKC6g7mk8EyyLauI3oLR7/Znz4i3HdGU8EVw/
CkvxwtJCl1FzCYEtOAAygpAYXkKtwnFC3DsAq5a39qNeW3goga7RWittguLr6O7W
Z7VdU932GGD2/vh6bpkYEcNJXpt7UeWo2gQuNvi0RBB7BekJ+tWFqfTyuPhsItJX
98vDrvO9keTQHv1uvhXTW9BBz2tOh3AhWSy7iBbRMrFjXPodB/RevTQXkV8pqNAv
wKd3p57RKSswYc2Y3Za1lKNiWHesL6TmjGhSoQileTCJIxb0VUIm/KGdj7Q3isL8
OiD4CBlobY5c0L1HdEr8cTTT63yDP4h0hh0ETpVuJDb67Rhw/d1xOfA4TvAtDfKe
+wAkS77EZGp2SdSToB7FqjZyfgXnof3vWBpAjLNsnlsyTCKNWTeu/NZw5T25tMft
N8g5CGP2DTiiW6EigAgHW0PgwrSiWfk4c8KbjQukJyTPL5fajKPiDNx0VUmbzGRl
8bIloFD31+Wm978fj0JoLonb377u2gJ8Wo94pVVcGzczagIG4opeP5UKqhtSG9+V
Z6aKx6lBnVuhUMPHlJ2MMuJLiAAqgZHmenq9S+6js1za6+MRmDJBSyvJlSfPmo3E
dG6L5oySwbSDeMstJnv7njCBvh8mfqW+xUjmFTtKFYIL+4V9gNAwjsB42LlIo81q
875NI90rhvXwJgWPlQv5HX7Ewo+Kt4unlUZIQlAeG01Q0rzcsIRjQGnT1nx9R1mM
5o9j+hRGHDS8x9sOv//j1buNcKzhJVPUoSETjR0EnV0cVDbbH3JyDae7fHpsiPP5
0GAFvBK81BQ/xYDb8bKUQVtDIkG77hsmWy7uzOSmKBesqYRFprpn3iuJwEgo3RJw
Hv6hhBvLBGJuy017H2kTJmPrIRfMkNE2ONhEomJ4igzw1EGOZcnrJZY/3PpnDcsQ
R+cz3KXVwb/119xm/apghDVMv26WtWTWiveW8UvZkfO4EBo7r20Y9dEmunOeyIzL
njPwfOOp1WAgWiEjH1CUP6hvAHLiX3jW9MeCor7moQCoJCJWasNIUo1fjYtVKUU2
JOCBo41LAN+6ErtRwta0GBQT6AMie1825pyAkKFOTwrL6Z4JUV056wzwAUUmkoiC
5rydEojDmwtoMU/OCGuvPjwYrzXVqGGEJfulbSxhmQgoBIdAwck4Y7LoOWaLuOGE
g6eqWevXI8+axS4hhmFdOEBouEY0+G0mW8cbLzZ1tif1FDREMkIvug2CDMs3r59v
rfeXtc+vT09NttElYtCq4wdTDazYuHskLc+2aaECPoc2oIs1Kiq50YEECGiUUmh8
Mh1YQO5ZUcJ8kYeFTmwnjOWmoMdQIOVIfPecaF7PZC5Emk7l9g7Yd4dgq2NusIee
Jhj8eLq8r48QCC8iP7jmwgp8Y3pkA+XgxkFRtkSklPetggAafW4Rv4+TewLtSWiG
YcmYvsMipckVaz8Z+DMnaoogkC/P6k1k24LScN7WSwfAWcvNCI5y5Hy1BZ4PHGB+
mPKX7+FCvKpIvNLS5XqoZcT2QxXLjV+SEB1pjbB/QxjV55UqGcgnxPwg3YEVzTaf
UYyudeXBrphiVFqiBeyYfUfEH7Z2WUKOn1DXToUdM1WWAISk+zmfybzW145qRrpz
+svEu5RBDdpGyPHLejR0bdFq0UXn/R2B11yKobfXq6Q7IsX83R0rwezrYG7lnZbk
GZ03Qj28l1+Hknl8T2x5fBMD5Wt2swPM96qU8778+4OP7LTQvSh2qAKrX0vGFR8q
ptl6ajTpuAP4dO4KcsS6SWgChuAS8POkccK3i5QkV2bo0NgWA5iKJOlFovTa25Hv
GSY6RgYIRqHztFO66Gd500jW7qYIGFJJnzv5nq/94OY1OqrwGL6bumG7Lx8GoceS
bKtKmF+VCgGgHa4F7Qs2Phv35l0bUovteu1/AqL0GD3B9nlXYsyQ5co9iHKIDp9A
UEgvSMtZDLZbJDYlP+doowZbaJPfe1P9mYz9sXdzdYGjjn0WY7yIS2/A9wI10e2q
eLvKt/pbsjVBt2DSHye85KHtZwPjdzUgKHAErTAEyVJLfK401Xcfp9XWbhLa8uBX
+tQgtCue7JzJOW4N1W0n5qqENnlT1/pvyUPhKwapITUWSBmjdof2QSw9C4mgsNKG
nHHJQo9IbKGgt4qjUI9SbC36xvJ2WtbR/RYWobKwxcp1qmt6a4mV2gyTJ+/+n9c1
HDWnGwYyMbkNtIIiO3KN93YJaXsHVjKUvpQ4IP0KaFTv5ueOqOW/qN1zRqk0Go9L
TBaE0fvQpZAW4TsHB/dbGs2/53DSaxaipHwyW3PujHhFwe/T2hXI+B/L2mF1Ltez
fGgOQPy390If/hpIjskg5nE9g+PZrz+JUPRotWF4eaBudv6twKEvmVo9uZXUoOcw
8hx/I3fZhljxU9cq4k2KlDWTOmN1t/mSUU9EyPwuiXyWuVBWwrDP9rRHwhOlLRII
Xq+eF7ilifvIGS+fpq1UtNE+ZCKeHuMy/RHNlDHYXkiF9NBBUmKqmbCkxy0sbcFt
0f9itK3WlvLDteWmSMlmx+5glUZcQ+dYyP2fUx3msvlSmv57LSV/1D8+mF+ey4h1
M880p2jbS2nNXhb/KlcolZhV1c8l+vaTm55Z/6F03xq0HabnkwiRtA0nCAxN2Y25
a7tT+ykwxVNQCApQ3nmTRBQlaLnVQd1lYbEjWG8GbH2zf2YwlocPj4Y+MJRaZ/Bz
cKTaXHtPN1qAeKchkt+rchXnzlELNKGymTwNNfn6xCHYi9peql8JxMSW6JxuvC23
OYH3mp6kw6Mm0jQPZ/au4bEma38ETR6h0rHLio8k6qnMZhb+eQzfZg4Q4IIdyGUN
SWYAV9Ax5ttU5P5LVVjTD2k8Isn7pYnXyZoVUV6LbsJDGqMr0iLPSOEh1RoIf7Jm
oihc8R9xLAHvpdiIAx2alfJdC8m7JHfnuyfSf6jH8SAG1cAO45sNAzkt+TC46JPa
hDs5j+OWgMdtmxxVrqwxWqRuLVA+iue0Ev20aChjD3xlsJ/1p3WckhLC7UI7yn5o
In3Y9uq0Qe+FXAP7rXHKHvaZRm1ZkzzROrytp6pAMkJzN04R9lOnUwOx/B+orIlJ
00uwhEbgzKT/cTtQ0PFlyUtzpYfFucxzb1Fo2HF6SbfUDDaUuNl70mTrbFGyE32t
SazA8Jev9Yk8LdeNn+o02U6nOOXwGyU5OvCg6UbOp5RcLmEcF7xFx7HqnR9sL0uO
il/rg9jxzugArvWLfQ8Wj2w61Amm7HZnUIjLCvgAqbjlXJmoc3o6tVugS/SGYqWY
4Xf7eT6VLHRzzcVlGU5juqEs2GnX4m5Z6z7K3SxoeG5ShameY6KFZAwUsmLZ1wdt
2bBeiJ1HXimhr2QdApgW60hT67QheboGR8roDMCmLhgNhkceyuQSRGDrlda+uDby
uKT6zduepmbjB7pfD2uZSU1q4VQebTzHFxYw3SVI5GuiFJDKoMMYYzjWwTY/rB3M
YTHzOQ61S9CGrKe/MTIagQkxyzYxt2N0/rCV+lqNz63zgDeQfSQQpO+gYj3udTlw
WjeAdidqZYD7WSsWj05SKeiW72Eex+e60ixXYDdOUjPUX1Cm3v7IeP7tChZiOONQ
P7llTH5csslOgRrgHsefhQEpWYfEyIJykWYuqBQ2Xfohg44ndxgDkmeLKz1O6GmO
bJhgOaQw02Mo0ETgmEg9mvV/2Yj/svhAtiAz/d7IhiMUIXFyRverbPbwQRRlxzgl
rH4K2rcI4AVpBxMW57RCb8cLeNaZCUAsvbQtmsUrOfim3B7vy7Kp4GqeHFCFIWlA
5n32mQjrP4HLLdsFu9dr5DVq/UZ1W0x9qXLTtnFnM08d7j4IsgoaV16Jngki1pgz
3pzoRS28tT9qzQKyu7Gv0KCgbhLrPdI8agELTzp+oNRPoQAyJEXZQoN/sswwvs3S
ywywN1CX1hj3w4zC3AF/RQ4zlU5klKeuSOAJzhwqCK0JdEvultmziLT4fjJ87ugX
w02K22cEGMvXpUk9rKVQ2MtwpntsLjk8Fj/v7NQdWqT3DSMN7JixfHnMxOmwJ6j2
ZmeBHjl9EfKHNk0A0C9xfWpw5lPPq7DDnfZeWgWQxoMjfbT3KGK1FJmF6CTDQ5wm
Mawmkc82FIARUTZ57ndXb6+s34x4qpHiLrT0GaMnZXZIOASodvEBzrLiltawrKWD
cT35n1Zvrhhs4Ag9uurYN+0+M36AqwhSWaNGJIFnbI2kBNy30vgOac0+sD3vOROq
jwlDBf2G2Kxq3xeKndvv7ah8zKQ8mUzppkyNKaUIAFJ/YgXsxC6rhmI0ZaUJOieP
iZYmIdt/mNfVIVOU3ullwewzylw32FVtZz1C0M6NoCsU/26BGCd/4HXG70NPYhcA
e7v015Vaai36untFh7Rp9hAdmWy94F2ti/PqMpneZxPRan6OOyTcnvSg6ArExmC1
G3BNCIvvvjHlWpDs2OTSrUTMnDeEtoEWzLqZQFpZvJu9kNT75dAqeSOE9cqpAJv6
nzgw6upUQByW3OEzBO/86X3qk70PDvcTTylKWC2/yjt7L57+5qWjwLLA4ujcFtDo
nYTCYWuN2wo6Yl2BODVk6XK+bI6u9qulVTskzcj3e1571+JsBJNXlChTiMgT1IPt
jqZiN4RTn219YOYQ4gaRq7bexTK7Iik+IlhFI5uFJ7ggotB733x4VmL2QQTZYmE0
mzkb57ambLm7Kr1HdjBgtE6ceAZJRf3r4XBujZBg4rPjqjgI3LgdY567LCRg2fkC
Tg+2dCTTrMQ7PwMghrEgJiS3Sx+I7W6X/KDW/C9KHV34/KbJxgm8IgjLvhBTLqLd
4M2rBxtkMsTQb5bBsmNGvRQRHvRu92B0j+UeHb0xPQjOJkxo1d+MgcsUCOeVEruD
+2BErR7hOhKW89ezQjU8SwCbfbzLyUxKv6p+0b84WNu4kh/0jQeBsmksKSR2vf4j
Agqn9L+JJYYyvIc/K/GUpgM8/V5wqTGK35xbJCqOpPBBgR0RzT5s5uqbDaqnWIka
7W1XkCiHm58MLAjMNP1tKMqo9MgcxM5Pc1Kl3u/uls6cy8KJWDRsUwOBRDpOypzv
DtR5kba9betCg579V+9B6tODnTVAAJD5KeQILM6nfeVgT286MHFIckd4k1AekkpV
VwI5p7e5HsNsrwfAcZsIsAgEJIxp3mG5vJzShbUd1bEwLNVt6KOVZMGvnS4zbics
luZy8uasIJx6QeZqHldMKbEkQNcLNJDsy6gryPIcrk8XBLmJUYc35epJUEgGmqy/
sv2rnxzIY3vuU4hohLJn6xGBRvixj4DyjxF4SmNJJwU0pQxgU1G7QJlXNSnuHGjL
lKAL94lpKeRZPeFjHzwQRYJ4cT3Y7HyhG41zO3e7mdu9hzB1iAqQPpXDnFGscd5R
NguooNJqG1KUyrX+Vk9o6FdC9uhjbxEbxON4rzKFHC31ExnLNv94ggR8CpoDOxcw
crSYFHlKR9dJnvcabyhjp55PZcQCWfYNZBAimjwBoWduhtlcoOWXaWM2XfLVgC6Q
nFB5UW2eMYEmVmjC+PY644Dc9TWTrrx8reIGv4Wh8A+K0xETV0dZnQyvfc8wJjMY
BsGNuAFYUaTklViTP2Kbqzn2g5WMZ8faJEJBE2neoLCKYfYBqKqbsDDTl7rVPjbD
F+r+HM5f7YcVdCvP3vIQw7KhE2Gop/2HHDJb2tpreSeo68MZlSotPrGu8jSoZ8j/
FDyFxvZC4eItBlDfn59p9TUHDbhMxs5wArpHca+lYBaTVJNPHXYuj485OsescmE7
pO7ac+IKQxXx2oNKE7Zr0FU0rOrz40v4KBoC5praN4Q0aUlcu94tCip0rPPu0XPK
mBJ/iSqPMn8d73Hv9CMAD99Jz42mZPC9v8aTBUwwikjSRGZ6vDjYAAS65AJSYP3G
UU4rqNZvw5ARHAy/jK6dlQsLcG52oflFvmsu1OsUricd1Y6pu4VBojMqWLY3Kvh7
qXltcsZ1x9iFMaLgpHQrHak695zP8g0uMvXUq7aDiCbHzW6wyE+LVY7r6jCg0zhw
fPD9dVqAq+xpWH7ttrhZGHFzj/PXET2zoE2SQD3tdzrWVJ3KgsuAZpEZ7Sb+yqlL
gT/+4tbAGCG5R9bBQb9AHMLtTkvbMIzXTEF/DOK4iujTBiu1eDpu7lw01TVf/qto
gQSd3RfvAvxQo++rWykK4lwCc8w1emMYj2VXTuwkXaTOUk072KKliBEPreDSG0/R
vcl/Fbqc0q3ZAdPw/963rBrGuczUGaT8fTNLWX3JG3m6kcQFNMZdjwlrMVxxHMxj
lJiFpROznXnRPOXNAQSqlcLNmovYzW5tCEPQ4gYcP4S05slmnz9UBZQgddAy2BRc
AExPXi4U1HZ4W95klWCqwz8hVx44WECW3b6PfPl5Y94r1DI8pvNBGhn00tPzUCJN
2KJZBhlwmbwg34WOqeTWINjK7oRVYbpEuEPzv0S68su8VySHVlGQcO4St1bOXpKA
x3gc/OcLKNvdfmoR5McYCp85b4y6f0BG2xtj1kPKCN+QYxJNPxy0kYq5DWnqnTLQ
36qZYZRD/XAFVJWGhLGRIkg2v628/Kphlkt/Old6qHUrlPTeH+kfrAwMyP0upkRJ
SAjNjQ7SvZMxBRiY/QgZyu3AYeIFuQinSo77mKyljXo1L24rtfTOrSJo83RgUdQ1
J90ZtvbsLosxHJ391eDVtIVLTW9g8aU88C6E2Qo1BQyv3/phdZMdx4ieJfQAY3xh
R96YyAKNqkuQtXsF7KNCvhJ62ZWYRqW+YmCiU7PWP1/tcmIN4hX/44Bxfx+azzSV
rE5TuSIetkdaP3qjTH1haHbXRAC1splIkJ6bJ13BpWaGJ1dudQ55zPrF9DU7iidi
kMt5eiNkH5fgiBirQHK6Cic/XsId9jmAodRvC1fjCl1pDDgEbRd1S8fffFM36oMF
ppFl8kuhdvCQ+PCwM373+/FkW4pWxMrhr+6g8WHY9yXJNDZg3JFyNCfw7izYhpOS
XmZPVgALB9V33x+uSHETGATPM2cv8dv41xuJccD6JNnV0awj7ZkY4S+ncDBJd67Q
hGTwMYM2GvL03cz/hWnz8/c61Fh2rCApgeUgZBJocdm4oPuKGfpySaqbkO+U4pmL
pZNXPkahSJYdw3c5HCNcIk/KA3lGpMjWn8lNxFXpJxPsfm2fyTlAdpbkFkOrZz3u
FAiOJ9p6T4J8eIqAIyMrlvHSRnNv9M+ffFr248qzZjqxHVnO/47CAM2SdfrZaBiT
5+aIHl6pmv3rd0kIMCZarbNLZI2SxyACzdqphHsdBhvUe3Es+dyG/m7jj2JfABqw
e8YWkGrXp8V1Ntzf82OiWMLnzFFJ5oTtniUpsbCuZr15efktN8yu/UToaDyBWjMT
lCDxgezQchWrRPaaPjD3m4sxfVNNBvy0kNcXRh0jIpdQuiYaFO+rUmNnVz/UY+H4
95C0LOEb5Fn3FfR4iwsJOPR+eXYk1t2mqgNtSFGUWMabeVqHW74W3py6h7AUuGcb
Ur1iqMZ3amgkVIHprP/UDWIIkBxW6rK3/kwR1rWK0My0ZXVXosvwKxLHdT5Iwh/T
Dq63id0/va8hi2ADQfP3Xu5yG9ge+e4yEnc813rEPXr2TGZ1P1sEmpq6Y5Bne4U8
tYoQBughUJf32Nf13sD/tkNjuv25Tzu3cdYekwZMioUSMOqnRNki1uOdsBl8ja0c
iv5Nkeh3JddrJkii1sEckKWF6wyNc81TkT6N9pB7q/gMasvpllu6Sifeg9Cii0+c
z8UturGo9fDrWPkMz3+/OXShxC3GfNNJRXvhrohkWfndwJPmGMpDFcIcDTPGFe/2
17ORo8LevmRAM5Dm8agyJkI7lKlBysFEy2CnEKANbKlLYFHJ3bx+rj6RVwl2stUh
6UU/ZgW323b3da8NHsDUIKUdiOgIpS10GaIkna6ORRKRiIwEX1Pn72n1GORddDNe
4qiEp5bVJupQ7OMtIplzMLuNMOL9ZMM+sxjhBIcRKcuYYE0tNA4VF6iriREMxOEB
IsXH+HFU5qYSZGvDAeEP+Ovr48JI/WUyruysRClSdsFkSghlHOK6IM7pZPG/suiz
GKXpAI8LRopAeLX/DvMKzGR2Kv1+KOCShI7Iuk7H6K1vLf1aHoQCwF2BBxyyfTym
FfnNQap5aaIanpACFZzzVqRmZQX/vTcSMwv96tZ3f3w/ACZr4qumiWPkujRi/obs
KFWobWK9C++RNW1CtaSSHPtlp6DWN19NiFcnSGvSp/cJ/TcgLUF2bJ3vDt4RYGuU
L7Fwx4Ch7HvbNi6CiN9TF5h06umuha5JXiTYxWZ8gVfIzsRj7QR1l/eJMddUjTsV
ksCF0++s1P4u/C7s0H2h871T7jiuTjQElqY9x7crRSzp7nAZYPgY05TGYHiUKIPL
gbQc3HI7NKnseNE40n3qy67H/FRbwGHx1zBInvjL+pYLFlz1hDglSn9E6ALXFuV9
oPTR2gK+S7EUsg6rZpqgwdq85Ch43GuOTnWzSxRr0LS+jROl+jKs6tS+fiffiSni
/D/bKcHG3UtNvZ33BYqU8QMRiam8pTlIlJilfBURx0pSlXaXCjgcQTtNfTn5Kr7j
b4Xtb6Ji+jyFauMLC1hHUY8WL2jKWXFfTHLuRwL2DrNNMHkHZ89hqeLHkA5hJ+ya
8i5RLS+NDihXGoLg512ay4WrBevEs8p6+TGd9f3b5sqdx+81kcZGc9EMFVMmqYDU
GVVF4oLW3vhNZbfkR0u+E1O6utSZBf3du+MtjGQecma4I142om+hb6kiT/ar1DPe
06Rh+2ujiQ0uIoz3D6N2QbDEyXFEyh48eELCs1RoJ8GhAubkJDsJywrZEBYjUhX6
wAXOMJDJgumKVzJ99UJhSXnmGBl3/8yLobBzbcci6DYEzQEwHX6K6jTf2OtxlOFK
skTYrBT1gaB6oJpLmIw9yIPBv3+RXposKxUU+Gsps+qBUemws54qYP9ZJNDXclOK
mheeof/SGBYtH1wGxCZTGZHDvlO9UNON5qsuEvzoXL6UM82jT3sSyJIIwLX/dKx9
eOdIIJaBWfL3Pajj2tJ6rV+FGvIzJR9MRA3QKwElqVcDV0iP+HnwHVcdKUv9fgWx
Sqz7K4Qzobzs1W7Pmp+Jx++j0XGvWYqCmfk7muXHvuZNiHtGE12h4HjvU8Bo/HWO
n+dVXXONXD40xb8/k1BMYipiSemWNmz3TxnSmytX1DFJjPORm8OmnL5i4eGRP/4p
SRJoyX3eBCHwmHUBN7eGfVo2zE+TBRQSbvxv0d7UUbZJXYznnu90FQ1oby0PLtwx
+W1fk0VWjvAX6fZYnI3d3HTcATrzWu94nK6J6JJN1H6rZVEThLD0cCf8fKXEqVjj
frHAZLXfjcPZkd+1FVfFCwlmBasEsw38OdUW1DHXYoquEeZmxkKAAsCp6RJO5QM9
E+qIqE0ndXdghYLZ1HPaEv06wabiwKssQnCTSF6261Zn5fxDUj0p8oFsH255CBlg
LdZmpmOSAMcRo7UzmSXZdvUFVsxfvatHio5G5BMtr5heftsi8+ibMejOEOurDGZk
xPba9UQHVAJogH+w2tYZko12KGItz+NARFoXMiZ8qoEXB8Diqs938S/+meJnf1ab
8gzFRx0KNRi2GqzxguHQjtSrKkAglAj+fzm0y2JNaN3vTQquo1YUmcmLMF7p239O
3G3uWvCo0WbUwDXiMAlX5z4p4qWWwQLSvi3eFWZ6bXwx9yMu+Yp9k1atJ5qbU0JK
ad32BiDWrLFLefxh38szKdZic1B2+MsnwQBPudP1XZTA8kBOMhR48Kc/A7qmc9IV
RX0QQ6wo1H9He7+ic9dtPn7BgspW1yE+fy/ttzl/OnPmpiuKbi0H+YWhoAWmSyUG
WIW1NkTA763JLjgj0BOKfyaztdYbbIEbq4CBswRnyfDUBS741b/EcbNUUW+15qsr
jLtxDGSBcUBC+njTkcsW1Ar0mzJIM7NEtF9MVpH1H2aH5isFYgua6NE7mWPoGF9m
yAg58O5QLS2s79/p/QNJAaecCMvgIceuL0fUfchwf1PBuqP6u3s2H8V7EguafNyO
polN0B1b5o5eDx7S52FI8zyScZxlE8Fb12fq7rKxabhS2cHYLQuperSvNUtZUdM4
x8wT9MY4DYGeVzKNGMqdUckZqZFAWc5eMK7L38fs7LlFwxgt7PMycfuTfR41GxlO
7F/TWwct5dNb9ibWwwYs8A9X0qMTG3NKAPibqamMLXuQS3IJdqvan2DMtKOKMD6G
js2Gp4XOgg6yVFIkJF7IAkmG5zJ5hTfmo9KpBwLKQ6F+ux5m0CiGgTmZMbdFN4W0
A/rs+P3+mW6wIVwGXZcgt54LTeMOxOC18W0oMcASeH1J29ITESiT9DBG7hw86dkj
QsWmLhzPsyennge+xeDo1Xz1JKok9MOHH3NNyJecTNuy1tnl046J5BGwfNpZ2O9E
Vrhq0BasgL8NO0dk+vvKmFapQjv24MCuX0GGVoGFpMn7kzpSu9HkrHdo1jcDRDTd
6QzxRzIViPi/rJa1tbWzwh4XTmqiWy3qXq90kU1YVgkdCWBIjzOXySWaJruJR2vS
VsRMPqxElFMO7ak8C310iE6mupynOsa4PKYHSBQZz3zdj33LOy8PQjul2r879Gns
ZRHVfi2zIfjHp659aLAsoF7Oh+n/XtVQ3KnRcESnQtnr1gBX9pJpa0uUmGClaWzT
PPrA2hMgu3d4GCM+9J9DG8QroLlLPZoZF1wNzewxzt7FotfFoEb2uJAGwRqOwqau
iPKz9AHC2vmaZ+COm/5/UI2ku8t+mUkGxy2/3v5eJAXOPxjSpDSOZDQ6SoNay16M
F1sRh0l3kVl8KaWL+KmZoRCjoTcNKhRMASYss9Q6vdqr4+gPXMUYPrkEDPqUxMU2
b857NI8IpnQQRgG9Tf4GmjLvqKViBgBGQ9DYG/xRwKnVycdFoYQxIOnsOvoCytu1
xTwS0DQUfRlz92o5bfSvEOg7QPmv1eg3K3p4YnOTTkK7r6MIZoY6htkW23QvxLIW
5YRjvOOu1fH3jGD1BKi3MogwmZYdMpYVbtirXh/j++fzmzIeGnjlKEBkxvbH0tIG
K25DkRtnARrM7iXb3eEQ22Kie/nuoA4Spp6LhDLLmbl7dd1sBfqj5Duixo7MLmD6
fCZ2hZl3qp3Lejx96sy+5xk6XtfX4DXUPUdXvlQ3hHimOf63TPOavU9zEpC4rT+D
CKRN7TDDU3w6XD0KBHvnWwnCq4yyg7P8FOyqy9eqlBnhyJWRyJ9u4Xt5OX36p8g1
Yg4OVrLFjGLnFbPXwrf1GtTvYgf9R1iNqHLDy3TirGsba1nO55c/5a+vglQor/1u
EXDwV44YBpVpp7GHziNHm/mGgoRGKHUbvBUy371lEbr39oipGl1q/I6pDRQ3jhL7
Ps9J8B5buS3CFAYAqEji6I/wA1oQxkYfEvtI0zG46xWyKEeNGsVWzD5Hacm5fNph
DV6JK0Yarmw3WBdfus8+ZbyXAHfNhFFQP6vl8wzv4ksfNv4s/WpB/kdPLxZPUuqv
W1BfsVfyOFMTfgqYqo8Kh/EUP8omZdOQ6iJKDNWLpz+b9fTmsWOFYEBPyGYuGoNh
Kj5LAv/cWlia+Q9XReLfUi68euLcMbQDeusvgClTEXzOJOWVH/dT1i5m0Z7jfJIM
yufXHtB0d3I8NO3fyDWwk9mD9g2pOwCjWtz19F9hEWSQr1MMsXXVXcpOJe6hTxrY
ErBXKMCySbt7U0Z/h8FM8jq4+1fuoV4mF8ZKmqTIEOJYugKRiq3+lWoEdlivuz2I
41+UNnY+Tv0LyS6Np5sr2IzD1FlGEV7FaNAhxm6tYa9SFXQg+ea2eUe3IfFPWHue
nZiMmdNH00S2ESA/vYmIC1JuFvcXBaHl+ycNzEsqY756+P9XWbkRZPW94wrqZAuZ
/rZ6ayMPiw4mlQRImPVIYCKhta7zKt8F4VmrFhKeuiyv8I/y40HXomogvKRZapbU
WdzaSTCiy0Q9hUzeD6wBX2SlhsXflzrV/gFBBDprTTw+N8Dwz6Fyruxsx6DU1J+K
qrym3LheDYYHykUErnfL1H6G7ZdpBDsm0/vLJjH5oS9hbhYlWJLQvVnyx3n2Hf35
risBQnrq/98lIxaLo/A/rDZs0+78rumkzZ94Pq9Uu8/LnKwuKQJISgYnWFs+CJDo
p2VMwq8wB8wFjKmeOpcj3+nLUWP52GC+Ky/ElzyED7+kP5QliROCyR/jRZgkXnBC
leQtEE7MbqpdEsZYApPUl38t4E3DVEVh/s1S7bgUcK4Q6VyI0to93pOgkfyOmlGD
XNraowKbhA29A93NG4/uuz+Yigxv4tjxZ5XpLi9AcfiQQSrs43z+lQazEpLcJuhQ
i3Q9ZTH7Iqe4jHC5tgMOIHGzHo7sb3t+Dwr94fydgwGYGxg3THncZqJB/E/mygXD
KjnKC725HKKIWwFwVdvwwM4o0aY0VyfAif6qvChyLt2MSqAtbdBpYpRn2Cbe8V0o
XaMGN4g1Vhlk010ElnOkCBpAmN1KYY41ly6XHDCIWS2ajgYaAEC3JP7GkSfighcB
yp5iQ3APoNwfIP6v6xv70LYszop7vgU14AVD0BT2sJ5fQ+ShLZ8A0I77UYQOOVgB
x6zjRTZPEs1bzdiWdO5OAy51dpIixXxhZY1UR+co2ISgTWfWeGZNFdYXEaHqXBVj
YhA0paSeIpEzY4LvuarShjJdhMojRmjqMPHRRLUM/GyddCsUfwg2IOiMSQqrLwh5
qtDmyqCDj26uLlgvj/nc0ngw5Rl0iTIwc8Mcqr8/PLo7E7FvJkII6LiJicYKIBTe
ZCHAaNlhu/l3TxSr/sbyKeIFqDnu16fkFUX+of730KR7CdcxIqMhzLQl//EDXZZZ
qdOmisRGmfDDCbJls/rncns9rB1Me+FfdgmGnDlfsuuZdg2V3x7mYXUY3Ty5avrg
L90lhSdcCYx/4fAG3qhbqdMHqDa+CUcoi7Fs030eOSViq7JycAcQqhL8wiD+WSl4
8O9yYLwbJ8i7Jk8OkGa9m/gKkKnEt7hXksUFBWdCkEq6/v93N0rGfObAu+AVbpVF
wLlREMKs4oDxaEb4Rk1nhjQPjIqrjsPCH4SzTc8hp09tRN0/hI6FRIvnltT2gOn1
rLnzcORw1tA5rznbP6IB4+RodVxzgOQUNbKm/8KTpwWY0XsA5GrDOFqofHrvZCa8
ydyEJB8aE1Rv26QX1Hxi/yYvc9tG1MNTL4oLQ1Wl7+EIORN7C4bhROmYxZhObPR5
xp4uUssSb+8M8uza/ZGWH87cGp7QtF5WDfGJbf3W7mn2hFTZeIonnEq5UbGDsGOB
SfxozEz1nV24QWjMNbAWxf3PMHBFeL/sfpHxKL2E1cLKuL3QJMUxTdWKQKxPYEN3
pUhlTs8HxOpJV0tm/cUzVAreoLfuAntnwojTgwishnck/T03h7SRJZc7Vv7D/biJ
juKmGfvwttLqln/sTWAH9NGqmTwhv9ceIEUxjbIwEkg6fxfYcmkKB2WrzswEDkNk
zet74P3QDAiJ7dwA+mnvbTsV37pXwMLWxlzhmv09hHsxCSJjzFpGEu4AAHDBwI3u
C7LKt+WB0KXD2Lnmgxpqz8uHqNFXhXOtc5teLsJMU4TXbRaZt6uErFCjCeHEhfkq
xos1cqLUQdEDEoD0TrhANvPcrPioKPWFp7bCVl00kw9yOlueeyUN/aWorU2UHL2w
BtYW6rfQaiLRzxABmECKPZ1Y+WIjXPEtdrYrIWduwGXq9GdD0ttOT2Idy/z/nCvW
iZH4o3PHgrVRHi9C7qspfoJZqfD6TKCthNFC3IXNSXMWVXzlnFJNkM/K0neR137z
ccQlija3B1izSLSSInfQBuUwbIOPuaMZTeUtrAq9OO3+M2l/nZVGxCGPiMdjqKeO
HzHixt9Rrsn38sdY7VVChoGhAQ4lV6zxffsq/C/03nJnIGoriGMi/CUYBmN3zb4P
4+voBk97/4WrwUJmlqucc6n5KO5ZuvSoFa5EvY1otCpMCpjAWrJqs6B7pfsd8Pq6
WKpw+G8hiz8eRMZUo+WS4fK7jKR9lmhpTGbD2RGboI3Hf/kPwPwcFRsUU4qoF1BG
8WYVSMpjNidx4fOIZgViVusdo+cXdCYjER02PYVHMqvdqH8dtHKout0dLcu9uy9c
/6IPGO6m6arhkic20unaUfNMDS9t9ysnoNxEo55dyR8otQ7cxqrErmdYvPMR2vQz
516/Q/y+4Calk2i15OA/fQj78YgxGF43Rzx6t1PxbL7pKNpsVyYJ+AtqsWeKPmId
2dPgH/dHqEahXA5A5t1mPfsjRInfHcvpL4YtxwdkK7UL96l1X4i67mjqoPnWEse4
bimnmCaMirWKmMD2dVPVt2D3SpnVcBif7hlGlnNmQzB30c+3eQpKFPScNDbhNl8z
8d3SUoNhPhYg170Km2IBFlFkYQErgdGEWQzT6dRJ5FKcNiKG6BVDSJxj0umRl/CO
6142gTgtjS5EEbXU/tvT3oPL3JKY3ZOPua7xX5bFEgGkI6wKMB8VlBhJjeIFiEp2
3mlErkMCW8pkTPlLPVh2P/IctJLRI4kM5PJUQeMmeQUDu1UMFKDaYLepr2P2TVHR
tRFtT17zFMEsvg1jfk8gfVfFP7Y4KF1wR6TGJ7IvCG2BiGGPvBCYaaczuQlieDZQ
KSoioztPjJt2l2PuyEwDSvwpgvvovGJcxVyye/ayeQtrzsopYyHmJduFUgClTtIv
xcWZLaMMbvU7H+Z0h0y+VV8kOgUPJyK24NljsN9Glc0SNk9SH+HTilYsaXQ1/6H4
GcY7hndfmfkqi2GFlLEoiny1nmd60m7RR2N4yXHhLklLKly6Oveq/QrHr1upZiBD
RY/Jd63XM5emTyysNz2NI5ZcqKz5CynuKffgFWhHZg+McSJAy7pmHNn4cuYmdhsY
Ye4W/ycaoxtR0FKO4yC5ItbsiltLB1MJre/04m3Vhv9XQvPf+yUaIkhKNWaoFZRK
15PcmSDumQ+IybXQP4luO9teQBH0GTFaZaQo54OHsmG4bfL0dyC9w0zDuwlXlvkL
eNKLaiWoXollxo0T4GdsuqNsHCUzBs7OlLyv6ECHUoO0KmRdKsKZZGKnNdU05GPR
G2/HXsIQE/MqX4ZBtWQyKkzOQYz5jaZCb4017aOxXykKiAyqctcp3hufRTQHT0XS
iwl4zJ/txfuT6RTwZlvAr8MSwer+k9DzxUMm32v/cI/uN47isiOreZgkPQB/OZG9
hVAkL2L5fX6oXF53E+j9Avcl8SJd10pu/BFDB8OG/o08Nn5+ebXPMPOvRNgXiGx1
6Dn3itUyIpsQbbwQvZoDNWEBNZgINioCLZ6/iqpbfoTubHCw5UIODGjN8DVDtMnK
xQEADaOXcY3wG6370GvCQWhjFosOizqIkelyZlF59GAT+zpV3yYyrUj/Tq48ylXH
/8iEf8MDzXq/XoMGfe187bH3VjyAny8XixEu2qnKEllhduf0rJW0161DBUbHuFfC
kueIG35NQUtlQHF+wvCpz4sVYNCCN1T4AZKl+LHbSHsYbxd9rUXT3LcZCOXji0L2
ergMBC6vXCPkijfe2hOkVQciTWEC/7kgQI9zbEM5ZzdiSAo/zeLDJL/m77x7g+L+
hqaJNX3trGzCR8Xm0BccrbjPSSnJCKmYDJ+4xYrxYbT91xHaF8MBicB2W16GzK+Q
FUzkP5WPjykNdg494DuZdP1yaF0fub0L2pbYm++gwQ1bgibK0fFPq1k8SGbdcVYc
5LyE40Gt0x11kxIqCBp2qKCtag3kMQ8SK/vnLSOJklaQoql2nvjgx8LkUUnrzrSG
iTlK56cotPCgvi8gxK0No2fLo5nZlXI2/vh00AiqDqwJ1F6yGenZuYFWxWziRIaL
BeMWGhY2iC2ffduyyHclCZ/5n4YUBUq4AAeTe+tTqsLGD/Tv2gO/0Lqy5klfpNkt
k6OkdUf+3Y1FkKjwANNve3g/9g+18pdzFOtSKXuVHRmaqeLUsgjVP3jYi8GSsLQW
AgJzp4zyEZSXHCzYSuc3OKUZElxY98b/VRwFZMg0vqfv5rBmdgYYMWG1xE6sdbSE
CXmoCluGZfJ01lHPLhdfLOjzcNmr8JiaP9FRfWyGnKyilDocMD+BlKOxLiPzMLIm
0vTWwB+Nym7VyNMlaWFJWee3C5+Z07iv7fHbVszCBKORh11r22IGql2nLwdFCSny
rsFGrE5Apw+3vd5+2edy0TqKF3FmrO4zCr5U9eY0RvUnPWliBx1GuH769zsv8D9V
9sG9mom34HVvszniPvGFcrkqfz1boxkEvBXdrAhSNNIoesXZILxn47s0T6I+m8bI
GBYxZXuwl8JVCF659U6yc7cON3CqN1+Aq4YyuniiWixczhe+clh8YJidLAJaR1Fs
Rex5fD4cMthrvCH8SW5P/4/DjEuVZhzqCGtk6YEvuyxhcsF5CEWP18lmaPj7fLN1
t57DODqTrChZu3fe44usEzMWerNI4GKTMXNwsWlQ+gkf0dA+b0a9LKIoIaYk7ywb
lJWdjZBNFj2wF2NBh6r/uXh7BNsi/jqRMlJkDTUyHhvN5uEGrU7rL3rGfM/5/bZa
qMwv/mGqam34Da5pmhB/qWkKlCMIlwtclynAq0Zss7BHBYT5ED0iZ4Lw3dNBes8S
k2iSaUIXeyYsvAwIFWQQ3FdLRDwmK4X4PNLFqNWXPnjL085FfDB3IgPptAwt0rFq
W/SIE6UCU1JGup4RkJDCfFW4yFhzxPLS8l4hxcpH/i4g5w8QKkDZt5C1hiyAdPf4
l3REpG/JmvlAViRQOyxu+KAjZMgrQLiJrMFNU4i6Ug3ua4Q8Kh482wyH3CiN7kSz
qsFoPWn9DmOUx9juJG46eGmxq9sfwX0HrXwIIkhomey6xXDp6wkp9n4dr468//2E
W39W7P3T6AgyVq8nHZTfpC03yK+ttzQJUVywAy6qRBr76LGMueIjarMStxP4zjTL
bfYAyCGd0MthTiPEXieZNe4SgevMQMxv9qReTNPyCeB/Irtl37uHX7jDtc2KE1ax
+r4VsBQ+QWuS0LX7BKAwG26FTn2pcYJQy9J3jpZrDA5ss4WHw1laW6+nBiwhsSRO
K0Ebk/tNTOCyCUkQeVtXzPG5cRyVzN2KTIpAAem1/z3CCGarxRoxOjNqdM+/PZBx
Ma4kPAEpN/h1n3/fde/wNwdRBuRM8HSB+TiVgJwIpjRfxz4UgieTX80jI0emC4vm
GRl8307MiUSmMtaL2gjPoPpqI1Rdzre27Zzbde5vp902xkV8x1hyoLZ3IP6KvPSH
v9VXBlJm5bo6kEyjfKtjDTtkiDRQtAdpSXSxcWaL+BA/+PxLv7iA5lXX3kFrxuDo
O6Adg6n/QGTvj88G9cfpgrg3A5h+7kE1qIHrWjbNlW608yIPu/xReoJh7jaHm6S8
tM7qaZKg9OPOmS/5dv1nd5poZqJOy8RE1WszqIOJuiSQq/TkqFy61sVgS1acH2ok
4KdZooHAdGecr8xlubq514jeN3vUQQS/E9ngI4TpufOtd+5XLcoBtgzJKLzMoZ28
71pwZF1UWQke3AL3GlNKLmN4c759MbtRuad68YknguGLnKqojW+in8v2lQo0YGPb
b7e6NCxob/xR12BP9esFP97GfYd6o0K8RaxbD6Yu+xHvcwDx0JgJZBqjr2l5fcyN
TPb0pdFRcW3Sca8bkBVIu3z7Qt8kThH6UGY6MWEFezb0Dixw+iynsocnEeQJcSqc
5kqz91/ObdBJtjGjtobRFFCMAD0WGMpF7fZVeuxAApkeQhNubwjKFLu8z8/wFzdq
LIPT+HgNQeGRF9roeP27+xL+gZWRzmvvyIY6RwNDXRO/iuOZLGG+NEzMQNdiS9tb
uFcGT1pu37MVLQPNM0ekUcFnALrJAmbi9c6T2GMnD3c7605iCPSq6t33XwMu1pUb
ghmQQSaAsuf4Lj5RNA6YNyGgfeDOsOh4H3eeKvSVqkZbKabsDowNqEZFLwt3Qs8u
tnLnnRjQTD6b2jfwzlrgnMgAAqjMT3EM8Ra7V3Xs+rMEU+7jKMBrk/O7gXpwN9jO
OOf8Fr3JOQl8FtpzKdmXOrc/096djmGkplBg2hap2oOi53S1S0hFBVu4zazswN5h
HcJTi49L/NtLVbWE1h+Ptidh+nGpK9+u8iDTzsVbimESLy3tVaj9ggw4I6D7GY1E
Xa69j2Gxu07YKRUuJX9eMP9iNXjJKK/grEqCsY+8VN4E4EflTtpQxIqFNEYQ4iW7
JXL6rShQXkPWQEBcTut0JoLBX6NZZtVfyG3UcN37ypI2GF1vAqdjjwpsJzNlQQS9
rc8Z/KaoILQtaq0+huRDvSlewY1otyZUYZYM+9XOT0fgXSA+eOaYIiqu5pRpp6gl
D/QoLfknfLfdnGS6vtCbLtqDlLGcCVERv+hmCjvcMkEyB8Mk1+fUPIw+pFtCHsyj
1i+kSMxoxNGoUbZD+U7+ExRtTADCa3RRUY7r35wnr2lxw8iG3yyKeI01TG59TLq+
2q1gXxTd/2jozF72JbN9Y/l94kBjUkx5VlyV+eafgarfXutMAhTR9xsXcEecySwf
wXi4mey0Pbs4fxZzLt49cdHxz/VV58SGnfC1XrwqxJbd1Lc5/0edk0CudBY7W/yT
9IlegbelT5rHbuAW3DTV/DpgnuruuS81fzhl+tRQduuhnalfdhzqDA+kF9Rlg7Dg
bLXJpSEe74ESqrWyyyxRpGyke2NRQsg3aB+fx4zHTqwZppb82DO5am4EDfOuNtfc
aIbHCjKGuwOESioMddOK3R8WewDcvx6pIMNAD6Yn2Pbjl8TtWRPtHimq53lQBkM0
9Ph9VPYRfnYprEiYGEVMr6phsVgERetHjOTter3Qet5Fx9mVgTuVV4dTdj0iD2NA
8qWXbK0f+nBFtjX8LGQZMLXRtj5qtUj8np9zavQ9AVP6nymVB/Hny/sE+Jc/Oxsh
f8K7Wbmmw/Oc6GYPOUbSVcEQScQtCzCjiAiicA1nNcZzilbwcDrFRGZvMFVpQZ3U
UmCqPFHPKeU359ouEyNuk18vVbpJI/J/M4OYb/B4HB+yvSPIJX//g8rq2CxzB/Fo
+tlaKmoh2epHlgLySh1ta8S58KdGCmoH+6Iw98UzFSNqqbAnCrtN/kUMYrJLfXWk
WABdnksguLXmkx+Jr5dSC6EsJms94b8ZMazAm6s69K1SwYt8dh1WM8PQ/MDVmnHF
MfqEdnXK6tTEGIikSFJ1lH/vNYu7GUqySqA19yPEhnPGvoa05b9SDrxCc13KFTkC
lo3xS6D6L1kWuIUtHOEq39HZJQS9FdicCcqRjZc2YTBkwbQl1UhvpCCYPcVeC96U
TpobthHyVrpadVxXJXDcDRZ1cckVboq/vHM5ZsZ+SOosuAtl3ZDVH/UUX12hcAaH
X1SbyA6/roQTwj/rRBF/h5T97adJFt1TqMiCvET3E/0q017UaqUv9qRofxEvVcOT
kWDrQ4DT2Rszy5O2DdLwizbACILrp3JWdt0m4Oc3GvXnJW8A/UZZK9tvQ9OIHPPD
A/XvUuxZUM7WBPRGtyM8sXGerKVwnriis6wnF/7helbxgCf9tOuFJU57b5gtd1C4
AxH0FzOM3CGMcBfZ8boozSVlIyXB2V+nk+gHztxtRtV8fvye6xDnmJwP1WAm2Fpg
lB9042gS+aN0VIAi+2fR7QD23N4PefL0KolXFyYYrVcxlyjABF82DbTFWFuGYtD2
XQLgOtBfH8zaeDROUPvT3noeWwJAnWool6LYXRNNmv3pP06SlAnRu7tLTJ2/lX9G
VfupyKHAq0A3a6+Gmcljff3G5BPLvSLJqrYLO5SGq9K95xLwK2TawmoppZM29RSf
MyQudH71+Rc+d96rre4fZOVwfRJaTphoR0sQPRoP/nxVFf/epu4qd0IpdiIf5gKg
KtbDzLAnI8odWXpPIXdD0TWKdZgreruSEQSaAtUFy0mZVwwxac9VmGDtCGCCBTsh
rcoyczGdF79kQOEYsDCvh/LZLEOONovAeK2eMrIwO0Mf3EK63qZZ2MQF3FAOMJnG
6GrW+vBvs/kuOeJVLZcuuuysYItqXuiKvPvYEY4kJJB46CWiZiGbeY+FwohGbaNa
KN/tmM3QD4VAkGfst/JW9dMftetm7QqWkvivBfGnRdf4YlaXeDdUN1CT9L6Sk3f8
hqrWVuriFpdp/X53YKCdPgZhuODsLIvqR1vMrFYl12a2w/RkBQfOCER8TzWqyyq+
mkuwqG74inUACg24Xyttb5A2fuXDYOjmiIjPJOMy4QtctZ/N/DS3RBCYC7TIuxS9
4qdhRd3ldahrMKq7+lCh5NMxhcPHynmxI+IJo/FfUW4Gph7crXAVYNpRBq6SlzgM
E0lGCP/83+pOu2dAayhKm2fPfdbw1IOQdrk9TfNqCp71fjS9+eixJw/Za9mjBPWu
avg6sKV92l2INsfLFsbTJb9Km42SZ0BTwDTVPmIUSdEyOB0K+bQdnarT+6mk9dwb
s6dE2xpAIin5ZXUe+jjgEJiuUq4qTraWBkuUWTW/xR6JFYUuRw2FQTIvbvXLDyw6
3HtmURaGUevvtxUqnDZrRxHLw9/6EkcXw0tv7dm+Rumt8VVSMgdWIHDzrAteGegt
ro8JEtctsy0iHV+Jr9jAODJ3EKfisdb2qt+tpnDV5MtXHHXRueaV/E5t66p1259l
ORRWkgn7Tn17rSBWt+EgwIOacGrsY/2pr7dbVquiW1cY/GwflPUKlNGSvBsdiJAY
OgZBkfaKobTJQ3Y2d5uxEDHlwGIlssM6H7fiHDr8hzEo0v3/CXAqchVIStRxFBvc
kOJhu4d7ZB+hLwblLvCKycqgsI3VLjVmGTGzmtWMrCU9OKT4iuF/lCVOa/HbZx5r
FGKRcRwT4K3KjZ7uWmZieFfzPuxdc1Rc6cSX/OGVI+UtHfdqjIn3lM/ktFKbHFSa
D4zNOJMASzt5VbrBuZdPkFZLkf4EAs92YZtfzf6nr1AY1AeMUsOQAQABp8UzGS2D
DiQFfDaOpmOLmAJP7NkGBVwJBsisHvG47eTAtEogBA0yLhrcjC7FosmtVqYO1/xI
8I0rTkYHFNoLV/9NFe475L2qSswwf0HJDSrgI/j41bOlElREXzeX9tLYLtVGLX4f
IIYEP/rM8nv0Klmg+60SjSl/nNs7gQATHg3v33CEVY+457lo33ZgTbSp/OsjXjJg
yFfcejil+CXMyStw7uajNT/bGKk9JA2uH/glycv/29n6Fxv7aIgW/ua54/pn2QiQ
mIAU4Wb72IaEkDbNtb2nZEgjYx2jswB1dHEBXXWyKm3WbuBaT8Z7BijKNBLV1lnQ
plR/hQwtoCiW/qBuqP/AS8FkqYfv5XvIPSYrIrBl/v9yarYz7YeYFIAbwWPhkp14
Bm95a5fuUMo+rdrMHxT9rx7BZPUyQF9KhK4qvZQ0oSJEtu4UZ2+YTM7LGXz2Bmzy
muwDUmOXNxSL/gz7E9IwnS6y0Uj9fFLG0/0zPohoGdSYa5OhTToTVPbddX3wry6K
cERsm8jC6DgeYNbLjydzmaV7+Imz9k4LwkIENRhTOiuYbzcyJCuymvFWnl9rBbhv
WGDqNnWr24H8oXcreujL9615gvVxAznkI3hQSbZZCY3zQiB4MBCBEkNKuaSWqx+M
SMytXQ0eA0mNChTEH9lN820G1xCXWfNhWOsPOIIJe1FmnFE7liUj+xr7sFLj1+17
z/G1E0HC31g0a5m6gT07bxzp0u3QFHxPFE+JZz6tChinOjjIKtfzL997z6r+HcOd
obXJtO9jAdWgIxgfp0tcqUn5sOtjSAg7us+9L4OjgRPkbF/d7PwKkedNuSX/QuNe
0TwF93lFY9C0yo7k9XKRs+qTd+4+jJvlXhXXYon9z5erHKtDmOQorB05f+N2L3Fy
zft2Ak+8mBxWFYX+U3M86ZRWIv9sq2YGg/6KfA4c6p7bfr9Wi7x+UNS2qURW5Xy8
hMFDj9f9KBTyeyu/ldFhVVhXl+p8iGSOtzjIpCp0owLLCOMR8gNJAi1UJRdOmFHD
GmgenMrl9xQveoe3KvIqrGTF/uIT5IhHJgPjnf4WsEEGmkD17NTbKzle+ijvgUKt
B10CCBO9Tu4BcCLs/yMajNesZi8/zi3Gaog3YGqvMcH4Q8/z5YVoHioi7qDn6vae
WpKJgp4qAu95bAYQX05lyqL5ef5yZ4n3bRmd11ctODu8osVcM01GhbiOyxxMrLwE
AKxssN0aUWdLTQnzYgXFVBPY2i5aadDCjzK8IcaoMLwq92t8OSBSf/9soPHIb53v
nMNc9Kojmi9M50lXRVECQuv5gBZyBY2w7Ooa2inSEb1rqKfAtDPGjgoDydGVOv24
XN3B6q3SKBp/bTDhMkROHjQDKN5OWdOChCnNbXY+AnpH7UZWs3t6DB+3IvjLKque
weMzN4JYX7PWscoxbM9Em2Gbvq6p27+O27Bs0tqoCj3hLBhYFSDbRukRgB/xp2Dl
V+T3j3tU0XMTPolQTDc0Q1AcpesZcpUiGNUkhSRE2fbU8sUawPxoYV8ug93GNu31
yvna2/hvUmY/vE4eYAtECUi7FDzE6AOwSSNCCne+2Pd1Fv++VWooeorXpZcpBrng
D0dG+vToWT1C2L12CKJpAF+Tlndc2cd1CPfvGrEVMlaAP4ZWU1nteMwTdbevdxot
c79LekANeTfJH7hYmiEM7P64V4hYhOMclGIFATpBjcbQ9AjZZGWmh+QtkYdY9fZc
w+hcmhiecWjo1lo1pSM2QwHCWKpQGxm03NUSmUGrp2ZVz3IMZPF4zdR3jnop9mG/
u4/evlJPF03b0MlWKJb/ONdJSQapZlohP1V5xHV/20QoZ/dfoXpsHIkilXnl5FWk
oX3ZR/I41dhtrzWMXD/YH8JamM6C3+ruZV+Uz6PnuzzJE1y6dg+4gfKQJIMcHyes
mrV99sQiB4sfX8p139t+NR41/JWuy3qHFRbI12xXOpagcrs6mWWkiGru8yNgQEFS
KjVk/IXTQ6/kmnUF+ABVYsMMWxbJ/3eU50hRqVD8t+EOhoIfD0174zsf98JOcvFx
pc3USMSLTOuU+9t8g5ZZEULVHe0VvPM7mRgR9RX+ZzhPQw9dJ0VDUc7gJx5bMZV7
qte7U2WyehnTjf9RjfuvlpFFNDG54A8eyjV2FpdWciIm5AbXIvJXT7pf4cIyYte3
8oc3zbI2hAFcMVliREMnQkp/A8oHd53soQIKalehmIkRhqVDHTypY/zpxAhT2bgo
tfyq4TbT64GbcL/mY7tATPXx6+6blYWIsUCx2Y6En2VVO+SSxMDyFdk6KpxJiXbo
uOp4Uvt4q8G7r5hzTI4totcj/POCWKxIdOu/Z6eOaHfcpYfuXQL5MiWaJf9kAXDS
tRZor8i//ysvv9SYTF4EW7ikr+i+7OFR77LMKk0ri12f1IZV5clvBkAjPOb8zKRA
xYANKRr6ujHHeB0giI1FBzyVhUZLnwNZm27XYXMtleyfwShqBVQ/cFe1/fsEUPkb
S0LsksAvO0LChnh7LfDzcYSqs/EwBdqFFsPPfWhW+zn9SAh3SR69nTfktho66bgk
ur/9GrxOSJqAS3y8EdcbX3ty414p7Q1K/zRZrcMuPa/PpTDL6QG6kPsVaZP7cipJ
+lUD0oLjtBaQ699Bgiit9T063vzyJVxcW/dvJ9gFABjRnmACf6LeKJU4fx74D4bp
zNl2ccmZ/uYgNwzXYVPChG1IOze1KCHtywWuWaqzhEe2PfI67SXSM13QTVjpLzqG
b8XkO3o1pj61GHeHJFPfvmPkmC8o+e03nO9TTyUkGtMs76KDPTg3fM/udnNP0ItG
8WUyvbz7xgfILaN9H0pMx3nQFR3lB0DQ4gcRn0xNkzQgRuBm1ilWDq7b6TB3qtyM
dNUhTHG5PJVXLHapjEajeBQdsgRIjli5LK5ENURtypNoYJ/xQ1mdvfpb+gygA6jS
928qIP6wzCcvCnsvaYLYroWUuXVvt1bGYOU0v2kwL8v6JZIh0Ad95hQEWZ/OANaM
JmQA1ddZ0LsOsOXtPothWwPPdQpdfr3OnJ3oTKu7g04EPs+FcyQM7Pq/AmRwuv8t
PsJOUzcXWgVUof1ogqszcIKZJARXbAfjozAeCsVbBBY2oFhj1bhpb+fsebiF3HG4
x+2WvZiZ9FMNAD1H8oEpUoOb46UVBVFsnj6hzlB9e2wNwibsidf23vQsYTJzn0we
QQC8539R42SF3vd0yB/sXXS9Xy07C96MVwnpvEIpdKG06XV4gvcQfF/cJO4FQnQ2
QdKR4YtWDMq272DbjCuuP+KOCBJBp3c5K5cYPQBY2LhT77Y3bgjGiA+7eujsATBj
1/UjMWPZvBKZDPXIVgfgKkL1zz5Fv3pNUJBgMr1BJGszXDq9MMRfI7AksP434B1o
lt7XpqsET18NEH0Jyqqde3VzJznWFCHSnbpRTKUOIzBGGTFdye1TLtqHTi/ZqvQq
iNY/ljUscoumEDuGOec8+IchaMh3ANRSnOvDO+oMik1nvddtMnMqVjJ4enGnl5I/
ENfaROFTjG+pX0YAraJ8NRz9OiPzUo4l4ozsrZh2DdqZK3PXzD/Bx/mmrZc7m9m6
Ijjyirw0Cd5ppDPuBsEELc4/vZ7PKTgU8EHMEa4K/IsqIRlCA1XblcaSvenxqkQA
qeN0GaTlgknatRWAj1rsFOg+kKgCoQaDTbBQSBMbDM4JE8cJ+IQKI6ytMvcjobSH
nfhOz44TtF6mvj+9npps26eRff7foBaZ8wXd28h4FObmqjOFagGEVUh9Bgr23K3i
dms4YcGiPgiMpFKfictsup33yyhn1YPZTT80q03vQzGyhr0gf0vHITXjgGBToEEU
LWC6S72zbeaJCkLFlYAHbMQAPJZ2yBD9TY3DnUC3jwml4SAonnGti7or0qj2yBbK
2vY3jC1e83I6rohvf4LlfFtnDakVI03A08a1UHb+9fuC9Ln1qUj2XZbfCxOwMjZo
luacGGef7QAslyIgoEj+AbHKkiOgx4l3F1IZZFhq/FvZeIe9MclNjQhAVrJwdXaL
S+KebCC365m1Vo6JJS0oICNDrrOcg5CP4AmOxTDc5iJXEQnwrkeFYvEynVAJ3JUd
jX1zQz5426WHYaM+8Xfxtp6m4PEQfuyQp5QH83otu5YV7yuEeXHToFLHOBZIAkby
t7JdMTcnbJnXwdLBpO+CIYe7WYISxaxS+t7DRT4TZ66YIjTPQ6DKIo5bU+d04ot/
r5Bo4f1ivnyDkz/37102gXK/yt/yO6v7peywRG4d+jJJn7yJPHq3h2UMoVpX+X+Z
3S4b6lc1G9UGsCQbLyOECWrg0WcXvnmvG2Q8AQL00VBA23A0NXyx54uLrHwJUwEx
OZuCpCBZTi6AIXU5JNXRJUL+IhLQM4Bj2VhaNaqglB+XicF06HyenP2RtYOcrWaQ
ZjHQV1YWmeERyfG2e38x7BZvshgLBIG24lLqA1cElgwrb40vxHNMCCvwocXZvWAZ
SCva9Oj8DLdwAhnopVPVLQbc5A7k+BludaZ/wVe0jCneqCQB1WN8fvUWKxAV3iWd
tOaptwX59feOFiedhG/qQnfJNT2uKDqrzev+4fADkhYPF0Wywfg6FmfHw7o/+15d
DPX2CeDOtfZXr6Qa4XoGJb/9/9mYZIgrUWd6Zwxs89hC59fDwWllHqYP/oa9mQAy
8BojeujOdoBN7mudQGSzAGdm9SqXRTxhT7lQcekdawqXIUrYRPoiHWzR26SITG4U
VThAE+XaElZiuHdpLrU38fMXNQt0t5TvehYlU3GtyfT66GiDVbx+6/o6hh1NBQVt
y/eNgSIHiSCjEUnJv1hqTrNgcZGnsJ28ID3XLqTCzHFajNjSQIK0F1aesQ5yPKNz
V9yJnYkJ+FW+vmU0dZqS0+23BRT+XZlsj6TlCxD2HxRK9//NDklY6pAaIG5HpGsN
alkNUlhw/UdjY3baoMdTzrSvsCxWen6Hd7iXM50BTUEkUHKD2NGuGe/gME1jJbV8
UpDtgmuci9MI9UKdDUScdLd38ZN/oKCp9uObFxZRCc6DUQoxh4JlBNm9Oln7tyA4
vgpyQGPyDWW4z1713lFv0Eas3qcGzeKwcpIi/cZhchcz0CKudeNcfmmK0P8Y4nYX
3pUnSbIjsqE0C+isaYgIaUlbUr/sKLXPiOOIKvBAsCxx6R6Cfa6VmCUg1l/sRAUn
dBn0VorN8cOb8YYF7QMlZE9ymKs+pYVcstGHeACiNa1sZtCMDKBjQmrpFfZYRTLu
5umAvAvAZ/9NS5jFW/6YBiDt5Scp+4tYFZ1UwyY0gf5+DLgjRT0W7GiPyAAeoyIP
DFO8kTDAgQ3N1c9hbUnEMvW3n8lEU2TEkhTzDK2RQH5ilt3R7P/Q+6uthaw5nrw1
9vKcs6gemWw6J2UHTic+f/TxBcjBmQtCTHBKZLG+YnYghl3ZmoeM+kHvERA0iJfv
c0Wskwk15dNKvM30p7hBMcaFElXu448oAcZM2QES3d0BVryf1PWG7irnyYjspmcI
hTR/aUFMXgu8cw7D1icRNw+6ZM+v0VTW9mzdCajRMKi3PuIAXNrpHzEWd9RDXRmv
iVkRaNKbbWlzL/6qNWaWgFG1w3NWGT0cYhvywc06LTu10GQsUDOWet7Z3kG5LDwQ
WeGDmZenLbbLfrjk4oTOrk53FxhsdymQIYRn8MCt8Xos3eqpZKsACi9MIDMcNe7D
RFFqZxPFhfKfXtpSmx4IabeYwDBcpoat3q0x7GO0xNnyoyd2PsQ/b72j2gw7zT4K
UQJGvKW3V46IlKJcv1C6nDeOGrwx5g0UcJajIMc6W/l4wt4KLpDSnsjVJF17/nLf
ojVSie0k8GfWn7CgITEQHyESIdS2VfxV5DOXuVwWTrZxvP0XcBJ0yGkC+5E9Ux1S
9cOX0X5uKstPZaZgM/M6djF9JWC1/r381KiLiVAhR+0sZnxYYX43jD1ijDnkousp
uXy7YZXi4QXO6TuUNHlkT+D8dtxbWHugAL/i1U+n7uf5GEy3v2bUb1dPUi4NxvNH
pnZnGKuz5GtKejeZt0H3BglRlIyrQchriGQUEbGRo9rVFSkKIly0Y4sadgvlyeMl
p98Fm5TkeusUt1xAs2SRzEcaPhMTD79S7dLeVwF5lOv5P39k/1Ty/gPLCB8/N3s9
T4amYLLLE0iDYwurjdYDTyNX8WPyTnZVpNt4MPAFTei9I/j1PEkhprwBg6HtrDvm
lMiF0kHAdMnVyHedYG+vbsgPM7SXkQt4psOp7JCmy1ZLGlQQwqQ8aex2voUi9kNh
ZctBCbqbjz5T+okDqN0Hi028nsoXQ3MeXHPZTkTfq6ZHTk4pVaP/YlVRtS9E2xin
TF5UkSLQxYJhVT90cxxE5nTsy6hd288TjUpdLzVzXNEZXsu+yJHjjqtyVkEE89Yj
VLVnj2w/hq3z8eDT7RTWkfKH8NJEwiTCxXNIx2ewV5k+R9fhRo/d+Sa/CTQF/GJk
BDyhKTujU3qusuIy5NrbrtQuqQtUkMHyfXwJo8pIGn9xA9R7q8t/G+xryxdhjwgt
xCAJhYoHogWzD99KOPjilKLDKS7hj/RPoclv3Ak2qD/a5dD706NmxA39FWpo2Sbn
7iL7BFl6dU3Bc4RGApMqnnDZT4KC6rO0dzzAF7xY5WvFNJA/FRRh4bMii/kZJ39I
oT0MVXbOpEQn1WbxDkVrc7V2+wOzezOr93Te6A9BA0deG7kHObegdH3epoypMfnw
68zClTiJsea24cGYCDwi9oE6MoEJJztS+6ZSffcWwJifqtMy9WSPRXwt5F/vKbdB
xNX8cQ+p0PqfIl+5CQ5Ns1p7S2maXePZSL2iEJSHX7adhb+wrLoZg2bC8eTzL6rD
94Z5OscpJwvHl1bDxk/cl5+z1C8KKXcsPMMvORNAPnNlZMCf+O158FifvN1DrAOi
KBm9q4/jYMbxRe58D5LK4AZe7c0V7keiUN2W0ujj27jnYMq0t+RdxO/w6TOW4/98
iA2eo1gUppxGHTGgt0ljCfCb9uYZMOyv8IZUISGLY8eRVIJELor1byNI/UIFe1eQ
EQFjHkqmkHbp0aLXYKRdGDs6EP3nYB2S95opmCfkJS8zzvOkveTlN3JiJL/9PCss
ewTWLLjVyiPNHc4Fs4+aL54E7oSFiSrKczvqKL3UwDWqsJiRMTOWqUga7mLIVfmN
mtiV6PbQcw+g83iLo4iWAf/ErJq+A78xv5zvcaPiqjlhfcZRARF/7PdR0UPFAY/p
PuXzPMmqOT/jRDIwkQEUtrOyH8tKZHfBm9owggiynaFdR1u346Gx4s7NZXwjyJcn
ZODJWSIdN8sxQaQZ7t9uRIoq9SvQRfOb7kmavLrxdzEaYuZgFOJUFf6Xg9Cfa8Yi
2g+oKg8RkUlRrweiiIHG9wP5kH7enYaAFSRV0BEdALxOHI2HAtjPVScLCqWcXefG
l5qcYYgrDm3hVJ8ud9LSTVPWFP8CcNkodfh+dTWI1req2BkIjlOh9MQiJ2ftBMvQ
Cg/08/sX+2e3yhXtWyyqi71IesIbltiamw3wFtG0+06AUupD1R3RQvXEPe8/MiH5
R7SzdZfu0S0aQSwKQZdnu9bb2zSCjbE/lwOaCk1cYNoR7/RgqNf2Mj/ef7F6V0ND
oxlDeOSkbj9qbFVLfi4ekTby9T/bLwtqMziXQ41jQmqWREz/91pobN39bPrnJcg5
X8DOkqTMp3+BUQJpcY7+c8YrlzRfkHIsjgnMCiQ1eb+2YhPUfr2L/RN1Obc32bi5
ckRlTr95ZiIuVD8yFGekvHc7ETdc5nXDCq9p5tPFeJhKOBnoZVaB+A5HPwLVfkYO
hMadAVk3XlfeN2xKi8yj6xU3PhosM/aQOrdVKywyCeXK5vn1zZdbgMtl891JpG4e
CAlSZXH8CN6c5FCh4CHOmTNM8+V9YGEmYHkEod73rMj7lc61OQKxrMO/r2Ufau+r
fUh2ZGGsqlew9+M+INQHUzwC6J7RdBNwII45+5/jVRnEQ0PtNArWhCrnCxN/h5gA
3xurvxj+krwB36183t0c7NrpjcTroq8rKueo+J0bfdyvyXwmuosg1Q+7aD9rUdSJ
Xd1X06N+iQ7QrLdd2c/dpGRjHHMrJVOTnYfTFPEd8nLLgsy7Hqm6DZJdASRmowFI
0Jx5tyL2riIaKLS17uNYCHHkN85IcW8U+IzDTZrdY1t0zR631EUY4wSxP8J1Zei6
i901hVWI2a/B/QCsAiR9Vu36tpTHZi0xVjLRWDo17r20bXhNOiIvjzXLCkhFalad
yVUyzPE3WRgJcTIeMFoa7Hw+UIWPuH6etx5bwhAmYvAC7CIkPsHL0vfeMa9laDg/
keKNVsqaDW+GqWXPkqPwc9HaWHTImYESEZ/JfrF4DzmKr3zUFFR8PrU/uTEr36g7
2S7LPnbRY4y1BqRBmf6iFnslsh9iLi3zuzX1rOFAnPfQ3LQZSl0jAwHzMCqJhFkv
1jjAfco/iaKhtAyDINWEQW9USWwM6YD2Tb5EP6d1obhLRmL9xNcgSMy6JJ4m84hQ
pBfUXZOrLbx1ihohJ7h84trHwEGLqW2TWpDAMpHV8vIEclfaaMgv24TS6kaZWnUa
PmyY3c1E438K98/gUFrh4W3CdELiXzWFMbSlYX/+I7OmWR/wHk3BaeKSvzLRSdNl
IbmQJm7CG25B2pc7/aeBVqtMJ6dGlSlj1bm/9LjOJo2WtZ8YwTmDFwfbgruLOtXA
fgntCMxhFkqbC02BOW+bA1agzOR7AYXb/BjpvqAzb2Za3AI++nbMJ04e55RJmUqw
WiZOoe9kVwZvkNpsMNNPXPu/Ll5bXPmFucx8tm6vI96SdiHmMiW2XdcNJJMOBdMp
7hukxabofUqkLAS3Vz3vPTaLDC5849OeFwxQWqM7HMdUxvtVkSsgU4X6trgXEo19
RV0LoEcu3CS2hyFGdQHHlB+9gwtHXZcYBHS6UgQ6na/pPm7RAguGRORinWcxH4t0
wicvL08GJeBaFv1Muqva5SmCj1ApF/J5YY9+qE1p9uQb5UBbMYyfTydgDeNvS4Mu
bbF9WlAHQS6SFEN0jeBfLWixXrvKBupRX2wnClVtEkMlkqpzHy7LbLVs408w7Wh5
EiuWQ62bwL7tMVYpLoBL+9lfSnyvgGgNXYEeQUv9wRCkWXhegV0KP8/OX4KDPw5K
IUwOQtaLvG1bL709TArq5xjYocReRRuc7OGyc0OY7LTaUwuU/zcV/mulAVY1nZ/Q
ciaqN7PPtam8CecmfkitGFDjqf7pOB8vzfXf/juRqeU/gaqFiSvVm80FcfWiLN7s
iSLZSiu78cTt5vf9Tj02NFXMY7IMTGRWTFF74XBe5vXuPfOLBPoA66oCSIXkJ06k
6p4UAJ3ZrDlThmThMGQyTL+e7fo5T5+BkoBKD8RLLAiaMOkR/0AJS779HHS8uIqI
avZXjFYo1YifshL5skFpovdQ59vs/36Uq9nlRRH4cf0zVOqX5Vhtnj5GsgPuIndm
n4XmqNm0WZ2c0vdNjvySWjZGaXn594jj1i9dw/rqJZbzx5nwPnq2QEc0necwDtck
M7B2BwNYnQKZZDT7dE1h7xvVCHy+TVmDRL3BUaXogR2ZKaaCxM7EoMtufka2EPUW
c/G5MXkU0GA14JCZyK0CW8KFyifOIiGvI9BdEqyxwpDYHEaxQJQn8xoL1OE+WfVj
F7t6sX/oOWHKpLeALQ9qhbOsP8dXibygB+MLuJI7UWOq9msPRkYEaIsM/fJPrjR5
HcMKWDnU5ZyjndrBCtlhqFxLqctUyOUnvp2z/pyyNAleNufEVjyOiT2VqtXk51cS
pRi8Sm0AE1l+v4brdq6gvdV6DrlZxCt0JEZiJdP+OKOKB12Wq9tQSrxdvP9oj9VB
O+01zVn981Pu43HnzYdLpvhYzH49tdF1hQbo+xZh6bgaw8tMk8fY+o+ErzsDe+yp
xpqax1ZWsA1B62ypVGtbfdJ7Oh4i97qqhFY25Lpb74BHhR8tWrv0ebrmj/ARBf6x
ySaweHAW3voUi4bX0+m4q3jYfho/xU3QBSt5fyNj7XzKAcD1cPa2wdu/zfdUuM/o
mXv8/O+htpbuznYDvsq35cIqlWpWW4U9Hxk4/govKsYcQS2rF04iD7nXVGXniqvw
ztVlEkUmU+LOiLsixtIDCzmEOdwYaILi7e5dP+63gm1hZzqMU+KTH5yTcab6/GHa
pVDvSDUKXdjQ3XcR6cX24gMmM1mh3iTEqM3D2sQQkJjQrmarzCq9+OBXkUOamxW7
WfcX+fB7HVbmF6LVon3QTngA2/D1y5l3pKSdVaFNG5HBkHS7XA2vIDMxLEyOvzwJ
j5mHWuACBbjQI7yV2fYE0dQPDnJN9QULPZO36axlNBGvyzTdpGuSIk6ssvgizqlN
G0wB7iUcpBpxZVnKVXKHGtjO0h4+CH4R2vlygqbav2gHfjg+eLUSvReqi46RF/Xs
DdBtWiA5b/7gP9tzzlqNjjN64eaBXwlYoIAVR+BpoaDHo/JJTs2C00/iO0S5mphL
0q1bU9QcCHGVjAI5PgNUpKr1PwuOi1trYmVZ4PxG3d2Wn3jzay+t99feGuCYJNJM
Xyr0loYXi7aUdwdtwtuzXR2/cbS9iuIyOjuKHjX/Ea3RK3Iq4sq5mN0QMsoOJSuX
i3tOgPN3qo2OGrsxMJIJTIPzJDhQFIAOudf6A2pKSAEWVm1q791NPUDx4TwDDF5U
nnVSqvIEKMUj3tRoLKLZD/bR9QymJxI8SXHS75wcnrb/Jx8nauC5XoS2wrDLaGF4
MYN4CiTLHkcyMqgMsRPK13z+UEzeL5wTG7L0hg/mZj3Tvsr3aNKe7wLZzafpZszH
ZL8DyrTdozcm2cdvUygud8sr8eX4ytBzbIL2jAkEXPVVr9hXP/AxS2+gcj6XLhQ6
/yq7iGsC1bi5rxHQxlEqW7e05wTxgSPplgwuTU4QmZt+jIXVNDYUTvn/L3Fi61Uu
wHkP6CDOC858SIWWtDiEbHIouH2X0DdGaf/ERyXN4ePUAfra34oB805r8MY4djQS
aCdIVCgp+Kt/gCE7O3CHLtQuZo4l9hkcKdu8DP0FIpTrlMRmVmsHe+vG2KKv8qIq
qYLliFV1M5qsl4OsOjv9B17Jwf0Jym9707TJW/7gAwXb2dSYiBXvayyl7fzCDbRr
WOClK0x47tYOnA2jrQx0pRupsXtrtL4aiLWUieIHzo0fAMF9n6OgzFGmy0DeXrqx
jjwIDm6L6jzT9Whq14WDdzjcvnA82zYPkmm+V8y/XVUuVjiFP7+usCTbP3/7dB5q
yhqKCkBhg9kzSCwanxKx1+RLBHa1+X21+KjgedAoyCe2TApuV/CuqwqRi5ZlRds8
dQo2xGkPlyKMAF8elIA6fYDj1+5B8vweJASehmwGri7ZFlq80NtOxQzJscC7sdu9
EcX/s+Q8qyUUDOu8Uf66wrSY/4xQ/IWG7bPU7rTW54aDTsU78s0UhubxDg1OdIrN
l5RoqcJhWO4mFZvAZ7/YAWNvAx5ieOp55KmTdQj00AkxG8OjoxKLIQyYfKhCL+Cj
I1fC0bAX8KN+Nyb2BJLiiX7xXvlyPuy8rAipGSj0GCS5YBM6p30xmXrIjG0ctInr
107SKkOnMyIP/L678VAyDaj241zf9qdbGNp1GhrOmv2GwEx51fvJKDDkFm2N87FH
rXBLdKrI0A0btkPtGQK2/OFiBErsMs2nH0y5EPKLKeOiPWU/+Mz8XTG0kT4Mkzoq
Xtp2nL1zAtluFpXyVVuvniCeBy7rogjO7DaczLVcdoC8SlJl8muFV4Vc8prDnD4+
0sERWjFVvDhUJKJu3+kJx7CPEI5WA8tnbGetGE1zsJywj2t9BJ1y5RbKxbwP5TXz
EHq+odFLqmgFyHnLHtmMEtbp9/5ASyKzqQqrvM5XVFeFLReHSg5mnboAHDDDnUW9
OH9kUUlOlN4ClHzfPBW4m7zvGwcJK1+/h2Efrx1DRajwDsmf8zXNbMNJI2YIDc2z
pJ4l+RcsBZmWfMnY2fgLKpD/T0TK355LByWuJ6HTHzM6MerW4CR6jR34cIWiudD7
ytHRL6A05V5uRuXpXNbg2lciByXerulgr+mvh/wp/O6eXHds31o0vhDmd89Zv87l
/3DFKYRZeD0J0oYJga7KpVHJnprvlVFWY0rOQP3BHFjfmk4AX5x3uUuoxr+ETL6B
12n9vf69ruEd4RXmgX3rImwwAWJ5TJX5jRYkGNcKo/lXPyhR9iV9mdjYsGCxp23W
UFRYev0fpu1/v44lDsthrVlhhPdxow8fTYBTGL6l+oXUqcTLftQrPk1A1CF59luq
6lPAO8/zJg9OX6RQTGED5IqyqYzaDBMg+QHM2yfVjWtNNXd4ZEQIUs/LgHCyrayY
XnILq5c84o+FzRqpSVDikHckhqI9WYx888pe49QWp9y9BuxOijlK1qetzkZVj6nP
emS1i5F2n/wxYYAdt94Vo2v/dsA+IRgzzCNsV9vdpI7phvDBw32TeT1rBcW58XrD
NAewA7xA0IJNJ5xN6Iy7AAXjkIaugZ10ss9OCbl/En9Bwce02HZbHeEEg1W7868r
yGrxxnzJFKeq2JuZgh/1r9NMv8tkkdvE3SRoJprn7ksqi8+2Ve1asOAX6wsXX1FP
wGPzi30WipphVpTf8RYRJA4MB+0lu3trB2JUozh33BR3VP0Ps3uIzfAGJAI6inIC
uTwNzUwQ7RIEtiK4fvG8OOXy4cwA/ir0dNyLs6EeLqYGSCJhI0IlAlL1gc3ArBpb
y+XWrU4haehCfFwkP/L/8kmGIzRaALQ6dysknaYPliCPjOwGiEneXMcchI2+gkKQ
4s/PlimAXW3Osn+vFxCdJz8U5ZmkjYzOxV8yf3DIzYQMomxeUFhDfEkXcsFo1TIG
wTOiCaqP2pDqwyNj5pzWwczkrbTcMmo1SncD5snFc/BP4SJsKac9OFw4CqdosGW5
6uL9cngjewyy3MuEBaK4jXRPudlAfn5UuBTY3Gfarg6PSQ6ukvnmw8oWHdoMmsoB
8ze4SUVaDTXr13l5TFjgsY0+xL2aA+Yp+L2a2VHuA7FyvUwrYjbJ6VooG7jV/wo9
YjjObJiKnLgzvEnmnvvID5+iUllUPDf2+ddyRyYv+25sUeXePixOYke7zrlhyIxb
PNoUKOXXJ7MDBS0+H4FP21EoUM7P28NMdzzPMSaqtFzRdwIXs2/x9AUMIWRAsLNB
nNeC0h+vaiSnxXFiz6kisnhXf4pe9v9FIIi9M7I1OpMh3oW6EbdnrigmdGXgVqI1
Y8fVmCPL5EYCXM9hYNrcxrAd2YSU05A3u6z67a6jCaG7OBDPsnxFR2dvDcX8euQW
Fg93LGZqnYmbZ+66HqbbY9Qw/wWjhkxRQRyWV5lExm9i4RGcVuqN8V2FIQewqGWV
bPHaQP3+jZt22pVaPoma5Wxi5yjvX9ZdH5lvyghklqccrgIQ2e4K1y7uHdBi8Q/k
bmY22PUL7q6KPiMdR7lekcbO2NClyRzgtgRnAxBV2EsdRKnH/C1y22VMyMMstD4R
DOMtvIwmTd71L9B1wynkEfNxHvxSQNvgdqAd/LepEMgPv+jmTyMyk06/9OZHn7+T
Ox5FugVLKogNb3dE48ZLJW7OVcK8DhEK1ATnRcorEio6WaCviXpP60pxVLmlfK1B
Iknmb2jI1yJm5J2LKBASmUvPy/6TkmbMpgPJVS2v5SUSez0rAXIZyxmMM62Fx9Vh
+9HyhQpohJjwbBKxF9ObwEwOQ/2hpIqKgC4JFv5V90agIROmONzeAH/spUPQghDh
/0bHyI2GlYhfebhKWSNhetzImv9c6lLGrsVzCH94mRmaLlXyfJbBW/3D2u8Vl8GB
xh3mqsOgmQeazkhhjms0Ea0LVbmw38OvvbKB7+Ily//4B0oYCrvfDUfBIW6JJ89U
QRTDS4IEydiNxTyZ24l5pJyUcI9A+5DnR6jYjJN/s4UtpwBvjfhTCioSS8fsB04i
tIJQq5DRXGh3B2Ciz8Uf+lHjayVnXcgYLqk/x8iCQnyGw2ddSKo0ipZxKg8f4HX+
6C64Ny1t/Op9oGNVU5VLzNRDmRVExx3Rka9tq9nDUC3HAUSSNGorZhifEr69nWiF
byoW1TnY4bL3zFeYH1DyXm5ahElCoWfek2RApk7X/jF6xHQ3gYiJidmynUh9rtb+
KhkA+QqDsgd31nCWvEIdiAi9K5sYb2WI4qCNoebQ533zdRIyZSt8YLEU8fKiAJUY
44OCGuj+ddtVLRT0T0SuKWpxY0IDDTVoGGHU/wAUirNRItL3gwWUnOj2IrEHeBaK
SCNCqy6q14RgfEqBJnSsDvaQcMtq+9w46O/YMACdtclRvr7BCL2f2ACyzFjtpTVG
PQWeEXfstOGKlXrbhJHMMkPyRZvLhqcSXf96oWnCN1F4kYs/EnxKO37L5regjvzc
OpaCc0dbNVpa2t3UP6JHE0eiax80HgdVM/fWq+EOCZfQ7PY96GdLjR4/kGswX0w8
AZTbgn3XrH5mg1jqOjFyE32+Gb9egJtW7wdwqnZK8uZRDbMke3tuH7U5GRt1xgfe
tam4b9h9aeLGQGTcCfc8VLE3FTOtx+Ovpqd19sL5TzS8eMCTvbqQP72ifSzfX6lf
WbNJaueroOKAasNb1g08YgmMwMfg6bp7qFAsz14jLyh5gHXnpublxyYjWt8dUKlq
K+pFQbnaVWAcMNkoaDXMH+8Tms01YA978EMTZLkbMlM5CHZiVaeZ88tDO1+NhuJP
7iYALizVdpY+H7HGAfbJfOfDCgffJnz+SJIfRrLeunE7DOCzK5djHMHnO4xFnnLS
jijjhlDKQGDDw5fGpxYMyq86cpQW03YVLxZwB1IJjpdgGU9akvXsxBlSuyk71JpH
c4WdJqwl3N2W+xpP464343gabJX4rR2ulPcTgA5Q75shJC2CWEfGSQxnhmoEAd9r
5R+G6x3rRv6x8CCgzof6QiUocpuMBE2HVSPoy4bsY9LwPcRov31d0PjGZ/7HCxN4
2nBj1vtm7dsIJgXrAn9YUNlKE+8HHTd2Yams+IvvZ7+hnCxOijyt4ePWhDTX/Mj4
XTE3ClUdff/hjcH8SfDl2WUpRYUS1zkUBs93y5TI59R3wrlZFFBn9G2UgrXn+9VW
y7H6E3mhf+rUyMB3HPSToCliwnjLKVqlZDZWNioyjWlYx/UZasIARsOTOo/BNg/4
GicQFrNYohUgkoVDxCpWEKrmCcDbSAFRmyzvikHtt9N3R8RYrP66pYGJNTtgUwMr
vrJjrOqgX9bpmniH607ZTrwnJWdOVYTjkzrcVJVvW+zgN3x5+GqqwZEaEIes0pXQ
vguyy/FSTejWRcYzyyyitkSMAukFKr1KsclC9fzfAa8AMxPrPTxMBhTTQBuzOGIQ
+EcINMO1AvkCK45O5idw78IX+KQ0a6uy33wuR+z1VyxkjixVXK8w3YNKwzRfF86I
IqZCo1zKY/DB86p5QaUUBbmvxLlAiylU4aIGhow4xuWvJ48vfiLvjRKVAv+a/HwL
sk8v7yylP13QV9zsR2zoJGY6rSHTvyfM/eyTz0WMb3/7dC59tC7Kv4LfHhFHsf+9
YI7MJm7PXupRlB9xZKgeHkZ4AhlVgxt2H9rF/dA9+kQ3Ep5eXTTX8bMiGID+SQ1R
NhcMSa2sIUoZ9s8JmiXEoNEv33R32IO4ZFAv3/vV2K0Lk86vYFja/yieywGPyDav
QfRDpy+ACMBlypoDI0FM+gjPwFdfm2UZZd/bXwFArMoJ4cqTm8fB1jnpnW1phxeN
/YD0ASKOz9Z0XcWYNJvtpOZU8VL4KDLD5AByFwYuZLYg/J5g72WO1wnoxNudlMpE
fQqM9k+k7nBIAC+m525rW3yjGpgwBh7qYyGnwz+/Z4t18N8u5uzI0zBFsg0+TGmg
C69dHrgAE8xbrF4NEV8LS15SJcsr1C4zBrvtALIBap/FIPGDpWoTHFjrfoHwXN/T
/wrY7Yo+QlaXXxMUzUmJgFcBGkjdJEtTUPasGOzIEKDjDWOZRe4QdkYJblA+Q6rM
Ti7UUIqiO872ARc0zz5/xrX4Bj801HaU9WVdJucERWiTlrLaDpC1xzBdPmWAg4oV
FaEshd3EwKvq7YYOjQArmldQ28H4bIldQPB78kGwaFGtER4GaaNS8mLQZjw4RomT
kqy9xuj6oIlq95VVCjXmJDgjxjpfXbUjMzBhhvmwXkPY0A0uAHRfQw6l7Sb7uok7
DKMgZuDdtGJihHh83HZbOQK07QL/1qvuPOe1a8iR7XjoSljqb4Z5NLb0kkYoyme3
kU2O4Bw+7MmyPymrNqIw/A442TAorkYubiEkm0qNka5sKauMbAHXgJtABSyMW+vj
miG/2N617sF++d1aNPAtMj+lkNGFd63iDoq5ixOV4cf+0jNNt9yXVuCyTZS/+/Iu
x4USHadhtlCXAkifAPIdJGN7+vih9QZz/EIaBDaPNDP9FYFwETKllhZBwYGHFMS8
J0bPjVWhAEIIDVTM2znqDQrJpMj4V7aLH+NUs6gnph56O9esD441Uu915lpGQopk
EFY06bzeReWGosmWKl68WWtcBzcEkBChBoojmzBj+t45K2OwuTg/JIPK8C0K+FVm
+761/AmpZ1w/p1uqP2KOH27YEw4B2S4kAhDFcyIYkF8Bqwr67t+vFdjE52I7lB3c
r3EcST4agmKdym1vIiFXrb6QS6Fm5P3/qp+8dUxbtOUxV2Hoaqc/ngTjvVTfGa+5
hDxNwInYLdqnPemWYpQ6cJN5e7G6JrMQeHDWgqbYUbQdfKnadpn+PN+TkVFta4Ct
aBaa690oIIWH9xXIxrn5S2QogaAJRXESITcuzRHG+NZPNUXxTowvDx2QmAFszYaQ
Ipxoj3OiIyzon65EDZOIjZjjk6bWNhEHjiTQ9z3EA4HxjLrSh/em8MZmjo2C3Zip
MN2Iuf9kWXRHJgbj4LDZ1dboJAp0RGQ/s1UGiCcY3dQfYAOqojS+rk4TdD+w8uHH
qiYxk4XnZgnA043CD5UXAMD0/DeFdRWI8IG2LcFfith0eVgBvJGobSGO6nPmUi7z
e+IhjaOYBiDhrASLkni2BbbvRFM6H29+Du3rdD3lCRL3VO8yAUSqMJUlC1V4xAwa
oKGYFF9I+Ht9CC4DH7gFd3lBT1EvdRmLzJsMtfFb+xb0TzCz/CYOH29bM0if9qnM
TcoLhGQ7Po/bMfy9hqwE7I4d42toatR/Cb4VnoBsKq1vNyJHhMyCFZjnK9wGU879
lLyFpGvFxtDDPgKxv9P6Kn04j5pkcwbDZIo/X1Tr9rCjvLy9ssNrL2jvJX3J1dEG
hGhkuyL9KUBGrZvktDXNdbs/0uOT2QX1J10zvYLGIxjf60yrduU62bpQt7H+uAFy
14RxSMoxwFg++RHlBtlCPdqOUrP5Y7TRdbZ3rKIf55sT5XIFOx2NXpcJSY14OUFR
6p3gRvYK0l/iO3hEd+9DyIHgige1AwX4kX2u1W7QOmxiiByUUSf9A76ufRcYhj4p
3vA5VAR8+x7Oa46F2oqjqP6KyWDLUn0/e9IZqwslfgs/rqhsTMPixS0DTQ2pw84p
Sbr/aoHKaGyNjcxdSb5UjxB88wJLlSgbOuzjmwp8LYbdY+o7nLlVtqJNXKU7c63I
rn2qW1sL4C1g0T6qEe+xCU76rsee0orLG/JiVX4wpQXlgqN4Uj6RMXebhLZK5nmA
8FfWa1lO3EGRJVrP1sIrfGA0RSQTfUKADrtpyP1PjmdZP2mt1ZZTuEB5z0K4OpXz
wa55/1lYe/eXO+eACZwXfczm7BFmB5kxoigi24+Fbo/M/vvAxC2SXPQB2OODXpS8
2eNtnLCmJ7aZM1Nnl1ASe1i983Uk+DXLx9eB2OZaaUoRM/7ZWa/mfO1Ui9U4WcIM
DMJYcW/oUoQ9yqr4zUgO3Dxl0ivO+4+7NRpxa7Ro7cx+dBXgPuV4Lv6g1vTyFLab
psTBp0Iy3Jjg03aAxbrZc8Sfw9EaGMP/GKfiARiVlEumFWxYqxWucR6YbAEJWkop
Sxc0CSmljJf/nuqsccEgSI/epNqke8WwYTlkaBnYl9mJuqETIUZ3MeEOHpYEqmYe
iXduP3jKwf/fSgS2HpoSzFRS2h3AWINMVg9mjIoURNycxg1dxrTpnpSnaodUexQD
i7/5+hwz54ZmHIfbzxVpn9RIRNnXiN1wT2INBSKxZQz0ExlAAXgxB5SER+ffhIgU
jXObsVNScEOGi5DbYXxeCczEsASul2lcOufN8HQBseJTyGJ0TkdJhAQw8NPYsFsu
A5E1m4UDa3XQ9FtSTh4SJFupz6ozz6Hp1u9LbqjYdNUFfQ4t8gN/5Tror3iM0OX+
vNDV1heMndcJJaiDTYlTNa+km+jvYrSpotQqwfmPNjvAjvaMDBJSOxutovwTRxTA
rnLgLw1NA6NSpLwBS1CjgVYHo3MVOAtcNYuozn0PxGO2SPBRQG+iS2sPw9fe6H6W
cSPeEfqU+lJlQMbwEsQFrclOKmEf9ub7ecCX6GUsRp8csKD5wdvjoNzKVDvsqvCH
ruYHS5RJq1iji5Kv5LMcaiCxbz2ex10R/LyELntKVv8AfwbaCPhkT12J7DTgu46l
lHGne9MT1xyn/uS0LM5bqEzyV31rfgX7GuzUPvOWFkySaYmph4F+itiTWCnOMQu8
a42xEfYnmIQqeM9L7MLuz2P8RmX21XTwrMfiHpJjYguPT7/vvJAcaIN1ykbw4Ze0
VEblABthaXKr/jqP7nQqoAs0QVEwlm9zPME9obI2VUUxW4fKncqa0MQ5w4y5mwMg
bIVXup4bnN3829+MSvW6IlLb9On+zjMZ9jTdLLn/869EREmYVN8cX3ygOpmeBIA7
aIuRG4UJM+ajAoPmSgV0u7f0+0U29ezxJwMUSx5dZdoGHo7uGa4yURR9q8ICGbbE
/G6GgHN/ART9xPJc7oip2gpIPgAAT8uMXwlSHvEXIPMnHvPGZr9CzNB3ZFezijYs
4ULqQxvzFcskDr6T5zc6JUzySTH6s8gqPngE+jQtk53tWoJAKwpi10bFnzcbUbeU
cE8zDN4Pck6xTJQ4Q3Ncad8Ns8IT4T+Ntq6rsOWHcNh2H2niUqNPfzBo94E4T1GX
gjHJdKocJt93h+ZBnlKage+dy0Ois//OLkPs7CqvawAWTzOHI3JMRUe2C5iS4gji
I1y4GknZXKlySG4V2rQ4h2+qo6Qt2Y/oyYt1GBxtK+S9NhsPQBycaiQttGqfilTE
ignxtyKbPXE5Yfuzq9VPFylZDXEj2aLoKv61R39SyyufbH7zNLxnAwJMGWxUtU7X
FwLvB43C4nt90NNgoCpoB11fJNFgcBcA3syTgHjjAvy82nvfrESBMR4S6lpPntTr
6/qmzaYai5sw5hcIPEfxsbJ6wogAX5X2EHH/2v+07baErRVWjZG0nMatpTxS9TQJ
vMwaaHcgac7DPSO14NDGbhNjrNMD7VVfa1WKyEd3M9KI7VLYHJ8RqZUpTQ/vaOqr
FreleGpbcEPLP4Eio39XcfRh0ettCN3v9JoWgYL27er7ujoae/1cxHiiMb3UBxUx
kT4hnpqHLFK49glo+Uxa8ttatIk248wNgFEa8hRpK86zGdQWY7XsAO4khgnTNknn
Wz/Lm7f9g456AC+B08ZgS+yiO6DVuXLNScdFNsZffeFQpUwIX2XXW4Ac3Sbp3h0w
nIfJm3KVN+U/Y+rq/4+3SV5VYoPOo4aLsEzSyGdJsN1L+c0TyfIeYWcVdsZnhAew
R0VzAjz/7ng5Hee1/Mdgj6VZCot46srSiTNQV8fOJ/VGAItVpFM+O7241WrGCla4
RcEz9lnQxPArcN2NXn2S/zR9Tf4xW2CQb9HsUzNL90Z5/4EG0Qqk1441Rd3tdflI
SiVKyiSPCRphimewhenoO5Y4GxHyz+VGRbOiScW98ZU8BeemWdhqjo0fdJxtUHiH
vKHhR3bnm882kRQ+h/zjuCqYNAPZBZQlPTozxeA6X+g+B7G3BcMVIJpoQTTl/7l5
DY3NZbyrRssQNci037z4xjZc2tqBILVfT9uAO5+hw9AyZgvFVQcW/s7U6p7wlH5E
J8Wh/n41/R5NZqBavhAx16ilA0PmzAeXyXNjCJP0NNSKoVtJlJCW2XZsQUDaJw3g
sZ8fIMr5U1bRxgmBppUPUXalY5bzOQjThitZrjGWDXRKrrocYqZuSgFotgDRFHUg
5X5g42HurnatFT+jlq/N25NfmEvClAKKyRk62QJ/pMbEPWJTfAIm/w5h6boRRfCC
lO0WmiBtUZ3+8nE6FTwOFvte4xKVotgisvW/2YxKEBzsONEziRc0QKo7EqtE7C28
VEScc3Wbjs8nVnlXKvPS+27oKWcpYjhfVveFAupH8iG0kIvp5QKdZ5v/hO2Jv9fh
B/AHmbm1gVrY+mUwNCTkmm360OQoWDSRP2U+VRrd+lA2VYSUkjubCmtylsto5hGd
gfP1w1qbKCPNTQhxBxKRhcgrpozIhawQ6LLd4QuhooOMpyGPKBGPoiL1szHF5V9u
Ax/XxcMmzSorgsv2KL92NKQ+TcItnk6xkqZCQ8MWCkO0VbOVY2HyugYJeYTTpzxv
yJovFUgFJUEgJ2UMskHsCb0ReYHptR6jfZzANQLN35v9vrPEQ8fVthOSnjkQtkx0
j4zx4nrOA1UVZFqOy3L1yNgdEmGhbXW41+8qzj1YCCyWg/J11wexaRf2XZhNcO5B
MOiEeDN9CNoseWzFNlECh+Wcf8XmV2bNzyENTc6CROfOpTuTihshfEMQ7OcQhxie
DZGBs4aofvhT2amjyTW/pAhfQMrzd9gMKo3gvm/hZzj0z/REQZz3FiLjATi+eoAl
C0HLxHSha26jPhwlMQCojFvymo5IIoGUh0iPzgcDD0daywojRtTJrd4dBi98noW9
+YGEOvZiO6IVMYHZsgs2AfbyjabE728T9dHwFwBLj1Z90/ilkhgnVabffFXxDEUe
6z3YTnrbY5terJaJRFTmlUH3wdLgv1wmaVsm5/Gsv94EmCxs98tc/hXDKVMDHsFl
um67jiOi6rzNV27x81z43BGFSnRtyoIQpYh0cdoSP7jy4yKHU4ZulNOPrYOdvuQ2
cDiKNxdlU3P4EmBZBxmrn1TMWkFTHrihdFC0Sf0yjvz/8Fq34AeW3lHZslsfR+5i
sela+dqDSQCHZ5Gf9QSBDIU3Lau6QxDdC3a4sfu9HApwJGJ1cmRG/T5mCwlqQqM5
RlgkNPST0+03Mk2ux60R4P956dQ/caCTi5Tc+df1WnRqBe0kUZU8L8SwbiVwaEFK
3+6ehBm2zAeTiPeqHtRpC+9NdQAy3u2EPkB6qqaXKakluuKpQQo55x6/wnMigD7Y
AZoDSYNnPrZstrZV5nSNtwqeTpWEc7yM3l4GEwaI0jy/d75q/6bJvFQK/gCB+PHk
KPJ9DjxP5GKFZLK2Elo1EzxJ/RUjjFQyO+32wRx+ZSi1coN7brsOJ9aPqZkHK2pl
xtxNxbP7wq6dJbwcTFa8wmq5hbn5ZL8KSFlLEuDE1kuVXqjb9aJIg59TWtAsvzqX
DfNESGi/8Yqm5qK3CHVFM1F2uVdUR4FVDzmC8IIs2pZgeSEWA/SGyXdMB3IHb422
+22XIu2BxX0YXRMEztB8bmbK1i2ymI5v9CSqbyEp31fH9t7ENIN7EE+hnOwuqWuc
cfG9Nr3VCqZE2Mi9GuF2tRerTQep32vDCGdj0pg/OPqcFNdKO54whbd2BkCzlcc9
VTzKldT85jA8e8cYpDAicV0DnMM/qnz/1UFcldQz9e0dNHjRU6ej0nkUK6AqLUkl
aTAIlCu+3V/HpMtJzGViwQJY5yQfwMHdDWFs2Lp720kLORJf/c72b1t6mSprzn3B
ZIjgDnBdclbiqySYSyUKRhVL9IoXSsuemthvSuZCWhsqY3o1K0Rua+q9MHBJ88/s
fm/tO/72JlzvWQhDjrlExE47tHgijiWufGF8pDGPwRTfiChvaWG0kmOGXIWyaoGl
sdzgX/vv7KBHRB/6eqhAs3BTSDn37gA1kI4115oRv9dxOLB6Oc5NZT+ArWZWMkWX
QjbwhnjezXRmk2PjIv4B0F5uHKL8PGwPih1GLwM/VETfVgKK+Y9Zpx1sdRwJ0EjK
tpC8TWRH2ZpMOri2+7lvuwhBKsTgoCo6xnhtc7hzyK2ezixiRXbnTyVMyrb+06Zr
p3Dqxg/VOeilZinT55AwOH3oqiE/YRemRtZsbc4ZrTQQCCR6Nxp7LKNTSwa0cCdR
8phxKsAWBj0PpCWNdrR9qjVgRsyyIh98ZZSixCEtWqYSW++BS6CN6VG3v76V+urc
qf2yX0/TXnNJxEgQ+O5hygpkalxEzjsShMbto4QuM8zNxJ2Xdoq0tPi3NQ6bLALk
D5c6Ls0716kYAQdQv+DS7PGYiuHJsK13ddDSslw4EbXz3yAVlSv+6pWh3F14g3Ju
GNXiKa2lae7O3/B3mRnjqHh5yYHjzHgpfM797ih2oSjPKtH4FBD/GCZjWxPODLho
9vKYHlVc3VfU5qJEoV/ElBqmQ7u5j9CdnRNKOe709fesjbdH0qp6BDNZrUtyp+BI
akx7E6WK+yntnytyovjaUWnCTfDO3fkTkkrw6J348Fgw1m7WFaaTN6XKSxzv3Zsj
l1Fk10EfeOu78KQ/Fr5G+5Y7AzvirZJlMmnl6Hj/g/09RI/qvuSg8eE5S5YaOh7+
0KTtejCjcHdGZ2yPoyA+DE4z9fzOf6oBJvVdRJ6OQhPk30XCtrK8d3mXzHRb1+n6
IvHDd+I7ykP5CqlhCDO91tQ3EEO8nZYxks144sje3TffOa48QmgAIlAYew2ckDOc
LEQt1UGbrghX7gNskTlc25TY4/ifkKsBvQeO2TiLpBAxtXbF/rmqC2u1DKosaADJ
8Fz6gz8RnU+2Rb0TINpXJz2h95ESfYYCcqOaUh5aYWGSlCsfSZIiamOHjPaOU5zd
PnjKR0BoVjRzhuk2hk5RU9hCiXIdnF51eInDanquNhGH5MGNqv2I23bxZGS8vNf5
yd6F5w0/xpxhHwyBbGzcdJl21sV9RVa8NoBi49/DL8CvRiJ87QHFREMWNYvZiOt7
REDgtapfkLTRTJH1jKv2qEuBpbA3NrRmTx575KFCl3NdP+Jk8innzt1alfHvXNqO
ia3LPZZR/i+0Iyyeplm6CtJEZ/KAiNgSXokE/NWD9H9pH8+QpWAyOJu+rHDUbzFC
pyPniEiB7Sb0/xjJbl5ToLUtfJxctItvRYwtiWxMlMa7/ZJHt0AJ+uEpfYeWceAa
bf6fPYG7zY//eDM+Etn+RS+/0VtiyqpaCai+TSVev+oTiEL2V7GvL5F4OxxfFFwW
4Wav9IgnCXmLs0hEie4l2/nfvken2zj+xYJWpdOii+Czr8ryvPSafzfplJgPIylS
Qfwo5NaT4tyqN/fLl4XakZkQaINwWBAYAqA3lxQrXiGHLN2zluxrqHkC5SQ9T7pJ
+DboXOKtfXAmRo8owOjSYFxCREJ39iECqxDN3wACvAj6mynIM0FaBCFVAl2edyIJ
FwB2VXPOyK5qkh3m1NRB7QqRItLaeG+13oiNnOuZ5RxMqEft03i+wMOypPUuCVIC
BIsczf37JXfX4ydsAj7lYLwc6xQfqGXuF1VOaL6wdp6qujvQZi6lEBwgp0V2aQpy
LWWG9pCaDAoQ+Ve+iZMiv9begxnT6+KkY2iVvDQkcel4eteKPzWCNgDRNPxtw5VQ
oLoYJl/TFxIndWHPjNvuGiHifBzf6ZecS3kbIRuJqkAND2mbY219L2PUFcapYPBi
0BAVogHqJZYEfo4qclG2O65Um9rzqtVR47XGUKmMYcYr+iPmm6r3Se3UjIhhXv3z
YyMHN7TSgymwtI8IxCGy9ENnn6oMYkD5VkvhKwP4CNRqee2x3QYLk9rC48IKzrVd
GLugUY4nVpE//X4KD/FsfM+dS2YQB9f/eM+cjHvoaLqIuc8pRtI2qpIiOlxcS/5i
m80em4RCDNMlahCig236VXD8z+QkakrEAmGxO66k1ftNAIlBkYQ3LjlgwU6BQF23
cvH6ySwuoCU+bqpGEz43I/NP/3h9ubbVade7Ij3migA63oZvi2AyV+W3ufJWCHNs
iso41/MgOcdkz6SB8nFpazk/sP7Q2S26YsCizIwx1fgRMKVKPuptVOLJrOCswxoT
4kawc9Dg0fNnmyh8IrQLvsosyL5BulOAppxPMOvlpxi8JRjI7w9hy0kefDfwLXy1
az99AWeM3e5ure6Cx++pe7+ovj5Gann/jWjOsyrhwi9hbSeMX5B6+ZfvtBEX1rTZ
kJAPWLvIYq4BcIUTwUzXEDdosFN+0i6MsnslCTFYHxNhBjAMddbgLVGPecEIiWP9
rjyra4PV7O9kXv5I/mrUQKyRhe4vQbtgJicM5EvawP5bNP6sHsOj8jBraoJ9Gz7s
z8Lp+zrnx4PZyh1FPLURNgFByO+QQRX6ZTKmI4BKfYdIkJhE6o6o52TAdUq12Bq9
ej0ViRfmKq7eZz2SOUvwnxywiNr8H25fvkr6sGDinYVQuVzAtDFOW5bFBFl8rxza
vXKrBYk8kd73a6nv9Zozcp2p7PsS5bKpslTIYDiQ+AjShpEbVgDxvX8EqPHhRqi0
GC4XqsNQchbbvUyKF5YKjyKdViR8jXehpyeOgLX2z2bYCbsGkzpYGKuqvwmU/kct
1Z4II7CI5FkhdcoBj9WEI9x73mhiMrDdVDqEzL31YjZxdhmBadmAjPBHoDsAnhtU
3+4xy7I8duBCRwR2etkF2a/RamzaKXYsiGDmnl8iVnWV3G6FVqN1oEi7zAZD3Fbf
bD0ajzpCkfGd5L4+kOj0bQjPKwoj2KMHntx9RAJIL+BGb/TuGVt2L1JAKStD0SuW
3q80nPzaGsIciBlz0KDvyQUTJ5o95dugSaKfGuzwFPad0gyLO6cNaUx1D1cbJf0i
Uvgedo3dwRo/TVvHLCRVesFy6jPWGFfW3rGN/7AMa/fmv4AYaa3wiWACjolSgyb1
ouerM5sFZf5QhbbudiTpTBdSffqof9ZZVMRD9oZw/v+58PobRUKmrWeZBGfme3fD
Ob/BmYbdxSeNddtmiSMX8TwkmESbyNqkK0c5O/JHLmlBZ0t/n/4+z/31eZX1gmSn
OfUqrI98myTQn3qDPzLbqqXKgtdaYzSDAqZklJldYBPsvYjKLNW2grBFTcRXlwwS
sbxxvVGr4J2nYB1uYLILlReXEFpvrbUr9J11WFh17hW9Q9jWsBjlXkaNOTDd5dt/
G7I6Jow5jz8OnREewbjFjjANp9u8YxdQpihpYUt5x2EiOj8V9dbdmnGvFiPhBdeK
WpQ1q3Hx7mVsQQqp89YthAo2FwWnm2vpnaDG4FX4Lve85YliAgldvazkZwc8l3/x
ATvYEVE4MWFWZrGo+ApQj+N+NKi9ZjxV37TJsBMvVusKdR3XLU1t74MbYWGT/4mf
TeZjOUxcQcxmyZkq6DHT64L0niBQBkpYXkrbPyJZQLEQgcxhVTGmgsZd+VcVa5sj
HlIVQ01Si0YwDTWr35ivxLEfnLIw5alW6LVDyv3QZ/G8W7IU9Es/PzoKw4MaVzAu
cqUPV3OruLlMdioAe4Yiuqp6u+bFtKvRN4FlHYzojFtizpDWPKSVQLIEzya5mGox
2cAzEEud5hd9rAJZe/KkEdiSEb1N4W6tPU/WUokRhJStWrkr1llX5nYpYkn9S+Z6
cBRa55sFqrRp57HlHAzPKPDzLgdeYfs/An53UWspjTFwRQm/YAsGtCyH6smMEP8n
F29tEzeQn9Yoc97dciX3QLUOl6KYMiwprm1eE7MIbFP6CXr/FenZvDmX+FoQqMHW
jUiHXmr0VHIfBuhiiMtr5QG8+BrnZ16muKDsZj9YOkfQNJ/lJE8gDPDar0ciI9f5
3PZ5zQ9zfozPcB0l+mQsssrMT9cNKWNUcS/EjOpIRf6LnIdiXuhoBGDoaM9+XoDt
AbQwMZTRllLWwqbI/U3DNb+kYNqaGXo4unwSuwxVTnKx5XJXn3EGaHSCM5UfD7Qd
40anHST67Zvx5D22ceeGAg4/OVSDYxSZVd6/MJBhRrvWIF6gOthHCLJF0871G/Kb
lg9BoGdOfwtyKsrDlxixh5LKRRHRV72GovY6eR/pV2jd+QFVJJyVisGaRhuNO7Sl
P+ZQkKZvqMkHtzYv9YITAZ0TZbbQja9g08jyDCiCEJE1zLaoVFXh15PNWN6GMYwk
NM4M+iDFseuxAlmWqnZx4Yc2qqAuIykcStd4wYeXJwZTwgp50gphormFn/02kD43
5ExmL2xUbqMMAyOS+bMVy5/CmZR8/6CiOKoJjghsR6tyx1ebOQSzRWFFbDSv65hf
RitQ+7Yk/4khPxfi6NRQN7+FfBg7mHxuZ1KYqSaUOTXc7mVSMCw/0wKjdiG+9o2L
d6vQLVBjY0GcDun0imkLo4uXpXr2L0ueEUb71IGPsynY1M54kp00RZ8QX1uK01gz
qlZTZKSvmZe00xz1GkSOBZRCbeUpPdLrVum/mMJhiSOXO0rh6KF6Lm/vNJ3fffvE
kyGAhe5FlUgDDyogRKL/s01k9vge9hXYwQwuXojHHCFXjaLirqp03sbZPIOFifZD
wvSJ6l0XxFNb15r8+hUbnUQAxxtpFxEUiqXEusmj2TPBHV1SorpiZnc/P2Xf+LyL
uqwlLbcCZlZEhTDKofIbS/RxZTC6fInF8MFn9CIIKlTZLmyL/lRBS1SYN+sgGMC3
fFLtiDBGP7muUyIICst7SCKCUhVtUp0qfIyx3MtntFHUIYz1hCphriWsemHfEf8I
SGacJMEWDWvvlK5ZhHfBxpaLi8kaw+XsRmaw54sk+GUIWwaj5Gkn0XgIssVn+pI0
w7zG/A/HJvuUGtuSnbYjEomxC4WLK43wBs53wYfQ1hIzbyeE6Ygx70LfUT10Izem
29x3dS5Y6L/jOXV6Wr+y8zzQYlQcCStFl7XQVELGsySAKbsehQF8nllHtBDSHHT+
uXfyvW8JsSXPDDDVc1Cp+I/lAPKOzHGWrgpNbdn+QPXZ9+v+vQtTAjfD6+R5q/24
dwJeF11kACqKp9XkqO2yufE94UNLyJXw0cfXKhdhnc+rXXjf4ii4uJtoIHHGC6Z6
sCsSKBkf/qeM/7w0uD7EbmeQPlnb3kZJ0MBNpruZOKSpjUlmbCu+QiynQNHMjSPq
/LzBNrRlmR7fEIC2tlgLOgg6jjZFX7cDNByuXmBXebTSmzw0hB/OYuyR/zJdlK7j
nEZOqMTEfXwCVuz2wZq06DDRVl2ZTB7y5TKnrleCk2yMbHVZE9In2YRsI2T7+Gl5
gfVtKKViQfrQtmvhfNj6Wx5XqNrFE28s8xKF6APib5beMFAs/vsnUh78eYP1xAzb
akY0DUNPiFHJ7hHdeMilfeWx4d9OgQ3CLD7vWE7mx7yvaNFdxUpFOj5f01zj9yXx
Mnzt3FWsihRVovuLt0rQbd0HYgRI0NRe4Rn54uUAQYNtru6K4BXD1N9ZsR7ImaxX
H8m4QIHW+/gbWuQHGKguVb+50+zuWJUgON9jwkJGv8RVpPfIJxXh868apGKn7k0c
T11fOe2kkzn3CjzMnuXnclTxbSDuqb2N4Perjq2mpGw6DdrtRkv8sKOzsesGGDrB
lX/xTnR5dDwGTN6hMbk9WE0t1h/yQohbe43TktTLHGggv+p/9GCS65qr1XTD/rwU
XzBBRYvlWaAh/w49utf92vpF3iBlYQqTtL1lOu0XgMLHDse4fxLIrYwKxV3MlLbr
942N/Y2aBSWtbclq3fYAuJ8CjdyBIaY/PqnLJJz4QtJkhjfQSwe7ocOboWwf1Sxv
jTsaFW2eS4+U8GlZyvTSs5pxonjQNXBp13q4iHvlz5x3wbdgDFxySZEjFc9jUpdY
MLOCRRFcaiDCyjq/pMjgjFrPt7A3NrFJLTerkWM7VhWhJTE6r0yt5RA3Ph/Mzq1C
Ez4sTWrCEHKCHszlx8FOqo1MD6dbVu6xk0JzgfwIBwCDd7cJedxDtogSmxmQ26rK
b6shK/N8Qezlv4FlgJv3gJShLsUGo4CYPY6+2EjypWqIesKggvdfxovNHrNWqWSa
r6Tb0eJ+ZCF9satkQbvd1j4QUh02KnLk39BbLJZcyLWFmSffyqSCEhTb0dxQmBE7
P0CoiNUxZe07+cI3q7vJabRTNTb6CQA+xg36fiPmSCGLqHbcLerkTin1zw351Pa3
znPRbeGo8KTPAYKNI0Mru7bSif0jil24LjsXDfJ1tPWdgFu3KMPigsI/qStpCMzs
0OK8PBQVgY0mGQZLRaSw9yxIZ1eMNLnF4p4EEp7laHpScJT2d9BawGADbdswg6Qm
D7qqhF0ScGDYHyf2E6IF4o+MrmK+2oY8LS4QXSbe8uz/uAIIVcse6VrP+kHDZdLR
fEn+xrjZzpywCwL07+AWRjnXv05oA4TDYEpFDUjuXqrQEL9/2xDOGI3U6nylx5Kc
7eSxT1BD245QWZLOLasFNlfS3NkSTxnKJOHVAxLt/Cn6nb5s4+/+pJQjhz93iqdr
PYkpS4Fr2hfkB/NeJI6KVzrpH+CKA65WwXTDfB4KZFTB1MH60dJhaDGk4XYSFEIJ
lPDmapkl78Q1Wl6ncBC8Q+kGWiVLI8SHZ5DOqymBLUxqO5lQzujOsIZK1ObgnK3L
qrG6vm+yV7dXeOi73ehfJGHpad5GpqjoLcB/kqSaMDpJiXgmH7eXaGWDnhjGOS6i
hr/41fzkbZVO4jrHwOWH1ApJOnXIK0JPI6YAA0Q6IUh2hD+m2fpTXfHp2LQGFCl0
wrTq9my4C0yxvFs4Zx7NzBD/iX/qLPCG13m+EADwnPtgbDLeNtcYVY6rlr2n4+jL
PpHF6QmMsmA0cT8D1ke+jLeZ3OtR6tPkZpeyHOzO+FRi8Ps9xwLFE0eFqE1IXbQ/
S13EQBh1sCA+7mOmn9k58kxCWEsy2onX99Oj9VZQexmRTvdZQX/9loI1mpNnZCcB
3NUm4FL8O8LBjXLJ4SC6v+k127m0c8eNdfplI9wkdrxlJMkpGyscQofI9JMTxGx8
vibvou4NxWxakTEdWXfffCMcGiDpMeUH0nlTJZF9HiLzUu4itMcs27uM5jsJq2Vs
CTP0siz+J6Dc3TVTmGY9aIsJP6DQ2ZqcqwuGRX60MWBnSsglulybO1BiDGn7WCmN
MxwxoidBemEazrYufQNNRrAo5pPxs/0AZ7nNplsZIoi0dL/jKZZHJyViJNqWEHjC
1WOD3YYHDYehnembgblneHqfiJEoKuD3sPQQ2wK5sWmjEQyonUjiLcgDQ7+ivEtS
2gPgMwP+uxhCejIfucz8VCWTcB4qt2PzRkhSZjZMMf+Y5vCmDQU9ZeilqwTBSx72
Bpfaw/SoERvIqwII65/gxzMpRVltkwdvI1CTNoc1u2A2EhNwzrYpYA8qDqa1KdFj
QxMbbRDv2SW7ZOcQBt4dCPQbMXj84q8RtaNGs6G2xvvmpKq710uN2cVZKWcbp1mx
/jbpPeaUl1U8zbXlzOxnNjpjwg7xeky7lxtD5kdvLW3sgGgCPG48W6/CHmysRKkP
lEeJ/yx7/HfaeT5PJRECBJAsisEjQ5ZWFW7DPm8ocHj/JmRSfg7sHUVXF+za+Ayi
CHBYaFqp/pmLFYNvgwcIPQ20/E4ql6gVFvDEpDUrCx0kzdflzUe3zo/RcL52NkUf
FdBTIG8zADQ8VsWgJGiEKV+kMg0n8zX2+C8g0Pw4OqyRfN8N/XI53MY3+4tc4aRE
Kws4Fa/kk9mlYTSfW9FyXuj4O3iwGQxTpXOZ9WlPCO+YHQ71IIFlbusk66M/YWsg
X1S2AvqnbWp/pHGm7dQDuj9L62LzVJ3kZ3A6G4xJpH23aFdGVjjqO4E/MkcO2Jpg
Wfrd8opWK4wKR1b+81Xfe+MUyI9EHCJsZk5B2XTnmJSx+/s9tGGUCOZY0oeX2P6N
xQTnj+Jio52PcWwdYVGCSINWgN76JlH20R6S4D6XSG6rP8pSk2RRgLlgPJlWKEe7
X4fvrnBpRosg12XqWXrGBZ4reimAi0YwH+We8jtjKzS42yLPLMERjHfGMvmE5sRe
fWq9KRQH1r97vED2WnPG/C2TuQ7WkyelUA3HDf0jV5howZHzphVNOlmbyge1UEvS
0NIEj/h2V/3881jppDTQorkSgOGe17qyevFrdYWhbRZVovpvd5oFFeSm/x3K8zrD
LaWZ6Algka+uNP+YU5xPwE6FCL3TZ9hFc1a9U1uymVZoD2gH1za/KeR3NeGw3ZQg
T3Ey5ZHZfwaY3l0zXkfRuSrbhpmypXNFkARL3U0sD30orrqOG199mQMS1gtjurID
5EjheVy80HTyjzUMZ63mbjIxb5DFBBaDr9FGFxwqoa22oOcq5c7OVX4+9GFkynrW
J2j0oYradOLK/prtqzCiSKv5JB5HubwRPKMfglUXFaPWctJlf/c47eDH2S7TjAYL
LbKCeG+SVVQFGgdzv2Dsm3FcbuORib9h1ptbKf8iQXd8x8AzChgAvKSl47adfQZ6
rJLvrOV0AMg1CAZuUyKysJR9tXJX2I8273egq0COMpfQY6Lj5+X4u8df/zAtuS0s
XCLw0ZymTn/ql3A1QrUIc4wVHxjL4v6MuHbhDhpaHJUJzf0eHZT/sbqeqiMQwb6c
1/wKSpPNW71Khk3v1tDSTwCXhgbwJ4VzgPFdNQvQjFi/Z/0dTIA+0hSAQLnBo3R6
1btPjGxhRF/njhA+0kGZ5lMVj7x+h2WI6DrzNq50vL1nPxmUJCkUCQIfu+jxVqm5
TtjqKCLpfNnoMinq1rLVu5ISnW980OASe75llp2tQi16Fjnv1U1QQkIXlPhrxKDJ
DBteUvbfPlCNdVUv3KxusT6G2JyAWP7NarO8qtu5R1KWCFIfVdhq2hE33APQ2tJb
MUKXjYkNLiSGFt6iLACaxm2Op24RNzmXSWiI/asuYQJhfU90yghVGCHqvxM+JnvZ
vA5rb1luZX5wvv8xWxYm9YOxcUfkLXHPWwUCNpZA0J6gCC4cJlyOAvHu0bCpO2Tw
SsBygdHyuz/rZqb5lhqevP+0gM+TIkd1h3eOOGUm4LbBmx/G4Tx+0Y7QL3oCQdnG
9l+tDk3GkCeHJfPemflWgnYOaWYw6vJ6d5Yi/Tzm8exlP4kde+unP6y8vJ7YrDWI
kOl7vQ+Hc/P4t3kma3r+ffLjpWWhb4JPtrgqTMfOn25CGJ/I07tK3867lpWfJ8kZ
o2hMTt3ec5GqDTZq1EIqrXBXMhCVjIVWVnbXu7n73ovVodPw7q5gAn+X9ucZ+bff
VCJXriN6sxmTEEuE/AY6PJhhWc/qKTG5i8jHodbA1ZwW5lwv8MNltrY0aCbdgr3J
Yr1mZ2F+6NrKPzSluhuSKy+JlwVG0GdZ/kJ2k9a19K+MUXUvSH5s1nJv0hH3DaEO
EykfWgo6k/kDB/ehyA+XJsb1f87nVvEv41pl17phnVg/574AduRGTJXLor06fO6K
3HoLibEqWXV4SHKBtEd16kcSqwG1oGyuLqPGwbToiRcmHzBkP/F/bh2Di7KO9doo
AphYPNkQJNaY3aZTninZ89rURMk4IP1Y7ynhyZpjgsWtaxXT5uI2FHpK0jETBtCy
wz2Pf+j1EvF5Lbj7Pw2WwyNxZ77fuqWFp9zglg2glZokbMMh7j3etvFR2HeavixD
5H/grxie13CE4rG8ujSZOEXtM4OVgFs91v0u1Lu1cAePLbMVy8riQNHLzGUkD9+Q
txCMQoYtKgIjqUUN9kJga2D7T8CaJtMrfaFcZABBRJWTbcVceVMODhsYUWZrpAox
RKOSX71KJWkZt0TEpj5+WJHgn273WqVyT0PNIU7ci2h2TNEjP+V6L6XLcyEiI4Gl
NACByCtgf8xlmQT88rFWTMml6NK8oHLV0UsUuxlTUZCpekrzQ0xEqbRAmtk57rUU
Wl9kY51IP+kelp8ZLo2awzjeOorpi4rnQH+N6UF1oBJDX8aySql4heShBOYag54a
hD6pS4WoluZgsc/KCIF6BIiX2c6sZgvhKGbkgsVbkItmijbUhIiTjK2vqGhpvOCh
XtH94So07FFsivegZm3aO/3syp68Gi+m7sSd/1XSiGgLWErPSTbgM/B1/ihueqfn
u/0dnHE7JDq4CmGU/rmzgsR8n+C1uheyO2YTmnNmoE1d/TE8Bi2YDkcfciHb41Wr
d/IHkNfUEMr5fd61tVd6wOn/p7Dp914vg0vP2ismwoBbmIIlRtFhr/znJf+u70T1
MI5vKA2bVtsPJ5DkXJu1vUImNF8lkVHECzndA26HxecX3FbqUQZLKzErDb7JhvYH
mdyIpsHLs2vis0Afylahw0xgs8ihhJNs6hvipGMSqqmPDs8oTBiCaxLGgTKyjKvu
/e3HXhfI5MtwlJfj9c1VCIgGWkNfgQcoMtnpSP6rrQ4jA9bcpjxw0PbVmZklgZX+
d3unArEJ3yjasw7gmrNmutbCqAeiZPpv7NvMJ4LerL6RD12dL3XMVDICrrm8jYRJ
8TDGTpFt7OmFmDbU/LH849fJHhm42fSfNe7XYWbGFHir7AFirITUoulnpJWBMCro
4DHy9gIYHRgIO7rB7iZfTP7ywkBCNg3NSguIF7YodiKxL+Ya4iur49IFiXtEIhyE
jBPFdstmQ/W3V+ucFRJJjZXvgizdr0K8wC1qgkxqN2tXJnqzy6oLUu8popR2/Fuh
CI7i51Pm852VbB4zXruYNIz5KcL8Zuyd6oseyaulSsO0BEetyjgkimN4FPhMJQHD
AVvJTl6Oy3qMqt6hnUWWTgs/z4AlY5nETcu0NhdLHgy0qFtB1IcWcmz6/z/qQSni
WqYq5GgZQAnfRQ3po0QHEIA4uJBX2md2A5PvxF/4Zx7OZN/+KWqq4j7GYVGqX1pa
Mr/ivPVEFkyXFeQxXJ0+fyehI3R48ZDMEiAFi9BFwNF3/dsmoRSrgyiyYHSTCj5b
RSdL3YQegCKWouevC5tmmRHkcvR4dSX+ugNuGt1r1piYY0sjfaJHJHVBYLUw4tC6
BOIQXBMmWBq9UBmzTjjEey/nSBNg31QRY6zchL1GGiRrBInIXXnkpNLsZfl1DudA
F1evzqxWp2QHE0WpG80XUduoUf+HWMfb/LNxc375GeURw46oMmuWI70xlrZGSkbT
QY74KMX1/PXUQqpNJMgta3GKb1lO23fpIaujCu8heaKSSGekzPMkvg0Q0Nl9xr7B
tXVwd0xCdqfZFDZjmCvv5YVy9JPGeul7xHdtLWAo6PSSSWDmLR+RCYmpV3tPp90Y
b3JbdHhAOsB1PhTirJXdXBWtUvmvouHVAbvGDnUupkf6mQ2x5lM3iuKyMwpqCD22
x7tB5ylnvGxdgrAVu+73xMB9NPfK799UdjPJKmoWTp+bUB3Tx8nn5wt15gDI9PoK
Mkb+OxYazSLfE5rpWDTW1SxS/+q5jIvfb3y0sAL4F+GzfQ/A4cTbjFopYxFL3XLM
tfUTyDx3i6VjYip/3Fmk5AaFnp711orRROVzCVjzMUpiGqRlo4uk07Kqp/gzvAlS
SvEc3B/uHGnS+Judk47yLc1LvnA+h/WYf0wYYw6b/ScVGHj5YIZHchJw5emSkJw+
bvsnPAn7CVrJZZ3GUNey3gUv86g1YLedAtHTHO95jMWXKGpyFCd2l9O7yeZJ2HkU
h15229bIjM1HejvHd1X2T2ZK3+gRqQgiNvyEEZ6MCh5nTgi8ybFB7QwRSjnQxbpV
9xB8pwuMV8NJu1Gcy7sFYZeomt6RJrdp19460aAxvv+AiZKENVUB4wEODzU/fm1k
dAc2iC1I0gzZwXO7dJJOUuekCiPLX7ifQ5ycdwiQU1FUR/fI4DYe8O/vhNac1HkX
fLpR6TtI3IIW7PD9RxwbLRGSw9uHgAiuO319A1uaDsYtHCDnDLmfi8K2HaLJQ6eM
vl0b97OkbE89uA9rBOP/U0jfb2BZTmn6C4y6lzymw3WdWrOMnFAlfStOjV26ARIw
8b+CcQh1qK4YpzX7Cp2HHY8eX2BrljtBiNWxvFOgeVsv4P1j1IIX1Gwq/+t59Myc
bSe9n1zjBaUl2HVCsOIAhJ+R1IhoGtZ0ZIzf8KMdEtVGExWA/zKqXdvf8SRtVLxa
iRP0Q3FJRYsuPP7AZhpqWpgi/hdp36JJ0EpuiXdyy2K33xnqWCfN30MnNJYz2SdF
SCbvIUlvlYvidpFYos+QNeTSRLH7kFEXMqhncQkD/LFEJhyqEoBdbV2r0CdPOLCs
pHi63te6gtlsZmSAx2LAYBLOqRAkrot+ROXsmnXla21BfuS9+mYluzYu/a7IzqrO
fveGBDYglJMQOinh3WhNzm01P/ZV3nSR4jGnptzEn4d77pk7v1V1nDRyu+9AyVV7
8Ft01xDLLAeuR6j0FLMzIowNgKtr5NhBJhascGUSW46QhzZyc/QfX4pGae1QPKof
1zPl1SYrAcF4LekC9tdPD/NUU3x3xtc207sD89aNgBbkWNf8UaZOjSchYxW3Fw9a
stYb8wlV3iXhIZYSEMfUOSXUNtHd0Lc2gHE1aZUXghuKgfO3QXdN3y4Tz4sHGEfs
nwowRDrKbOwyqC6IagGzVPTRFuX6Y8VSfFwYXBQPrjLP/zb07oiRbyuSF9/8/f40
dsTwMrOZrBGmy+g4oQb/Tg1vXI5nlTx6dYagi6wIhML4RIKx4V+t5ByQrJa0UvV7
spYGkY301cKxXFZP82UrhjSUMAiGff1tOeIUWNn3vMRyCNcgB71e/fiey+SGUjW0
vsJzzju9+Obr8ZSzdedNwhl5n34IiKqo7tZF0W2rruRkBBilI5A5+SxKm1/neUyh
aBoWuvYLm9fvAhf18zcC3ooaRhB7n8qP7Qvjgss7UeGBx3k/ROfZTlDkgr65sf1R
oUQz8mKtANvTHAqg6fKXsYdgsQ/ESnwvFBLnaKiaNcLNUNPumCFY2Ot8mXy0GkQ+
vj783M6/R5IxVVhyJ98Rz22i7UNfzkQFBRNvgsatEs9xMyZBIc8VQ9hIgnRsvYDE
hZgTPTbTMRR1EHfE3uB1YUx/kB3c01MlLxqTvPgQmrZvzRN0bgd6jEVWgacc12ar
iTtIH/V012DK8EJ9g2IZKpyFxP+MhHYL6Sb68GPHZdLe/Ry94G12sjSC125DhhkS
qFvB15E2pBRme0nrCJ1Hef/ixdFJl3POpBQhgfXY2haGGBt//tKRHGy2fdnOhrn5
z4b6W0EFbA3PIkWP1S/Z3MljYrS8xtfl0zTiQUYtcsedqDYwnlTDmto6/lSM2ws8
UNF6ExKG08EnDISRvIvoom/SvEG8CL4A5To3IY5c9SiPD1hG9FhrQYoEhf+Ia4hQ
QbIMQ0V5koA1pZ/9zD0hB5tbs5ks+IMd0oJ/98yxyjDqG/JzQgdHCxEweVfLXF8n
w0ExXkTPvBdfWaDkG3qwR0vQpdrgTtE3IRTSuQqVJ8Fg/GaqStC7xktnXyJZjknu
dRAWTZ7LiiLj5yheLNoGxppCvpoAjnz6etwiNjEL6RL4CVP5niKv2AKeubT7bU7n
EEhP9lNQXtFzHWZ+ToQcU9ZucAylMiHB/iPfjZzdnG/cl/ZMyBUfIF9YszO35rID
kZr5oHxQ7IxKWqUWOlE7fmGnOu2mwSVowiF4drK3LYEJ/Js4xWof+BBwaR9tfRAp
3PDP1o8FioWOs2t4jB5Vpz/RxvkwPy9WJCS5BRz+Lz1IGxA+vJmwpBY34NIn+YoX
2lsOVfEWECDL5p14kF004gt6b0+SvxcrTH66BktG5spjqkwOg/pXSW2mCOsmvaXA
yCoCqBxyEjiucbrDJf1PmKC5dgbSrKAnKxxQMNDTX4gRisuIWnVyc1+TUY9ljmQ3
0PqQjV6MMHty94qEfUok4RSuzBJdzV8tMaWANK29TDtHx8PiIs7m1vLsvm+/+S+G
8gefs/Uf6nLCVtZ5FyTx0QnwWWWxC8oEYAnM5jLbOie1ZJsy2cRCx8/K31rWrjKF
mQdJzUd2fMYfCokFoAk9QhlIcSWD6L7LMQz+FcHGazN23b4cYD8ACnEecI8oXaF5
h4W3zKwdLxGczTyDH8af2Q4xldpKKIwowxqQfdVPibhJLEfSe7wingDuhnXdGlSC
zv8mLD+8xdTLqxTeP1B0f49qfpjmW+5MJPW71AuvRZru8KpBLnbt6uSoB9C9VucK
XzfY6uu/AzZqIZCnHyBy8kZnm1WECmzh5pM/wsKgLv4yW/KJEpCUOMB6fCPF5ZFu
ESo3JPXqb2fPoSIXuivXQl1DjaJWUfNeb1WB6U07DAmr8A+kGwDJp1ZLX76PhFxF
oUVVA7nC6ZIKUqSg4Y2OaqqCKs4Uxt1FoElUdnEzTyem0Wkesug1K345ZBNKOzcm
UBMvwq/Y7ZlzQ+nDf9hUGxily1K8DB4gjZPuEij5h1d0+DPwyVFhvTgI9NX5K1Fz
/TDzK7mkLJb2Pb4Zdw9IuEK1ImxlbZGixoA1gpA/Co3yzekDTI5Bpn8j+EiBx2Iy
9H7jgEUFcXWEh7km1QbUD0eVYHXJqgexLYZC+v253gyyB3B2qhL0co4HKkI8+l26
0TK2v7qRSUzqceVsm9MUZ8v0H9zrzKScdiy2/6/850G+d5NJgM9a84iDCP7f1p+1
+kQXgg3UNIJvAEIQhrmwPQLRvgyvrehHL2OvoN1TH3nayWS4mhkNKYeMZ/VSUYXs
1eHZOyuCgOQUttOYJCeIoeV5HnkJkSNRjdQ+RH28FuT2AQJTvLIUcoDg+LQ2hH6r
+U3jlaiEZKAoTPK4MwQFqmUZXNqXnLSC6oCSieGJeK0gTYUQfE7cPR/cllonsoaC
0s3EZchiVZSGsgEgqHL3PduFwkTfgXybdZPdnsaxQCV7Y2iuG+UqYSDUltw9KNJ8
fgGeLvAzDbCZaN3AtvgOY20qi8rgkvCjdfCgm2EYKQWLYYssntpXsWoqohtHsYnr
b1/G3ode+RoVKw5xNThwSRK3aotb6GduWxS8fA/PPwAtSrFVbHMy6rVElNnzqTuW
WxyFyFbbpFqh2ixY7LVXMcfryaE8djC7LIavgfppOdcakLerMoyIdTlcPUJXgUJu
13F2/fcoEDKtWrNnxcnz9mFxi5FkHTRFegSNCQ+bsSzUWIIBBSWvESPOH2wnJuRX
1kRSftKod825bJ+iMl2DIJUy41vbf5z6UviTcoiuUpVSegnrPEXQCtrQNqowvB7q
BO8I+ijnqD489+dmUq8OSKtMY4X9i49y0Eax4voZ/mvqN6S/UyOmJnpW4lzu+YTo
NOLB+OwWLvkXciKtxFango8P1bEn+sDOIshNovp3zJzpTwkD4cS1jTO9niA+RnFD
86kpgSF8O2ktkzmV4jSjnPVsUPnbtlXaStixyIiZUXUTw5tAIRxU+ly5bPeAEWe2
tt4KTMlZi8M0pw0Q6L7wphuKY/rmiOGnSzcNfHrL4tV2IaSdJSNBaSrw+F9EYR3L
OHANVXJAX2oc6p5LenjzOE50W3FzAGCk13Nz3mmxPTN0zlG0STXGJNFwXK2LF7i1
R0SbL65CWGyZjrbAeDu0gmWO9Z9dHn6ncN/aQbyDr0MbeyhHpnSUdnxh45ctToOJ
KHXT3fYH0wvFrdbGtjKbm86iYBdt2PatzFXiPHJOXiZgUKZVoZaPGCd7Ep0D4zPj
aJO9RMGsAQz4DhbMvgTiduVBiWfGoVqeZ4kJfHghIfU95rdKgBFvOrR+w36+9vP4
OY2zIr+qZ1kcDJpd6TaICyObXQmWf4f+HwXX86FOIoy6u0PXtqP/zHzFq+thjNMX
nbg0sFF3HviKs0edfoc7YR302jOimZOGaEi2Zh+EMip+EYVNcs2gzDcBtbaEM/Rq
Qt02OxtvuzZPQd8l1YBHtm2Wucgtt2NTiT/y4tj+yGSJEj7gTgtr8X/WtQrcAFzN
ziGAHb/gum9cUi2/TGm1gokmaPpa3z6TydcAbsqwM0r7Af3gg2kzz9+1BtZ7F8z+
eJ3jz8le2FKwglaqbhNRDWYBp/f0vuDzhdAohniiTeI5EcM5WxShJs2mcHDCLnfN
9yTKfyGgiHVS/mNzEtJFz9IDqTaVv8ZFkExVRddxlSxB6Am4em7jv6wrK+pMYK9Z
betrgXBo++psafG8zUjEIPT0abw8BUxkd8PegOr3bf/gLZjy2pvNF7wxAh6pmnTv
HFpajrQLfdQj1qhHPrJRtKHl9jNIwfy6TfdEWNslJ1smj/BvPmsbW1QAiIe60hCa
QJKczd1ttRScw11akE5rxsshu4pY+6SnkJqq0BiLPHUppt4itjaAM3dAWACzGtP/
AL09TMpa1ZsiX570DDElFagfBa02YwThUPhHP4sPKLgGC66Z53/BM22n6LDK7GYx
9slEXG1v6rH//1p0IBSLpzCVViefD1W1nmoIKScdL1z6nERvgcEj0VcjNRHzXBio
Etbkg8NU58d30Dyxf2bNuPcw3QVwtmxdGBNpsvNt7E+OhBhAEOpuZ2Tzw6oBnyTj
eghhXLuZbNP6HZE2Cq3UPjg0elxFMYoneWKXQ9i4Z0Ltt3SfmZmRyIRKBeyTWZ53
xPGiQVtQDM4iXOLCr9BK8Jwt3hOJrl8cywVVvinD0mjNY0XS+Kod2nqtJvMVeSq/
wTgNmEZRac9k9m71rM0L/kusFqofJzCVqf8DSw+WcFVrsQxch0/pRO2GUdo63+Z6
Sd8Xz7BY7+cppl4dEXcXiOcmPCpBD3ak/p7uGtittqlJLvhA8pLl/1A9SvRvhi+N
vERhVc8aR/wzN0ytUjVN/gQVf966NBekxgDVS7zcYztI3X6UsrqmHXWWXPLU0Dux
BB4fseAQ6ZDAA7V9GvFsu9kxLtUPzfXOCgwR0PNeCDOpUII40lm9rARTXfaFWOZq
25uq6PcW5HUoPourmDxAAALJPntzCLyhMLXpi6SqSIow2yQyFpI141Agw7IBleEr
/Fi2+ycO18vVrKBBhgs7p0n/uUKgSfjfvQfGSizy3y06KrKu3weKz9e0JA1LlAwV
19+RdpRd0hJV22xbruhzzxmlcMyK8KeWeGGbet68SJydnI9a8UD8xthq3u9xtRvI
2Ey3R107lHITSrFf1j1Oh9XYhegaCwXhu9QhBCzb9GrdFxaXBvAfsei762gXRODl
rDZ9S4JpK7DxNK6lKKExeGNyn5HPufcd47bJr7R/whl/6QVO8VV0x5XBrb67yFIw
OD6yeSWYCMVzDg3/4OnjOy8Y1ZO2U1cu9/YdkQ65IJ6MX+g1IuJkZPUs7ebxB1mR
IPKVvUIgWQWWNmDIdSFDZWLrq7xcQU+1z3X14anLvm/IWMf06clThCvHU8tIKc2n
Ot2FjWc8bWo+2RYF5fTLWzPsrbcr5BoVMKrYIxuHAUA83JyKwbqnqV0em9jRYTEB
V5q0dJuv5mAIRNRDvSWdBzUGJZKrCq8TaCLTqXVaz3QAAFVev/YdzwF1QzagIMNy
ZWK9S6hYAeHP34Y+i8ie/x/Hrr8hnaHlaSjbDMdEQSr5yIIvpV1I5qPk9XYc9XSs
wFc4FqF9P2Ce1AGwCMXhTJGIKMnaqHDUaNnQn2b19oDjyPlWhJoNZppvnhBPydX5
JPZrMVJLF2TYx5TZaQuAi0vFeIwNxuuOXJtUl73uWf7syeAR8to/j5JNkzX5Y17d
GUdHkW6SrEAYjYGWPmUf1BB8BUjnqMRa0JyJDXBBEVmQlHVCXiuE6tFPiV2mk5gn
eFbJK5Y0rvQAibmwV49e9lGkIXHqwtJK+xM748aI7/SWVvGedkjIPDvUN6H0zXqY
q6RcF4+S4EWut3IqMgfLehtUDWuLAAH7qojAqVurSflas7nGlZJ5U8Mg2LW2ic/W
KQRO88D2P/qhr+P4qYu/5qg63fFBGrs7U8u20xOAcCx03MPjuY1fKnd2bUYJqZIe
GUy7LRLTTTGu7GMOFa1f/ilKqv8wVS8uw1gP+dBNZHdkcHuJvYwikC6Gq+7MJrYd
SMqDOITlcHkWTrnCA9W7SQviLMEiQnJbNjx35YVikxC0qwC9pf/fxe+RjKe8o2xI
3psB2JHNxnzlt8FVuTShrYY/5lhx1LzSlfFy07RTd5IgWr5Ezz2MmTJMfCyMiKJT
kspzjuecoCg5RqnHVNpW2lQ7K0oSh2+s6JIiq/o3jqJEWGyFCAmCtAMtI5GEF+Pg
ExXA8YDZxCzIzSd3SWv5D1WnOfagKZ/wozyR6t9LyEEABJ2kEHqyuvzBXrYqqjPH
fywvgG/te5getKIjZFbzmU2rX7XFqumNdPdGp6a1QPT9Rs13OkNzzYQoWBfhIr6u
IPqgQFdYZqAbX5FTOLAaictcIDP/3Nz8X8uggRvPjgaBmeDvR95R01eeWgaoNVjY
7DMz/JX9sb66MyoO0qYl7H9bnJdDElaBWSh7SaIQ4qKVkw3h7gIdg22skw6SaFvt
jxcNeieho/eC2bLO/yZ1rg4AI/lj9ExIdCtrMINAko9vKvXLxDhU3Xd447ONf1BU
MGzJMMofNzyaAZHduzQyrjNvz1ZU5NP6W0eUochxGhYwT17Q04eAkhvLS7LUOX1E
hqONjTa8QRk6lmJHl7fAUg/wac4FtXD1fTjThRN5HgDXpVclIggGJKuo5z6BtLSj
7LWHzWdZlezNnptM9NB8jSpS5qhJOg4K0YuXgaVJiy4rCZPAELyeW2lA3JSMswPH
UvASFDZ4Z5HiLuqZzEE2aRFGhsT4y85v0/AyJEXymxe/UGF56uFhZWqkgUNKUN/v
oRZEfTj4I2TqijibwncMW5WdWMdr30JpeVyIM3njMiSHWjWBIMi+M8YbAXKln6n3
+iii51uIz+4N+qD7n1Nv03NLO0Tqs8Ynev8S+zaewew1CK/mfDQt3f2IT91aWR9B
cVoPKrOxsOhdM+9wqGJswjxOmve3hhIRodznjdKbnwS9XvW9lHv3hb5igG49DHAT
iX6rhBFhIiWliA6XT43XxBqjuT+r0QIQ7GP+0V/Xi+diLbolW8FEwGKJrdCNfxd0
b2IyaEx3n9IkQVY9nRFuuYpRlN2gO5borpwIr5xRBNWlf7TgotmC5glFD7lUacLa
Dm2A5ZZiAIpGXBIoVP1Yb4L+9fgNp3khoClDFaW1v8q1jBbHuToAVRBdgDrad3Rr
mMXnbuIFWT0A7JSyKukUJGC+IhmpTcGvbVfhMiSM1KH4AvfuBw2gzyyMtAcv1v2d
BBmKXoMXw5hW7iz1vVHe28i/Rn1c5fHynQvNUwail9oB91Zx4ki7MnZhA/x2OeSO
zuNgjABhjnkwROP7VYe7Wn1HM/v9aRYZ107eahz41OgnpvvtA5r0y4hNsxG0s8mu
zmEtusg0otnZqTp2HLteHrtOFZ1bwEKEAoCtnofuWRBDlFZ7D/wODeW4A4znVwz/
zTyIlNz2HcYA5Ca1BxDQzRpIuf7dLxQhJ8k4GKHLJ4TxaLtXDpIUqJEi4E3zymQP
exYP1ekzlw38BAEFTHU+rFFO0bfrRLp9v6F9LL/+jp3VxZKmh4bfwDNwFUX3gzp3
2riQKgXFe/e0fgjURV9Nl+46NnQqas2eZgyK3P/LlsvbtPj4IxZV2arUnHXKa92Y
gFQq/18HlSHH47wnudLFpgex/XZ0WU2RmkfU3vd4rlGBio8Pf2Eyr2AWcJMc4jO9
8QDHrQuJ1yw7v1jZG4axy4bwgLO1LtTbuvy2bAJkvDgmyIiIXX0KRqBG/WF0Iawe
kgt+uJJ3jjh2kfi8YNXQwtelUYs4FuoUO8ZP4N/Yvdrnw6LQ25HhCqTvwgbsmUSg
/31OEW1ONd0X4WT6ryT2SdSiFnrxl50t0CWL54AULr5hp/G5jVFk2U45+Ic6kPTe
9c8/oUYGiIDbF1qToUkP8sb1EI/bdBiEpvVSu0DnVXgEmXDjtvWAPES7dN5ft/o3
7IEtP58kaXEy64d2Ger0hETA8/LP96QcJ3/ggWQmsksEu5WhxM2wR67YI6cHJiSA
PaT4V+09GVlyHvVlnr1yy46kurMqC+L/2AJJfwD4dwJb3pw2jugpUxBK0XDt69Wn
D0kfA081WCaxAeIkC/bYhn3hcqVK3Ml7GN5mpy4Y9kgBVu4SV6PrUeghnFb0Y/24
kWr+x/LoN9GC33hwre9yzqEWbmbQQTeKGCZPILbSiBwegYba0jK8kGGjk9i3LMkG
28hysAhCNpqRLRRyP2gC5L5/zZRCRt8idOlpTwfmz+yzfokROHpOAIi9MYyJ4o5Y
CjMaTofkp50tZ53PhY6UFGHHHZDY0Grkv6bqyX8N1R20WgUfjOt3xyQ2Kuan4xq5
xutvUtWpOxDL0DwNWURk7esCu+RO69R/RXunfMpfpOC3hMJfoUEKpWIBDVKzwPIu
ruBd3SztyNAFPAvjkx1eQ/gaBOnk4IjVgFbBhsrv3ugo2f1VaMApR8swTvaLMN9b
QDGgPRe2St9KJet6uVTjJV1ZYq6+osxr/hKFUYom2peosH29NU66We9Ohh+LXxwX
230QxoA22YerJx9S7MCNm6mk+BhWltBYI2DcCczmuThiy8RfJeeubK8VPagu5GEK
GsrsjSLApOZbqccpFDn5uaNRFd/jb1seGJ29gmx8aSe/FuaIM9yzlAekLHueRQsH
7bUzI3dTFEz1BYPmW8PeuEk7qgiVia+HFZkadish4yfAHDesa/3IY4hwgxp+TZ/b
QQOjF4OuJjjnb7Z7H1kAI8TLWSQCV1dRAJkRtynW/oHf5+71neOkCEPDC9S2TnvN
ivC2HE28gnZt8nQgwnRH5yyUnK6uX+fI9Hrim/YFNHl5fNY11XxUWTdfSLLvdjkX
fwFU52gVyWFikolzhTvxD/GI1FmEG7A4m3LGV6+xiSVFLUcx3m87fWwOE4m6A/T0
iRwjl7/HYumFDpcfWItt7Fw+tQnugV1ZuC670e+2y7uxULnbjvORsINfA5Sfk33F
aZJiRV7mu9IxdNNkxKSJGFpWac6rdBplCIFxqbFAB5AIbTqLzih+vtBKTR0vKYnJ
RcqNh27SJaEHphqqu1doYZXYXJrOMJSnszz55Z9rRTii4BRzUFnK6hGZdCYYHLJL
v+xLDkVp14t3a1rni63hQ4SVALwHlTi25pSVrMfm1f+zFjWjd8G2+9dbzScR80Ir
v8IeAmC6dqOpvwD9ReUUIfaF+IITee9JBWKHwtrzCJUpsTDlQ7HYIWGpUeqDIwCQ
aFLKiFQLTmZ5ZKwgF0YmSRyIFQjLxZlO6e776KUhf71K4g6OJ9mzvyKoImouekqy
dq1msYOiJRCEf96Fmfti8BzH5gb2est2u+EezukfGmY9HMFoEv0KeWRNkokvSou6
pGDv5nBhpENSy+C3XTvnwQiVnXrHFrj6I+Ci78WgEEXrepNQc1lF9kXTTpaAd8IR
3oZ/BldIgJRVAMlGBe2jS9zb2QTMEHBrMnk+LWHpl1hbqevtpu6oT0ehSPZ+v8KI
twn6Ux5csKlHEqIu9k79mfS+cB8lUyHT6/5VCLDA2/heg0wKEpx5kgdlpcap9WF/
RvSi/jR2gc/3CdX3LuDHGwQwd5ZA+qkFkwHZ2Im0RqFFbXZoxPiTdyI1tNXX5233
jomF91ve2NqoFmgVtU/bNDa4GGa51r2ZvGpFw/MF3Bxo9A25rX7qO8p6qxpBQprD
uLoEIf1RWTCkWa5TI+mG9Ij6r3Cqx85WLSiBS3j/oMnCUP1LP7B710pGKi3WDI+s
VqqiP06sfeC3aDn+QSk7MJkke3e6SR5E3ka/ntWUZYjgmses4VccTCzXhCDbhmWM
Gvh+XXyHAHy94KTeaDU6tONLtkwrF5UT/s0FExxn4OqNWPF49S1ySvHuLGRDupyU
dlWWSlrGeOrw9I5cCkoHTvtyV8nN0cUWxCb7B6Vt4Lp9oWHb+iTu3kOWtG+7R+n6
of+HOc4Mcf3duw2Y4Dr0a5gOw0IKCbppTW6TpP/zuYXwHCY8+gHgd+jWoN7VhO9G
MTA1dSbvcsTKaSV9jw1BAGRbEdbjKhwHG9A0TCuyYGJNUK6o5KJoEw9E8AK/0kyu
00QDD6OEjbdz4J7ZnCkCZ+52/AG+2US8panwqa6OFeMTT40iW2H/dVeJomCl6J3V
DtZtg5i/IVh7koOdrMK0S/ngOZbsX0Gr4T1ATaL43qVpWdZlvPxLxN1CfLxplPBJ
G3M5/BgIN6aSkwkH0jUHMoUkUDMDIWWd1OEOb5NQBxI+Fnq7l5zv9unkXclAXGGa
Sr1kcnHVetEx1O8VcaOJr19nJWN5JLWxeTa8xnI5O9JaRf6RDHFjpeyNEy73KyQZ
MiWrCeBM8Rywo1N2F8ddcWxjO831CgtEuGVXYA8nICFHaqGsnkPtbfqPvjq1ye9B
Rj7jUUfD1JVVtHq/qFyLss5ulC8vcFJY7XrwwvX2qooGUoTYHXxPeiXfFNIdsjFR
mz8avBVsW+cwGs8WxIX/ikhW95gche08d9X/a1MGqIqan0pBrsmQNmznXv5UK3qq
d0eZcGJph32HkR3NV30SwElh0k5DnzOOyyrqMT9MKMNF7Cf4Hk8EcoyVgebdfB/x
IG5DXeqY/SKHlseq1UAtJf0T5t2+Ah19NtKdzy+7badb7Yqik7FRM5bAPZJvnqSc
lCPb0nouHuhpRWRD5AFM+Xz2mdvqBzl5+ZdXWsN1L3tzmrLDVbKcj5zA1QWv9GUA
rVMmvb7Ia54bLuO1H2fJLHrCBTDAPE1nKGpoO4ysor6QseY7E8Xw4OdlhZF1cU3F
UtISlvRZe3F2XOFgqR2Iku1J5h6blWA49ggAROr8LeK8XqM2Kf1kRsATDa92EXlO
/AR8Y5DsdgrTtzEtaQY853BR2WyBRRDSohfPldT0g87rj0sgzC786kCjnQde4g0L
1x0rfsouSSqyLpfUZcbXKLB/nmtxd3WrEqrD4Mf4/3pR2CJKP/8MmnZ2Jg63vPS0
DETxpPygaYKz0npJcZTwF3jqHI54VNwdOrBYfTbqBDhn068zfI8+wOO7LbcvwzBa
+pkWsJTyX2GkXYssALpLxySJ5LPUYsKFk9ifHFyTL0hmcRw0rkTFbeu2I4Fqha6E
TDvlPGHTP4WRsMiHfRuF2bqdoQVyfhRnX2eZ6jKA/Vo1WmR9+GO1HWt7C6jmq7ca
i8aIxwWqwysiyXguTCzEQS/MtQOE7Gymjli9EPybnrBJ/vhY6+zGSFPSHMRHlx4V
TvceWY39xzJKcUbxkw3aqsyADlQWC1gjavm1v94MEC7b3TvfGPopELg86eLSzf9u
n61nI4oC1RK7cj8Kr8Z4+elf9OvzKi4VRH/WrOyj9lYRjIalcuLTaEP5J0WuW+6J
JekvPJDkibGJRIOWSl9GTuvGTQJioGOJ0ohq1VndG61JR3wEg5Ro/Szu5qW3ihO+
VyFzv6R7nEh79WTwNgJY3sj7uW9bhtFbfjI/7G4dkoL0qNxaN7joi30C0DDysvv1
ski1pfG2O0DoYRB8E8gOMCwEn5l1pLOAMl2S71uGMqARQZPPN+8e8SCgtgrmIos7
D1i6bRBtCM/bu9nYNfcvEs6NFHsIykK7nMKvrTr/5pf2HXCPiY9c2AtJMJtW+mwq
2pDmQ0cK1n6UHnzKRbEmNyN7K5FEkKHkVkW9O6TG8fcnSctsotvhCauC1u6L65Nt
47Q08we3MtXamUaLQGZcIoLw1aZQbPAMOTW8LRazh/RQcay2o1jOliEYJ5O0Z4+7
EzkJrD2CH142R7CP3298WEXO9qxSAFKXNaZeQhBY1pdXfcOav0k8n5vWAcEbKaJ4
apjjL9XbXJ/YnRNGZAWJ7fhfVS071OjWd17OUUWmmZDtLG1UnjuxrfKuZkOYPm+W
01lC8runAnWF7+EoMpp3tniJ/jIa9kM8to9C4YXESZavVq5PBIC7ATGaw8F9MqCQ
mpL/zJ+hVAx7l2HH4j8oJCOrW/Sl86jdWfB+NjTnPR/NmWBE+PWZdlnMDiSmiqci
WG7djNctSzsB3OJBeclGTsCZQY5n4XASMH6wGX1XrEnDNSAJltK5/hxv/nQSyDjj
DvgN3veOA6+Q5RM6+lHLH5lm2f2tG1TA5dr5qmWaORH+7FiCaf3l0pqU6b0fRmp7
Qxdhi7jFtHoABdHOoJ0GTIFfsrfazLGAnFDWDqaC7UJDR47jAWiJBSbMFrJeXY1/
7gOqLKuRq7a4nDZ1yImrrf7MqiW9RGxM75f0bxN50c0uZtZmsucs4vqv+RKMAI0j
nU50uny/EivO0BzGxNEn+O+YEkBYvCuApJZqkO+fHRtGh6pLUWPSw6/v2sQYjpBh
wKDbE7IxMer4UZ4dGPQ/Cxp2CW+K+2Q577LInDU1LllvtkGlU2BVuh7eM8+VQsDr
16QE4+ijgonMN8EznLMF2ahgl4IT2V/GEAMx3BerU9dcttBm74ONTz5EuWP8d9qp
9mKXxOWGCyOfR5VMH80ARj9fBSyMBfFFBDfstoPlA7W+q3N+lsxi+o6OUzgKqtbf
8K8z7/xF7Gr7YlZY1+PduKj3KqvHMR5DOW6Ftssmwtb82ef2ppOWDur077gJMOm+
CefCJDiSIlw/BLqLdMGmPcgsldyMlTWNOjFV2BsRqDyYTBI7Ox4mWs170pYd7/5O
OjfukTL9WdEhm1pfY2N1cduILOBQEpzlol5WiJiNDMd5/BzL2DF7Ek9b5JFUnZoJ
jPA4tUzas7VFJret6JfuMqbEIM96Aq0rGtYynW65NhFjT9ug5KYa6EyGwk2uPhTM
OXmtwUZ/4GjKkV1sqpPjnNDhGRBN2bmwN5kwVwd24XgbUsVLF4joxqfwGVgBnVzK
9Z/ZUsZgUzpwn1UwGV4g6GhnL7OG1KAWMFhO18C9tjyGcpAz0xMyAcOYq4EKBgqv
s6ab5H/k0kymx3ByGrYVNh2KRxAoH0bfXUyj9O0kZPOr0rVAAUkAvU99uVi81o+f
n48GEFA8c/zmESdGGbmegPs4SrbeBHX7wzasrpYtYp0bHA+k2hO8EWSUYUaJbEam
P4TLnxptFd3lJtwN+Hr3ZIyM2O3CTD+dZgNpHWfJEdW6fNIqlPgsDkIcjrjLJh3o
s5Jnu/gNaJAgBizbsh8tyaeV0Ii133PCt/DffowpRjjf6OdayO5JvrCnkzoxmmAM
srudd0l4eRPIRlRO7/fldAYkmjN7aQPng0ZxB48enCzRnPbT4Ti/nVKCZa6PgkG/
oW9tij52D7BnFIrBPo61vWn8NlJxeR53rFFGvtjtLIsODOIlkq45YcP9RebC0Zga
39+ADy7mHYliuXnwnov01u1C/hq9FKVvvsF5ZrgFpNkGn/DjX9I+RoOVJZFUppsq
sg+gvgCsVcxUFgmb1tt1mofW5qvuyA69OGJ5YtfR/JQ618OT5FC9TNhv1AEVi9XF
ueIG+wZ/c8+nBz0/FZe24NJMVcMSXCt4dNMK1hCAoEIqD/WG243XYVKovWeHyjrm
sedEnxFIYxa2/wKfX9UTJFhAbwHpkGZdL8+JfNgBTTg2nw3Scjpbn4ATvpa+NXPo
tuOCgE77m925MUkQsxnEbGuaY3mRmDoDGZ3+zGfOIVxP3RWu574X0MDO4MR8oOkH
LclrIIV7eVrSo9P142g2xRu1eSXIcH32mUv8x9ajutpfKnF1DgvQOLOguhUOTmmm
jqM4Jiz7LOMqEFeV9y6/9IUvEXq950Aiy0ACnu5IA5SuzQoP2jK1KwaTymQw/SZN
OunRVlqncXoZi53H5QRIiNXQvvJWSIogw4ordJiIembP2X1PuY+RW9bAC4c2zKdn
1Fp7zb6iX79eFYRmija7DZX9sqHtp47jjWDAOQ7jcCZMRoris7oc2eYHfPKHaE4I
RfrFfMclS/j5hnb+dHxMDip+Uk5wBNnLFbE4RKK3uAQDqH2mQEBj/xb0igiTzK5c
hKF6+NdXFIYBu2BUdv9R4Az6gArfTumca8Pu0MDdQ0SO+br5xNTVANO78D6t0hnH
FkSVcoLZZ3ekoJKtu1lJE7Vcm2L4D88natVR3VuJNUs51CiMUu1PVDWONgQyKko/
XA2q6MpSGN/t2T9Mx7DIMgcXh92TyMv22Dwh8gTgbXeGJteoUlbGFs+P3u7Wobhp
SYvJQlAEp1cueESXfnwGPUkUFxts/aw3dZrb3Og4r9mO++kzlsFTYD364iayCvQn
mScYJ4PBTNRekYftERhZqS+lg98hi0MaQR6EoywUKZq/X5SRD9+DG3H7B76Oqck7
p3bWBKGeaYKVrvxu83YI+rEIXO5lQBoTGOSLPsqAcQICBlKDtLzU+lJ5RxMWdqgV
3diYTwqW76ieJ+GLO2r13aD0gqTW1Gw87Dj+d1H57J8AWOBMh+UlyGUz5Yz7uT8n
l2r3ULqyY0wCncTCUIYWGUDvXS1lfMprGOA1UF4Oej96mxxol2eFL2SbEOMxPAG4
NePUimaxBkMCbPit+VwXzBoRT7kQIPC9hp2dxkdOjiF7BKepRXF5z2W2nQNYGEVE
xjcE3KdPQBqf7442JxBOC8r1PpymydekmrV8n2kjw1qFFyUDhsnZTc8EgmjFsw/G
esDfr9SwaBcBdml/cTPo6D63U3mtl7sVKz0n+M6dGYLcLpAhHZkkHqAN15EsfIP+
dwH9udB8timhh9OATs0UeWVfrA1F6etJ/jSlSkUjVUPDp9etR9EybTm1gbILY+yA
1WvireGlfAe+amojmq6rzRxCJ/UAbwQ9aLVC5HcjV/SYs/Rb+4yIrYxanHhAAWkx
iZHmB+F/ayNC5kR4/f/BIwez/3aPaOHC5HWAzUSEPP2HADNYH2Y8sCrHSs1q1jQk
IHMZeJcvR0Wy6Ob0ZIQpysNyFohFjWi4j/4+r2JS5YN2aIo6gDtuHCkOklMJPyM8
iRyQlANB38k8pugRoF89VZE1YWvEiXqZDWOhIumpbNHWsBDOy0/43VWtkActJMoz
997J5MjaRBzP9M9neGjwAke1ItpI9KJ54bRba0u2zC77b53qFuT5X7zmLcAk5TTk
vX1NUW8HpTbnrpSd9ynNMDJVp22mOqJYeOM9MNQErgpyWuy8Cgw8aw9lOEvq+h+O
QSK3kzxa0ubicpjWeVIFnEumDnGuPRitNlh8LxycCbozkVxEJ+hvVWIHtJFIg27D
gpf7o2faqWVwbMMewGk8cd67ItsITZe1ChfyndxyXoUZsSqxXoAM0rOad6CG0aUE
pU28Nhhy33ZhUcjZUswIcZPPvezcCk/lp99OopWOCiqMiL4LIYeO5Mq72xFo2Wyn
0vwpsU2osRMcjV5pSx/s6DQK23Y+rCW/+tiVSXXDg+dRPv68j/cNClLMwMiBaFZP
vmFXS8VTesA3i25fML+ui4zFOgQBminds9ZUjnCpVf/WhHWzbGStCdGR/x/jTdek
AljXPXdsdmu7WQ9dxRBMUEReznjDiiiOonveyqa1knlOslFrxx59Oc0tMzOuhPyg
KGyuNlETyLZiIrVqq1F51z5ivUEXBvY6wzEphUXaW3FgPvAtYmIvG/+06WzcSxV2
mceSV0psL7VPNE5FW1tOslsvJRFjnw8G13B8vvoL3hAlqshXkFnrfwYyyudPqN9G
O9IOFg+aMylqaPkKYDYUPLIOmlNNHoeIlT6fVnZn1w5bePs7WfgT+Fk+JtalmZz6
UQBYn27MheDe3Uv4jS1PeAJkm7euktI3JlF9xjiXubJk3kESI/9fxxm18rqonru0
PtSQ3wNiyIaPBf5TCGYtgrRaXT/nr0nZYpPXFm5mRagHBjgZBtQZmmg5ec+03rdQ
D7kCQFNLgRjYA5zOjWDwHY6e6DwFMczjTn7LqYWTaH3qliGAKb/KwTnHz74xfVdv
/T5mF/4gzVFgyI/WR2ZnqmX6vjq0PRfQOx3xh2ViBo3L7rztRtzN/AAo7wwQwrtl
OUbn/HiN1JD8aq5bZauwvU76u7LHZCmKJr1XZF/4N4JbDwPw6bEHY4WG8ZQH8Sqm
mdgIWHUmXWcNk04BKf5gM3TJ6ZDQ0JC10Yu+4v7Kvp2lRoCJ8+P/IY/5hTnn4ZdR
tFR5eGj+WFWwNtd0VGRc2WQREwOhMiSbYSScrhcQ8gXimiIfeVCnCQ3OPmltU8Zx
2wzuJrpZ8RRZ1/AB2A4Y4u0ASdUYKAldXFVvdqTcbpXJSbAyFkAN/yfru4ZUCAjs
aBuEp1DneMus+DKHw9gfz7OCBcS2+oTquY7WM22hPLz8aNqxojnwPJjPvfdmNgc5
f3l726BFNCejIO903wpn+ncM+5xTXd1srLvA6+KhYEDmoMTho/WoAGaTOuEq+dvs
etONmd8LRrY7F7rm5OipuFjaaxrYxr5dewSENhIpqV6XDrLgnPlYx5YRmRlaGfBJ
DoXoBLmyRdDyalSCTBMxkM8v2NnAjQubyxTMXweWZpa3i+IM22mt9D/SWsvgxqqG
cI0S3vRg274eWRvQpDPjWuA9l6dsl+MAAfZuqiSvP1nhdTtt0Z2hdqS5gBCam/LJ
aSWjw7C4Pca0s4jfL7EzB+syyjSl5DJ/j1lyrX3khGRAnVcc1lJi81FGgFxztpAX
aTSWShLD7RWkUz3S8SGFgNOHRAsQ89+7HFu3seSfw1cE9EMWO+EtawLvucm7J8UV
OnbZZ6qKxJrTlwjHh995wMjoRvF2YXFCRd2NMvhl8kEk32yWJoRjJ5NTqvC0ChaA
978ys2ZSvK/YZ5/4x4fmpOm6w3XdYwlFOUJ4b59ZOLS3PgWbavGN3NReyy92apHT
KKU4M4na3zLIDOT1e0hTFAmflL6eeQMfOhxPX8ZzWtsUnphZO4R5U904fo8J8deE
Ua1+g1IPx8mJTq6TuEQY8tbldBGbRDtlRNOuS/BjrlyUYLSUUCMHO3EZpgHaCZja
7hu0bd3azF1iScnp5DjJ9LmJtjrth30wdquozuS7haB0Jg02L+nKB3QMXsHTKnDy
twQnvvOfW5iiE9fgtaOA5rhkZC82qTUre8+Xc+9gfQoSaUfP7z7m9QDFRDzF8Uvh
LNS0IChIfEEOt4BRnE9yPLkaGt/9QZ6ePFBC78ds/BytJ43f2FlWxn8ahjvT348X
Fj/21pOWeO/mVZDFd3hJyq0FDSjXh6TUPcPmkgFI1vTGPq50COGX55UD8EWWj5Lb
Y87LBPAVc72HItlgkmhL1boVS7FtyprVW0onzMekjBPKV/dmiD5b6upi9Wj7yFSC
aJiENyhPqH7mm/ERP4wg9rq7nbpFzH735EGeWSse85bnqAgKuAMgZ+W48hb35NAA
kDrIs7OBc2evsRSZ/aPyVATJDGQmP5Q+X2NIFYnR3LgDozlTx2F+FaGsG0mhfhoI
dOFssiuu7NR7WU8Jx/84o75u0sv2u1Q11lNDl30+c7faYu9BeXIZJtml+tAzgt9p
ygucara3X3znewInULTFoSY+yiZjZvChCPOhqN6BBy7CV1qx70PE7wGYKDCZMH4J
ftqzoSwlOdGp3L0vK8uAY1kZl2szgJNJDdfyh2FI8x+4AyMMdxbxcnPShCsngMKu
RP0JRBurw1OP7MUzoyC0o6YrYUJlSpZ23aF48W+Dbb4jcyIfYE8eY15qs4IdYRjX
AHONAlc1FH+Cx2a2jxuin+L2yK6aojFQ1I9JTkdG/BayKouhSD+Kp4b2S4VVmZnl
Vb6fxPtAcVseWEIBZuoAE1UCycNOkAgKrceOiHmkQDtM8lP6U821m0xTkqHam7yR
98hvWnndIv3Rf8z4PFKu3rPlAYYFP/EF6fjXrla3TyK1LdTygdkI4Wixbf3ApFPN
Ouq9dsbc+rX+M/epx1AJ/PK1JClZt9FUXM9A0IeI9MVLVUO8RxMiupScI5tceoyr
bYfNpzNlQqyamZpuPI5KMmVm9rtC/S+Xc5T9g89Kolnkf1zC4pUI3OropJPvJ8J7
ky3jeRZdI/DUqooUWcrlM417HFri0lWUsmUROc9N3D2vl0dtQYnve68MQiDeDiMr
5qukVNGeGuWgEWiQFuWgiTC/sE1tZbYh+nR3P5YjmSWc/ie1RYU6IAf1VjfXtyD2
3vKbJmiubiooxqyTmixUZAz69NSeqg1M0x4fKOe8IXgxCwSDLsHj4jMIHcs2X3qo
H0yw+WMuYMp8YT7UV+Z0ah+YHr5bkoSW+s5N9lNz5PhMGKfN52jpnrn6FFcf3ANp
cNgjOtf5GMUp71+8bIOcFoMEWm6hvTW9o2PQfQAXH8nR4Z0oKR6W+LupSbfPDBvq
EkExi+yFJeVdfYYO5VAfWi2HGVTGxtGG/KyWsZtV5FbN5ruI64EonLkCIgIQFzDO
U5XvpLG1U7+5vxircF73DzknWsoDmoSOqjL2qX3xhepCy1C0sqSzffp63CUUC4+S
iWE2OZQXZNOTM0r9eAXn0XHV4nSfUDtbce3GBbBDry0q+nPUEH9J1tfgGQdxXBEI
NlP2fw/ahKiXjIy1zHj/bbe15Y/TM0+ADxfrj51L3b5MCquINefzPCwrQNyR/DHj
nO32kAV+WQBQ5DYE6TNUuUhYAYuqNusxihBrEyXsXjyD+E+UdNQ/iSi5qcX+eYN+
kkJKtzhNmbVN6KKE9cQuTGzdt2RceQp2jOOFw4Q8LD4mEe+//YjU9xImiJo28y64
f4tNJsvyvV+sn8QcFL/TfjNNu/SQHhnZqIrUr2mjjk5S3ZofO4f8St7qS0MrUsCp
EYB1/65cXtcUvnwqASj9K1FcxuT3QLOArgkMlm4z4YgZr5giXwPK6PjrTfiRntP/
UMWNDKtyENte975lNPTLHfEefI9Wd0ojiqAdIHB5Fj/B1vzznGSeItPBLiZSNNbU
Ye4K1s5UNP880OXpeQ11hgOsn989RzrpEZMhdYN4Md41D4JwuLgUBEOXIDz0wbnV
vW9HOkh0nK8EeV24bGQ2fio+l7OZxNCuNPDsRyWyG3Ym2bucfc0bmoO5XDL1BYkk
tsFhcnbM2uPMDEmSDuWrjlZAE0hiYIJdHcmFOkipkkjD2Q7DRWKYMdOIrhqkDaV4
ey8Fi9bYh9FfH0WeZ97ds5jd/DfHcIocd4llhzSfOLymsmeDVpJaZU7j+TVrsoJv
yeoE3xX8aUaiFF/BWK91XKSUZ/fUxQVrvMwiFN0KuT/ljnBkCVGAzjo5BPYCoSva
owCNstRVJQgWtUXLmlKTLZ0b4DwO+FNJa0xPzItmDvVCUg7+Y+ozZmgN9tq8BpKl
W0iQ2oZ/28+fb7W3v21Nih0RgZF1gAoqWU5iIWHFYFnXxKeDxUxGuyJjmkRpMmdP
Jwj6cthgae69QPYvHyEdRkOcba4p7vetxMxZT1MSChGn9NDKDMEr4ojm69itUuNT
f94LdxcJvja9+epmcNkyWYeZadTXEdRsyg+4WTLMKDGnLgGTzCIw7ubRrB1WhUoG
aJumO8L4s3sVoO3ELvg8u//bK9qKymkpD4+MqpzvLBDrWRy+p6ELqTZFRu9jAEKe
Bwhv2Y1LdOft5S8GHd0vRVnCt6E/TyhyD/yNLop0OPDNj1giUsRsRNzwJVaEb41R
RmHg9/slRkG+m/+zfoTvSkmZVhHlrqhtmWlK/seDbpq/UKne+r7phiQbuOekvpKa
1tuuEf/wORsiJZz+oShmk4EJoXNYMY/WNtz0bZbv4M/bbuOoFKsNBQdVHPQPGRQO
L1VJJ+/sLJ9cfKTRTCs33YyVHjN8YKedI74/RobVuJcLJuZJF0+ruri+8B6kxfKj
40nWpQY32FrIFprxJ+uBegdnbvLApjijJVsRYqR9kpaOJm676UzlAswhfFqLFCSC
VU7vYccyY8spk3n5N9utrccaHFRdFIozKAmki4J6GiTHkv4/fSpHyODT5rFOhUyi
JGCN+jwpyko1c4nf7TSr0O5jYbut2v83MIWGdk9vLAPfeTtMoIxDrD9b3noADlNz
uPYLf5qC7ASUXNIPVHntiTdtrt40G2Fx6rQG4JfSHRGsVbWKt+O40lUS+AfOA/iw
aCE6VfA87MQv218ERO4fwVpRGukdfMwauNMCCw62NiUd1gRkds1PmBXOKha/fPuV
EZ3ooaw7B4F3gXnuY45xLF2DYTXfo2/ZblUwTGAnzDJo+F3fgQRzdQJ2Es83c146
D29dFOUcN5/w3uKUfQKg9NW9PKhXY16mzxZ0+uRD+xYx/Ihxk/2rPi3xtp8AHRAP
cWnvwyuCB5gmoDAkFIa+gcQX4tdbC788fsQWTw3hIzYw/RjOpWCtMJYm8U8tNvG6
EsfgB14RT7fydLe/RYJAJPvesZ68wiIZns64qIdDxMW+y7Vmd611doUnMy8uc/OW
dhbwWp8HbQdihE8xKgj8Ic4nZqM493mtN/KBXbvJeTAcubLJNOfIBFapAlW6dgz5
/Qypt09L8V+60OgADjMBAhJpcW1bpHGGiKnvrIwUCeKTK4MZQKizFAeNVFEq15za
XbQPzUpInJZJz0xlgm6jZrp8+qhU09RkP2IUR/IvhIb+vErvEJ7cB/WmDs4RYOAB
sf9vB8AvHO+TXYSE0VlcxE8WfMUkPItMt0lkWhdBz98eso+mMOXweO9D1JlsBwTF
9NUZPVPYdnUB5DVNmq218XYWVkYnSyjugcsApCPeeUeqmhlsD6JqXBSZhEef89i0
NX9nYvSxWkLGEHjuSa7GFFrip9GymmxcG+ncFiDZ60afSXH52Ab8fjsQJmUfSZ62
g7Awzzsmjtq+lszRkSQCn+TT7UYKOgl6v9hqkxaSqcZFILcYwyIiDoDGCQDaS8u+
Sf1ZJpZRoxG8tXnuXnRUsV+Z3KX/+ucIxLDuPNBrbAirO/OnIY1BB+PejAG+keO7
fDSmcYFXhwwIPPTYkp+vCS1t7y9qZf3waO7/KM9aFQVXKsBT5lpblfPziXffbTHs
sGr3LJbX+s9z4zqHKMco+FJucJNYWB4Fa4MAaGWPdiY1m/TXVjwnJ1hBSfhc/3I9
wm3Z/vwNXOA0429ePUaYk/RyuPNQDieGdvOcPERCqPf0fjrRLHAYtIHogi5534WL
+UjQcTzsZNf29ETuU97IktQgOpkbfLeO4zJK39GktTInS5xwtFqGMxTWd7kR6Vf6
cs0p4QLSIXsQjJTjbonc2QxzwPcUxthd0pQUr59wj6Cywl+TX8J9YIJCMzc1jtFL
dAfClgeXRXC6AGMnZsw7V2aOro84si7bvk6vbiiW65GBSLsQu3KUHBH77dRJ9+Ld
pw7T2XEQ7oFD8ic4sFFOE8Z/dU2+wcaB1KuW1Cuqsh5xgk/zMAMoWhojYX40D8em
U8Kn8F0mEaXWj5kEDjQ4xvEQF8kxfwCfVykpJ5w6dANb6k9Gn3e4UgISubRzuu4R
414JeBK1nJXJ8RsXRJp0EK08G1/iBAgYEOdxdZBjN8W2TjNBqbvjTzZ2HlGi/b+n
jU3guf7Tmv/BN12XLd+EM8yYw1Aq4V0TUWhBCdXQPnqzjnjifL1sqxuOiFBqGK0I
OkYNtLCh71e2ArXkyS/nxRNBXVbgmrDQr0KVlIhK4l9zrXYaxu76VTxZVudf50Pm
EmhzF0EvBxj9TiiSP2L2Vk7q9g5cY2gVRrYGQbSPHgTK3wGX5XQNlisI+Tb71i2W
QGmXzp7R2ftq244J9DUBkITEpkbcu2+QjxOMA+4fQwAk8B7KaFbxQwvd739MnWG4
ZikUR3vj1oG+YlqdFDJCmA1MqEjPm/LgayZGJCFIUR1IufQa/P5Usjtabw2PtpCC
4vsxmTO9qUOIbrOVn6pILGeSyuYx0+NG73TyUIoQ6C/joebVyDKzq+VLJrwPT2bR
e4NQqZ17EYnMvfyutZ2bFfYWcXOid/4Mh+EnYjnt2hQuEN3kmJuSRgV3IeVav8Cy
XpItJKBHfTy07kK/cnqk5+JV6dXVrZIrQPL7mqGQQNF2qH40P+1DzRMMDJNtOA37
8FnY+ARYgjPPyLZCC4OK7O98qYKAjZbFgR161bcoxVCi3Ly/6t61Khq45kbvu97O
+ZwBgFoANV26qWdsuHDJ/wAtFaMNQZkpghb491609FeYlWoYNBza4jpG//GCq6fk
JDHOOnCsU9H0wQyRQETfD/kItUwzwvnmaj4eBys2Iy15HWvZ3gZaMusO1v1lwZ8j
nL56kNLBaffjzVulLztMrXnteF6Sv95sJ2roqG6+VQHS+0DMi+XZJjx/29f7BINy
6cq8+IE0UegCbTCWwaFsD77qazTue9xTS4DpUtkvPjWReP91XNtYzjpTYBPniPpo
wIX7y1pWkUs9iPUnvRS5otz2YElKX7phWSRGCWJEnAIM0SOkoBC1qnJmC6NePJFi
CCQdRxS3Ge7O5mcXbZlkme7igP8qRWi2rR9lJ/SxPTWQW1tiSSOWtKkouVvVS7kp
CXdLTScqt/ULsemAifjCiAb8Io+HBDUKoZgHUBFGNLXkCUq5qpTX7FLPBZNQeBXc
hABkNznvawXlgxqOuWnhFpMrkaYyGRzc2pNP0T0ITKVsBONgmu5TKmE2dl59boRN
pC1BwOWMSNIZZ0hSe3vBR0yxH+aAEToRZmC9rLs7z+B28LQQtVWAQ3GkOAwFoj4I
iNDU2u5YuKnX1ojmn+uAUl1FycYgGDVrIVYYNkdFsucWz1sewFRF1R8ac3oZaGpZ
7cIFyeet7A06Ul/yMmDw3wSPVEvNqGHmKE4pSHdsdwn4ExEEPISpYKqIv+SGECE1
nWCdzXNtVd9smI5DB+ChEIg1pzE4kIuFPYytzEf1L8aHRgD8mPQInK3DO2FvHvjY
9QkugnkOmk5cItJi7vKYSVuJJp5H/7Y12YToouf2R419r29z5hN+SYlsRqnttgOM
fgwzANWTZWuD0FX1Dv23nZHaJ+Qun9xcf+A4B3jhy7xKas5ehVSlapeNjCRh8Igo
V5VNS9XC/GobZlwFqJHz5TADtZKLa/VHOL/l0yMOS0U0pI/FSJwg7pzR18xyJ7U0
4OPnE2/uR8NBDaR04/lPV0XadRlNnW3xPdjw4Ng7d2Q2X1t/kNz7HsnD6RAY9sTM
9DyNbiakydQcW4qi8kcyo4TNxPLXUei+BCG8ftcEhGPYmHa2gswzS1yvTBpeSAMo
LtHn/5mXH8vKraF4UhZZE/TRyDH84pe6m9QniHwnP0q5Bdec1h91AordNTChv7Gg
IQMlXUciZirPsGP6K6CRsmfUpOjik7RQCFbmF/XQBXJeVnXOD8444UwE3fQvThDh
tocH3l3oQqQOIAFIj4pl7030RUANMtO90cOu8+9RAKRUYJ44odHo0eLoKz/6KS91
KiihTlOEvo4hlQRXA3yAV+FJV14hCJIptY2bQKBla5U1BcXAVk3v60W99g8HY1ZU
xSdVxLAbbbIuM46WIt17/8kkCpyFx93ZcWLwn2dVjRAVei8xkU8eM4HRq0YPhBaN
DHEIqkP81lSi+gHQjiD/k3YW47QJu0ABbo1VkwbgMA7SN5xin5HzD3MT5Ygb6RYm
i06OXVf6Lb6X0wuENsx1bgUBsNyWUC2JhMgJpxDvDdVudZ/MjyBc1NIyLLHZQdE7
P+eVtutNHH20sf6YxkfYxJel6tgbvAaTCX4qyuJl5IyId2cieUr+ZNeJN7jiEFVn
RQIkpe38DPP14cYJ0wqS2GVm2XmA+Ld6L6lwdGpegEVtc4yQEer9rko2O2c60rn4
h9ilj2NVfCBveFqWOgk+I6v4ieeCEnu0oTpBP3oHbfdKNFJb43eROQJNQXJcBBuA
fTamTNVpqgt5KkykhMB9SB40xSHmP2xJyW8/A7jJY1OpiI3LqFd6sWKXKrRvvfUT
vnSxlhtj7niWpTWOmg5aI61eAG2W6Wj90B7eCcUFXx12OuoKHObyQlgQpSYcAphN
bR66DBo6iYmAm6UFxqxBCinrRL89Qv4w+MBQPRrf0oEGN9sQ2vlKhbaqQL9dPi3J
FllyA1QLQpeyjmuII6kygBu4Y2Jf/oWVrmR7jjIviDKGR43WbFRT/9lWtbv3n6v8
cv5402SOjtN13L+ndHL7iAEJbMasOnA0jLch7u0vyl41RtD4USntza5Bc/eMOLDf
6rpaZs4MXQwJuHXaPSI8CvvFzJ6DsjOY1czLIwR17E19ctyJGAEnFKcb9K/Ai7ex
Ad+1NCA8t9oqAob3VkkmXbgRiAhWs3PEEV0h7Kv9zoIzy+NVxhkEuaFKjAApLLBo
ucFqOEX0aMM1jO7T+FQusHGCsa3ESU47nIpbcbA664iDlqlbdVJYzZcYAxnyyW0q
P5B16GrK8Olr7tZLExWMQfOm6pw8hpTOY61YyQtzJ1XpwIBtIMMxjKBHh6+N75A8
ewvbdzBXexn+bn3Ch070R8Wb/XeDsL4AWhlGuLxrzSDxweRB1MBxDsCL3+MOIEbp
3mWS8ZLt0cWIAhkTgL6VPYy7Nie/4eThIPpm4S5dbqQpFlZn8kTjyEkkhb1koq3M
BDJag2ue9QU3O2HcGVC6tMkA6tXiVHK+HrMuwSb7kLd5f2fgeENqer+I7dsn0tSh
M3kH1ny+41HltpUSQmpK4qCb6ylwjHgMBUAL6uOdWNeyqvp2Vm70dzNg5QsmV/pI
KbumrBNrP54pC1138VmLUBebaHziBOIpOsjN/ojG6HM1bazmumWx09QcknFzpMly
kJ6k7Wy0TgzgpwBj07xYYEq23kDtzbMGit3iclQKrvXsWq3u7mVaKfmYxeja91fC
mVLrKBdFvy9YuhGNtoj1VR8L2KiWe5CJPdJVWCR+XH2ghpJ0iniC9HWT2NKg6dud
ARE/dM1HabVxE2RRBResu/5IEp0+C0T5uLl7rUxhnA1sDmpbpBDEHsBPIXuzMp6R
WOIFTJstlM8bZMKNq/0IgdRLMvR6pTVygS4x4rChA8GG869FRxnFuzKqPvS6550N
s9ObTs1mwrkDgal6b4K8zfsLeflwxwHYn1dlDZjt7b9ksjvjypuPxFWbQfDJcQsD
7C7+t7YGCAQz4N7HKYJFQdQXsGgsj+jU3d8BTLJ+PzEW5TRk2kCz/bYI13uj6yML
F9q66AT3xr8NdVbkEv7r9DL5i0IoanVV7h5cc0KFGYw2nOzfEa4Id/8KawIy0UMa
SjiFssRzW1Uq6SpdYvxiOreoxTLK7V2pJH6xtQ3Wlmc/60/bCpL458piZOoSIxL9
LoNlqpWtZJb1IVFGiOoPVJwOw2l6ZnteFJGAjddS1iMUO/uWyjstXkaNIoI1PZkR
5cgc1EUukLhSu6ALjKFyxjaCcICN6OHeMdybIXzAZSetDC+RhWNmglFtY+WZiVbk
6J2KHLGvPLrGdpY31QMJeMwbXFycXNs3CHn2n2x1iRT3LeV8LIK6pxktCpY1tZbv
2UUQY+kLW1GesMZciH+sUoAThdk4e5edI5nkoizNBx0WPLjT0h9xQCilp/nYGg1q
TSUu4DS6ccd6zmm0fLSQNp3GAgS2RXCJW4jZwaFaVDI/mlcSAUaJIOtlXsLt44S0
9k7q2Z+lW3rIlmz/vG5Zz34Jc0DnJUdD9ekDH8NNCOI5I7CKgDkHTcmOUJEEh8Vy
9kp0Rnk+9rjgwg35uk7LrQL++3q4oHs1778c1SrJbndTdZ2ukqpIeg2pD3JnUAjf
F2MFuL83cf/2ioI2e88TgVk22P+gXZUb9zhr/X/9gbrDAXEE+USIdU6dMkOJ3Cfu
aOUmzWilgQLPESUiLfs2k2lSWQ8WERILy75x9vDPde+bomlLGL5a7I7ZdUN19cfx
8q5g/whBqzopmfyOqQrPIL56pmPsN8vDskq/1qL+2ElLYGI68eVExbQ19c++B9tH
nORm3xq6iw2I6aDiNy48hTkpBSn9rPCtlUPqPB7u6tFC/ZDvIiY7NaB6dH2aXjs+
q/VDW/DT/KunmWo6YcO/zEUtwOiV+mGu/NRx1GGJVmMBpAlqXaE1NUBoPHXdon79
nkdDxr7h45Gwg7Hc2b1zB008o4gaPd+tljpORyCRD7wlq+lUe1wg8KECjy2XuKQI
pmUOFNOGq5AOhqqJt+P/gfbwwbsVZh8BHgbz1ua/JT2/dfe3EpmSGILYITxNrfeh
j66dT+z3o5Ss6Z2pePZx0TnYiE5dcWZ+7TCUf3BIIPYjp2IP4TFUR991X32MqQkO
l2/48aaOJ3mRFoMSgtymlSAoxoOp5DNNSvC+zzAmJSA3d3aeDSGaKc5f78pRof5f
mFZHP8fVFPr+HwdMe2svFKXidhInHFNKSSDhmKYAmoeelqFJhCX7Ha15cUEcDR7U
J2HnWjiqwCAZWMS4DSLgjqwwdUGHHnaROGxS+MTCa3HfG1P0JLOyl29J9Ui/KRzK
dqjPW2h1lGwohX1F3YhKFn7cxvL2x3YpBWcxRUNMbVy8+IRdHhAuXDGYTprjUJ69
xQlssMFnXFeRRYP1u+JSq3COV8eD0HdorF5/Q5Izlv6UydRu+ruzfqkobtKae+2u
i6+5NkbkyGnNDlNsD9xOsZ8I6g/GRH2yCiiJbOCmllR5Hxsh3iYn6mrZQccVD9lu
n2FgShHHM+6PV4A3njfIXufDUxIG65xG7UHvPUT88pQgXmrZhMZjbBESelo1mNYT
l92F4yIVVqeJDu5EDy01sYembKrDR1ReI0TNofX3QmKcsOiT4ro1CwQf9VfqvhFv
6i+lDwr8sVbGEC+12FiJoZHPgkQMQmuqs8VWz8rrAUcLdor0+1kAmCYmvtfXwyD5
P14pB+ZFiAcFCHYfB4WAv1FZQUm0nEEjDIZjFo5QGg0naTfcoFH6RAgyQfksUH69
uE05uDSmc9Pf25PHGPxaE4T4DpyZKwi7LDBatkCA/crUElNCgUmbtk1DkQ380Em+
o1anMhswMBkeudC58yF+jv89FTrEvJLGAx0dGX3yWJ/BNFojN3MnCRqnDhKAJfQ9
pHyyagdruleul0S/K72533gACxIdXYqV5MdW2NcBvFBTEcpaJczm8dKipDtSrL91
uHD9TYpSuL36HSX4YtBbqTZH6f1yxN3uZBelD97pv2+hAYuy7HenWCCFo7s7JJBx
3Y7O8daKO8noRKX3R5WvXq2rZEb2g0QsxWLNvNo/QnYJLGmzz5Af2uIM76yxQSwf
l2qx9z26NuN5Jgs1KCpLUepBVWKSB8deis5gU0Abtc/iSjqVJgXICgMpbK8ODYn7
5Zyijc9YtpTDhNVuI0QZZb78WEVuTqQE3L96MLx2VqAFAJXTxnAi8gQ3TIKJQE9S
cGWeayMFMNs9ozSgDeH/M/Eq42K3roY3s/O4s1PKLH0z4QAgJ6BK1ORqNQfoi29k
fewFeh/AHK/iDR+g6x+sWCDcdAh/3VNDD1Bs+uddu2nATgReWl01Ncfg4DiG5e0C
waU8hzeQcHwKTnQhqRpXCmZnK/R3QGM8EU4VZpJfPQ4LkRyhww1vb08ItRiQdJ4m
4MMeNG8rIHiFMKXjpwouKDpdOzJaRz7e/Y/XsFuYx9hUUtWL6jgxy5De1Te5YM+N
BO/8EbyMDWNL336LYPIhK1aIPaI8n8d7W1tX+YSv79Ee31dPeMMSTxKUv1iXvEmS
fdsTM21QwWr0cBadX2BNOOjGHZe37zfuEPT08VcIvorrJplzdR94ejvDz4GiHEzv
iYDilh2VJ56+77QTpPLA0/8dr/4UA4m3JZDsAsflq0pvrzFeaRM8I53YRvgy5Al2
wa8WJDYOtNrUntC+mOvlXkUyGaE95+GCRR3cnl2JYhf7a8BilFPOfDwvbyOPxoGl
yyyo5ta6kuw74GjplGIM8DUyxWaMu5dPdiXTYFTrUtnAxm0PUNXHJgmDPWWoIYYM
Q62wOs3vsoRC8BisHhbXF0+8sHFtqyQjXFEJfODYVt8ZfJhZqwuztMgyVg83hlk7
UT7cy82syWGc1jSsWXshIKpz6fQaftz8NMuQjGN7HViWz9sOb1LFVDGZQIR0gmbW
EF9fCGi5zVDVz52AeGMpoEnHjqTNpcj7TP//aVmsUv8YEsYzyw605gK4pA6bRB+T
D4OwyzPa2HjyY5lS3888QsZZAdbAIVkhBBqopW36Zd9lNi+fJK8Mtjfdudll4IlG
N9Yt11GqPPiohqhUTZx4RR7QNthUqqlnabWx7k3/pYErg/fswABT6fRMmG5Pv5Kp
MGbCG9TREkxChCfM4blU3fGvwjlVE2kChuwoS2rdzM3w75nApGaQxTdU+w1QMSoi
hMRy/VJbFY+QaIQiPzLDpfNVn55D3G8tx0INM6pkEV87T6FBghQRdUMkRfgbscfp
lASLASGDQFujr/vinkWGV4yffaU8ehAbvyaTH8O9HFBoEx/TGCpzIz/FOTfZU7Ce
9OFu4QVycbWAVGIfrffoN61eBH8sba1DIfuCakFo4Sh5QbL0UC5R4TNC48kmC3jM
ITKecizOlUR2ehTDG4RoD2wqyB/DV6TW0ka8B2mJ7vGp/sJ7R6OD0/iAuIwoGRtp
RdJ8ldYbt/JPXuxFk6i8Voq7kmQYhBjHmgocTqhkhiNYfZoCTRCB1lDymqvSYlyq
r2XzXzB7ALUBqDfO9cvNQolMaBNy0bEN7Pe8Vb6uXxq+8a9CFgGtV6T/zzwFS4gM
t9jxUp9b2Wo7eBaOxJ6w3wexZZQxUWJHnu3G47/Pk8xbUYIVPqyuQsnhWW+p9Pj3
up/Lqwgv6EU97R7OHHDWNrloMwQERoKB/P+ZMkiFs/zmR79pBqVNIVK72FQVJXuV
xxpNMSXHyltP4tjoNSuMeIllwoBAWqy8PqijM86NBDDWAmScWK8mFujEpxFD4YfA
8ZY4DXMOxL5Gsr128PHP51Awk4h9M7CvXG7Yf+ehUR3MyKeRM8KUb2RH5z0VfwyJ
C4qrDhFYLjDK01fBSIuy99GmYsw9auyc0X7TgGuE1GcRuYaNeSJAjGIVzYtPqxs6
IPOK6375n2X0B0psq2ChE8yUhXDIKTUEzQtDmsjvA+SwHxnMYIEm3KiwhCl0yDEn
E6rju8HrJ4Ld6ECAuagGkycrSLkjI4Yd/htl4Jdy0YRePkyjuKlwFm5xJ1DeeL2U
k/ze6uWuvLT494r3nOuMGVQu+yMnCZaxtq9P2uYk5NcdirBxyDqtlzFwlRP3MwtK
wVTUKmEsRXhCBWOWRQRDV8jKdnx2XOqRDULgUxTWwWWXjnA/Agp0fQi7qr3eTVah
XpqZgmOppnFFzRj3bKQJLGcnjEtOeYZFEUCL+JToIref2RKgkAlSXbr0RROMqDbc
nlb9loOvsCHYo2hJFhkrPxjnaO0vOS2IvBggbVySeeuLb94uQBIN1vcPd7VIxC6K
QZytt8gFSpzCq90LtdeD1ZhKSkmpVDkmFTyGKIqoJactjqFZUhwtWwIrdNu/xcRT
G8OWC3+77dF3AE80vJsJj+kYzWd0dszvxDLQbLHpiKkL7nshOZ+vtuyr5F3BjCiL
cEtCS/U1Pcdxr8M2XO7SnCmnDL86+JcKJXrfEzNLQULTuNUhC3ZeXeeVxbinTSSQ
fuaXgHmHlKTABkxX0GKcOuHxxi11fLfPluZGSCMrw+oHO5GjiPd6DCWoJsGZZvWZ
XR33inmAesnGGSbEH88LWo26a5nz+R4n1y4iZIl7TwLT8uXVWBdOQXjYw2pFkV8y
Y5wM66L5R4OuPmP24/X4ObkwQu4kRiYYQu7Z0tLN5ayjGtbLRTND9Qrn2loKGdEL
E6LKpddg3l/DYhR3Fiqx0B+duB3aRVT0jZDH22DSFRDqnMu6cU1J8fNoCxl04BtG
yZ4/9YKY96b8Nl9TFZkNScmapxTJXgxu4zrDS+NPdRnT7lC82EglOjFFBqt3uMBS
w/Jrek7i0/p7TvlkK1CFiC88H0ZQcbfgPGczFc1WF+tf+kunVsE/3bT1yV1w4Rtn
MHkrIUKQQGXY+Il3CSbh9wPcpMbTSdqx5YXQL1CW0PphHmbly9BhkmD2CcE2e2ux
70vBiotJTy5QUKkYaYSWbqE2WO6bOW6XuTzNdE1iMeArJ9m2hcfLVx+t+uYGzhPE
q7AAsUKQrl97U/iroszw2+F74AMznqZzn9XQ574N8C5cDC/SzjV0tdTGpPZzm6aL
FievnIIuPtCuFNNu+07nHX6f4n0PFASRnMeY7IH+NTuq5BwQyTI6Hv1Td7Mtgr3I
EyoAijsdVwxiPT45zM8n43hmQVXRLTHmbpnYS32LZ7jYUd6/CW4TESbPvxIjBALv
A8VAIwl85q8kQiX0w0pTurDJ7LLRV0+Qa3sKqmyS4NNBbdoG1+SWDmJx/4HuJLQD
PelAJ1CXV9y8slbfyQapl5cOxGTkxLfQLK1hiOcAWGPJK1vcGy7ItsxpNr5ZiI9F
9JinW+/ZShj+ZC/GNlxxiAdE7qtG93Nan+9BVgeZpeeWBvWtn3C9kBmJmiT3cl7j
LxSrXRwUNEBriK/gB7Xj0/41FBxe1jRQOkPx9wFCU0T/eraasc4rxruPOeZVu6hg
pTWEMjI95oqn/ZqMEFVJjcm4c+nOlo0siiRPWa5N1jnRrRMt/bCUFmOos6jLwF9O
eFy+pqgBb4zsIG59fW1OoKcL33nTXizOBC/2lrwmCAlJ5D1Ql5MbmLaZ4v7oeR3x
cL1qq7z7mQFhlenqbw6aaLjMZdTP7eRReiWb/OmQhySmrPdRN8RJhOyFQghToN6d
XNGCSlvLwpnUnVsHYd1EVbqmXP8z89igRukwwo99glJRzhUSLkRne767gu4hJKhF
ovGZ22g9kwVpfMIkbNGc/sYgVTnxCauLkaHcHijXxNcvV0lu+FFXcjPiotwZAZUg
pgcd7b5gJjaklLW95AODl5u93Zk9835hjvQuOu9ZwtR96cvGgW8ZDSAc4Wa06iXu
f2n/AzRez9BlE7ghAteN3Z+xyDrW1VeDh0AkvdgirOhEtprnvHoXicoduZrzCPMk
4ieYF08Rt/MJg7qerg3zL/4kuIM6YjqK5Dw1O6RJFx1R2IS1iNSxQ250Qh0GALA6
wiJwT9yT36HFTWXBG6xR6TpdiszDyYU6nN8S2tQASouyffQYQ3T9NWijfSDyWkVq
s72CpE6V90nMxIB7gzPQQ4Yp/gIJMi7MmJCK2iBc4ZMWLo+9NCNALNWCfmjEIo8u
UYQgsve8BomZgrlMStbDSUYC4y31uwtyWNBoJSCxLtwrZ88bzNw4a6bHj6WCP5nT
bS2xm4tOO1/DxjXCJ05dZmXDb20JnqAh+n76sNk4PRQAWPCZYjbNfVrKiUp2hdNh
wwtiABvJKBWtjQF8XOUAbXX+UQGhj2+9X7b5rvaQ+jCA2arBXWTkXWn+9epfisdW
fHpF0ZgLS175RATaiKRRxH+jaymRbsOY4WJSki3dzgyq51xkGFKpZIk+LjogvZK+
aBuYYIo98Tqw+nzB+McldG9VV8cX8z4UqgevGlJgwMpm+3R2xyZyBeMy0BZXzwEk
RBvHRm2DlnIH6oHQLr3ZEh/DNHLKjDPXHEqiOmLp/doU02oErblts4o5DiS3N1y7
1lBi57h0crLjxzxe1iiGOjcvzCGp7EqWeW38z+H/ltIOXFJNP39LkxVPDKuBpmbv
G59ar+FsvAhJpR7pGFEemFFk/7YkK1mF00Ul8K3NZ50oIht66YlhoLxQNV+yLmNn
llnZpMyCbXTXI/Wet9su/JYlPv0gFjN3O/fC67LGpm5vGApjbiJJh5qqdunm+qGs
dH3gZdD5jQgXpHVBCog/QK9E0zGNzHioVy6PAs8OE2ITIUxJ+ivkkdNCP1FE/kjP
CSxZjiiQOzMEdxgrleJcqxdizvuYWZ2fAq97JNDvFLX2rfPsU3My6/Fex4k0SKOI
W3+N31+G3y4NC8f6Kvso+apwNMQ2MnB1vgcOFXrifFVinckhOJWZBOlYQVO+dZYp
GpB88OtNt1zSQc6v8tSfwLeG7YvCkefzbdlPACk4Z2yXiAFThg0UWdtLZVKRkK7n
hGgcrc6Pf6zn37SjW4MrmCqqVq1MJ84dzvXyvxtxIP2qtV4/7FiT0ChM2JiD78R0
IktRTdWJzMrLtZZ3O5Ec7cWHkZhiLIHMVg/3rKzDDThxqjzUWUE6w0a7whvnR/9C
MmiBnzzU0NpTuILDFu1jDV0c0jKi3IzFUyAFUvQgxeFrXfIhTvGXyaaexFlSDmol
WbPQvKk6o9VDEYXSWmVkdgJp9MDbjJhgVsPcRXAQ0VxRP+R3292pyj0ir50y28GQ
Gal5JJp3FBc3A80ecUhbhpzAkgu92kyfO9rwN8+oiDAMLF1hyQT4W1LRD84+WXdx
TLVksH2Wjcn7DoSwmAE89/37R6OmM10VyreZvoCiM6pKVsWLN3Cgpr/wwizYpGfO
CLJMk+Y9MxkG1UwOxxJPL0QIhWiF+U0tj6ghwGkdCkBYBVAZQWU73TS4+JvNonfF
UeTIltGNV4MoqiqBcE5kAL75cRs3UeKBOkMHXUjDIzoX7ujaiPKUU4MfG1v/Zp/G
kZMR8BY3RXxL3EXnS/3NbK+RMGlpFY0mYLJQRzLaYsPc/PUkxoKWNyntsUV2zK6C
TCof8pw0s6Ibt4aGY/8kJ69R92UqH/NpptvQhjOE6SgPI/ntUkYHc+aMn7keJGQE
8y04iMn7FoUf01AgU/24e6NNylyy/gUmDtGGcTUKpmmH8Sq5mIiqImQLLi15+P5K
m1Ogqbgp0GeUa0TJYEb5PYUzLI01E4LA9D722ww6463jjvvcx62E4zcXus2N5oxm
o1iPj+4/EYq8BnCGlJgnsz50gGWpz2v+iYVwBPpt6xkJGhB5se7We+Ff5CaSYUHw
nZCagVokiu5Q18xip5HeXrAzRj1XZghj4zkfAnTAjCh09YVfGt/IJeBnnf6klyol
6Rvyp/9Tr6GrxlTwRe+DiCvmeZj1yjJ/RTjuCZ0PcKVanweGBrKjZtFTZuNOmEAp
ZWmBW6GQePQ0WbTZ01fhCE0lJ1A5e6+HF99S8SKDF+uBNXQtlvZu1vcJ3sYG8bC2
1ieMaB1MeM0VvFS7OMxEqbPKy04+vZOyT1fnUKqMDJVQszOmXzOgGaqdQe6L2Sd5
1WjaN/gfKalixg2kc6L2rxAXAaNkgbKRKndzYKTMGhHrOY3+25mpPUc64D5NYe0t
HJsTFiq2k8VxDDHEepvIno/5HreZpxX1wLv482sgmpVT+KYS6qGH9EnTL1KGS1mZ
xGtB7sdcme4JDOkDI1nchAZqPOEg0A61n61Jx92zm20znZIZvpqDnITiahyCxOvQ
CXA0jm7C8P5M9eMh+k84r+qlDXqnSg5bQ3dYUMYznlIEVnXnn903JH6VqYaozk1/
lf7qWs+wSuLxhMfo3Cnr3F1OgEQ2hZN+rcSoyZ//AWYQyYSgkuNomGucrxN/6J1p
GfqC3TNziuxkkKG30ieWr3jfexeYz1dW42Jq7Asw5VlTjOsXFndH8npXhPPcmUi1
cl7O0YAw7UzyNnq3DUCN4PoGGbDM+v2yu+3UFAcTKITdmAf2+QCm7a4nibjED78Q
1V9QGsTjmM3QUlJ+Ix88Ot8rmiP1XjzFG43J+E0XiEmC5YXN7Ke0I/IpdBmUdQnd
l7pf56SpRm/uejsF+Tx5LUvw7ml/TGV5iNdoI3dPWs0TP0w31Pz+Z2zkahrIJVlX
bu3ofT/SOUCPaVRmctfPaSd4QFnn487fmvdnRx6S10FQn9nMwHcMhs6CJ3DmAArP
IhLHejTmyULoX+2fpF8mLffqqWruD8QSPrG4W3CUmNoVQkWdwCUHz5cOUeHDfODG
ybJxNQ4phqER5jIksYZAF78cTO/wwjvM0YWqRW6IIEjZ1EWdvEmupob+JpDAEipM
svyABfSi2kZNmdH/lKEIT57KysTIgaKrjdCEkGv6VC3NHP7/TgctJ0l8VDCIpJ/G
fOFRBVv49cHc20ltJMN0wZIHZV4/rZgCnXtzFGyf6Tr6amNHpp5xZqDPaGOWNQzV
OgOqx8GPLRzpiWcWTOwwHlJpVjA9VbZ0N+swt2owN4WZcrk1r2DX/wKiwluFp5kE
XDw3nIb8ezNgKvo3mWOOb3dKMqXqRGnnMISq6bFB3DwE0rSkG6Q7rAshhDV9lQ/l
bUclgV46lqerLy0ttuQIa4ZYUycIDn1e3c9A2mUyd2m8M6jltB6HpO1aDRd2IOYK
J6McL2FKDhwOAw0P+F2YRu4WZfgeNx4PCcnetpTW4bvX9KpTMda6Q6jYjTcQxfh3
eKNQrj93SG0SWv7D7Q97ViKG4lkVVl+tx7oLuKkXHk40SnauXnChgzAPlX8YLSYX
div3jUQs2Ev+lafIMmY7G53k0UipKP0nZM/KSP1XwsHnsBA4dM1QL+w9N2VofpVe
4EncM48hz5C5z8oYgkruqYxFhoGYiW3Ga/liMQ6gtb5mwAkBemiRRe1OVIPQV8Jx
RfXnUBWVIsb3NOaSZISeqEv17eTHm5jnvbQb1LwOQgNiuT8pYh+PEc3D9ny4wnYE
hCT5lJrq74OdFVK6Z9pahhQ9Sry4t7raws7TYOnHS937LkgiFaGWVtCsUOI1Cn5D
33N5G8z4Qo/1eg3Qx1VgR7xJY6SEIEOZKgrx+4knDqQeCvYYrr9lCda7I8faii1n
mnhWihhQbld74KKkYL8CEycpH+JoDZvF1GUsTt3Fzi9CuW21uPN+qspVIt5HJU1a
M5OEBVeT46qlh5K2Dp4auUIitSUJXPHk2gAkn6EIE/ZN9h2NOScuAEASedVktzkg
B5C0xf/khAYhpGSxW3rpb1ZarSlwsNjvLC0IERlXWpqQIO78ununHwJhbA/x+zA7
QGjfyvD18bWq3ooYmGPp7C/WRTuq77yCO7lzq8qC8wr+YOwnVokLdrvAV7V3I+b6
FikZtolp4CsRZhDj3lc0str9h/WI/1ib7bZ1IMrHEywr3ry7uj2/VS97DTwjMRvy
Ea208VxdYgkcwQc+Z8KhRi4HBY91WiBo/zlrjz94pJrZ5l9vpxBu2x25pvJP1IQm
lmBatmT+MNNcnRmRtSjOLEYHox4ZlPKYFKVl8zEPPQuNPAmCIo4SVlM+CnlDltjN
F0Q3ILWfOBeD0oyw332YOCWNOU7yB7lbNNqYz9oM4P5oQWKYu2U4YnVDE5SjPhMC
iVIeKYB5k47p5SkoQTsYQQAcFJ8+FKobRmbrh8WpbhZmK3fQmrY6TcDoBaQq9VyZ
NlZ+B/4mHeGay8xEzHApGu1uL3Q6CTk3bIx92wyng27uLnmbxLuWXS5bg5NsrkAD
04AAeBW01eqAOzYwSSeTJGh7jvjKmaYLIgW6PU9b03CxmoqpkHiNCpKZSAUxrRor
Lbj0XhsZ04I/x+dAX+Ff8GMeHwZpOHSsIo3Ajt9q2Y/j5p/rW1FKy6Q86Z8B59Hn
mk+VHqokaOmPf5JKpdzCAn/CyY5gYo1jDBr4WuIrGoP1Xu5jojdAfo3Srf1xSqXL
eXCvTpzjQP1TPGM5EJOA6BJ6QhewkF6p81Nujp/+Y25HVnOCzA751rwThzJBMcdc
Bu8R2HQL70Aw/zoI2tAKFLkyxXXJIdaw7IguylNnMV3EfloTn+aUROZPqa1urxsL
UjENi4Qqo7XcXhTP4FkVWrd7iplYSXEVfiSMrVv3Rl4Mv/xc41DTKO/UIf/hIGFw
lKHF8VRXVqUaOtfwKNTLfkXxF2jy487K6KJGlYj96FEDhyxxWM9wIGdxSuZAXC3M
kL6BiWbkW5r/2WkfgB6K+p8iuhn1/zS/Ym5edMyacjttVNYs8o6pAL3JpM0n1Qdu
bf2pXtBCpgWQwSaDPmMDLiKoOockaSQqKrrLWCFec1047ZztcLTvIv1jf3YFeKe2
LB4H61KNSxCSQbykjxdI96CuDR9aJB2+0Si7MwOaM4Md7ydQSmRArxbSdkOX6qA0
Bezx28wl8nf6WxjtjwyP0ZdO6Uk0GvNmEgS3SqIt4YqOrka4AAmBMI1FHE/Gr/YB
6OM/dlmWAF3WMIlVUh//rTy81j8YdiBRyWj1Ho54jclyIzP1V0iDMEq+FhieCdVO
98Ra1/n1w7uLxNgXSSQzw9FFsJD0Y+ZVotqMTAAenvaoZ9t5QpFMGNSdwfpHjDOg
THhwxeGdfiRXp5XklUSDx/Nl8C6QepI1gfxYJnSz3x0k3SbTZfuf5nhwfxFn7p98
SatCqgHvBGoRSZecoSyPV2LDu5RnFJR70pLDS3wrkI4bVdYWcQ5lLUlwS4EKdX5r
aN0Tp9Mo0pQx3BHgt8IVPCfVbesHXe0CeaeO+8/EN6IV6HZd34u+hflUTSgNgBLn
vRqoEeoafdz8qPTXTlJo542nmA3fmsPYQZvgs8YSWhZCAphRlHv8YCC4GJ0/xzbw
Jb3B15RfcJpo//Nsx48s957JffyztJOjAuHgiPUG1+7xm8xcU8ysmlIUyZPcoUFl
J8boKnbgVBBnjvepJyP9uvHV1fK1K73GB4fbk2pNaHJSGWkyPRlO0JsLAz2qcyl7
4pwmFU+0zRXF2lwVxcUmf8spwklhfoiv9Ie6Z1TA5z55636nkKwc05dFhWBxHhQ1
p8ABKQSbofDH3BZZFuH/wppt1zA6FnoCIEVNLMuqk8O0qEeAbCTfby5wP987mwOf
XxN1oP/J5SREoX8UQq+6dm0sq2E1y31fvr/9aktep3DclN4vLAFl89ESGedgw44y
RwXVICkul0QMzMe10r12f0K/uax5+ZUkU3CRLNMybTssqmdyF6bzGFJqqdiLcFJY
UytqtmLaBfVbmGgNip5kA+x6bpa9f9TGf8iIz3BucPvxfqZKjsWieC1YhgK2dtzW
t4XobCVIapwW5IURxgNAXNsS/3mwysfrQDRcR2A37aQUExIM+oKvqQM6TQ2gdRQ4
Xt0kQa8vBjg3HhraMCmAPmbqQMBZPK/zT5eZ4eMhmchXi7k2qQTT5hwQgek44VPK
LQh6djRAcmqB52x/UCNQ/qbg2ZwKSNLQYEkCPgWdSkE11PxcLenrRzUDjsj/dm8T
XEkJdSoODUsXtSEP7b3njUYmG8G8LTFh7GcV+uyJ34frUjG0PNWhBcTu+457fgdF
poPoYKYRUXHao8bHFBsTHSIlpIVkq3HzmsVsVk9xTBjmlXUF9fHSCLg8aCzIvh8X
TuwESM6poCxbh0cy/7F9VTxaSZ7SD5q4zulHhVXNJdMfHD6hkcfNq5uXQ9fVA2fe
xI0Zg9oH2hdZrpvS5eZOChdOMZlq2UsGRLrdA+qGfg5W56CEry25wf5cIMuHN34w
v17GI0wLA4SZrW2YevamZILhlXYXpe3xg3JoOyd2kXGItKLB8pa4XkDNEi+WpLpy
qiRMRM+mhE+q+jqfs9rt3OPZ8GhVTGRftF8LJ9A6SY4xGpY2OVgiuKJBPCtVULJj
D/9WGAbNfeH5ed2NSSWXrh/QSxuhbxte1S4fKvcfPqNMfGY7ynr+IGPjMMgD3RyC
VR9WREpo5VkN/8iFOHSy103RvEUlUtmbIpFvd1jRTrglv6zFXFA/BCIADNYsE/ti
VuzlzTIjweIhNCHwSSj1YFz2ZAuqLmdv2g/tYwT98ZEcScofYo2W5oHuca3dM6KG
AEzIlkHSlFpE5xHPq3SN4dbvOj9R7uA83YXNXepca6JPbF05d4b84Sg9q64WTYpM
usuhOWRpPZVjHxuZ4yN5EHSIjqxCS47GFWCBgWnlxiT2F3hIfZF0J0q32qhn8XBj
2KsB33sZTPPD4HGa7wiBM2+CWFCH975peZEU2m8Vx4y06cz1x4JCRt3Gnh3L8R8G
yoEHlmwZEklwO9qBo4zKpyoOAVqENKHYWuaNe6Ax1w4y5QxZVfMBlU6+MpIjNgzC
0m11vc8Km0sDY6O+SWobfzvdtDrEeyReNt8DJzohzw5oMkCivK934G2/O9d+SWTh
eyH4ravxsO90TIUCyRZ591+oig9FMm4T89cCFjFjW+jJ7IHJtFmcFomoItqzLnyw
T9dCLF49gror8HuyMKY3s/lmROcMdTAbZu0mrCDq8IL/oWSvz0KKZ+CF9YB1XgpL
Xt0EUCUosNEZJAeHqiOZBQFu8aKKBjzWcJT61NSm7ZhcqHRM1mHYtFtLhUZzKT1K
qj/y9M5pxXUMVn3+rM+ettUAUqhDbQIZgixyEAghFa1viIjH8Bqe1pRxvmgKLs2b
ld7CTHpSI+Mw68jMAid8m5n7kTirIAZ2JeyN05Uv7IeaqyEuT75wYSsgVWLlRRJ9
ihX1EcXvVWPJVOz142HuIoulM/t4NX+71YUIHzaEpxSrxEV2MU7jE6NRwE8TrYxa
sDwpYEjRzibv110DPkJMxWBtBKqBtoj4gPipyOJM6g8k234hzPNpVak+cMj2/X1X
3SC8bQ1Q/xSUiCpAayMyXEDFVsKVODeB5yev5P8ZAy86Jnzno4e45XOxiNRElLJx
Pr4tshhMMvREUGS49eXwBhoHU+aWAD0BJdW+rkPiX0uij1O0td7o2ESd8eoj3ZZY
TIWFZMr7OjWNgFNGLgUUoFLMCKpu5lXuR5Lg9RGWebmZv5LnrxGs/8goP99Rdaj+
4YeNaZGI3mXERLH16BAKYwa4tzM+VhBMIaqQ6ggZyvmW6n08407KI9GsChBAOcZo
FcxcA0vxLGlzDE6aSWkXZTbbC3uPdiPpflPx8Vl48F67VZSB54kiiTRjusf/I0BA
aIO26oUdQbCT+JdAeHPrCZu+ZeBdKMa4IfwCj0OKv2to5EXkVFMfyydynlsGoGFX
SlGMNyUQ2ocgVKZnjUCvKJXmllNYeeXT/M/qGJguwx6dTrZ92AnKsWJpKNddqpcX
u7jM+h+sYTEfTk3Ntdj3VudNYYHC7VudViF4w4XwS2Ww2xZuPm3tdrH3d44bOePa
NotbPQ8C1ixIR3Mpl7wUFG4vhkOGUjt98TJGwWYftnbChuuNwQKNimKLCTf3i7O1
QkiWQcoUuUQeSPcyz+Ic3pu6/hrNlr3rVZ5yB0w6wXOpOmIai3rhYVv2eFAZ0b16
n/avFBomZjkkKkUTneVfy0uDtSdF8zwUyoazkLJYihFMXkBm44D5lnAGGKHC85/r
GE+H05d7K+QwBiM+wRIp8eHALNifgpbiXH7QWdnz/KxNnozXuOJ2YFm67dy1ubko
R0KrGVV3CkBGjc3uZ9Wbsp/seaBJIqKElBSj1GY6lkE1cIigveYtb5wVG+zQjZx5
G+L5qPZSUmX4fv5A04g6g9GqnH8Ub48PM4o/wQjcJgL6XGAyH2GBls/NVz89w97r
L939ls0NNpQUAkddZjrR58dNIW1uWEBObhkUip/mWN/rJEMM/H9C+R+VnBQlLf49
4sLcBNinpWmT73iWih6yAGyiIB/KsQSjqs3uq72tBJ+FRMhpmYlLfMHPdKMreDr1
CkhzB0qyZyGTUjEXUjYGxcHHSbkNyXjkyglHz3RmLqEyOCJQmz9xwxrRb2cYzcje
PApZvLL9sjXTrd9gvgGF0DcI/Sukdb4+LGylZrRbpE9Guen+sRdd2EPX60jGJXbV
IjJOrscwH8LI/wIZSWosrgEoP+zORvQboxxM+h4AP7z3IZX92XEO3sQwnPG//k9R
n5igXfmmPa8drA9p2NV4jZrRAv0Rgro8PXdHR3vl+g7orLod+38sjO8YhG9tQrL5
PqDPGzZrTdax7hOo4tjeF4hdAYPt7r622AffR7mRwuhsVH9tnQlHgbBuWf5dYrFW
fza73GB45Lu9IifocWUvV+0fxG73knu45pxVQXwMTzegGgH0ALidodiUfSyOIwAw
7/oLY2XZN9zSaIQD+LH5dcOjDxDsb7w7iCmjjUIuAUjWvN3d1uwxcr8opn1dbPS8
AOUu3nfAnZMp13xl6aL2xbheFHaoeQQvJSWznki9MOiCQFC4WGzDWyFl5srYmSTN
UufGwVK/7pRJiJFN3zvUe9PNF9xahqahGMqKHpCcoy8kwuIInQzPqbkum81j1dGW
k/RP2rROGlGb8avbnm/kcr0pJkWatELNn0xPqn12B5Xas6Fo8N0XAIk/vPpshEYk
+5LXFWGXeuziLWv5+tgY+KsHGvzGnbWa5E7q514VWylTBLbSIAqoe0l6gA2Hgj/f
DsOJ+teNYaau1j1KXimREPCcIZKMGApCygw4OKYkFDsBxAFHW8ikGmgwBGCO9FPb
CAMZzsqT2pTuh2WbwU7CkRJIfQpPnz4zm6sa1KlUuccNZnh214j1vBsHp9gK9w7V
qwpdeFG7NS4X/1OU+mi+IjuxvRnqPm9nGuZ6lpPvUuzKcDsOWv2Lhd7r1oBgIkYD
ZC0aFJZgxqr+aB+0Arm7ePsk302rQ6ILyzDJs+TuUuHHpfyRv8WEBssmF+FUqXdU
qgkSaUMvR/EalDNYLFci4wVaj4YsU6yf/OZ+XvblmiRjGky9ffMq2366qfo6O33N
RLqkRMYBJ4eF8lxmL2AAUV6cFpJuazGXuQjYAThC/tm1gHhuc+tyNoV9JbRUSbPH
l2uhQdWz0xeq1cIDGWhibjIfFUQZmuEfg6Z9h/MTmqqyF2TB5v0AfHuyzuw3weW/
zvrYXDSuO7AWgeBhNwapMQbjzpjVvwVv3YL0oDil7+N1HYmyOZ40Y9hY+mDMGevb
DGT0NFY3/AS1I0M7zhFV221Hy92Lk8OAvI1N9exyUybXOGn1n4I0VgyqsRVLUYGI
TlUOZTknTuquWVoOLjsrjCyrccWaYpupEpQ2Cc5QToHsAGWYsVgt6aWNlQaLuTbq
ou3P+RZ7IrgKhK+ai/quMUa8OgmBWRc7Kx3cZ2QuLAeacLg43wV9nlrnNpdmWxTb
WlnSESsSNUaCNuMKXU4xN+oiWYhnBPRcZ2VRMDrLa4R1fG43paW1i9tmFxZVOWLL
gc62sU+Isadmgnrt/iJ/vWfnP8GG7jStVVkx9T+cnH+V8oQY5zkU346Uv7mGZV1N
/05qoXHKGqECKQ+QAr+nf5VXVvnmmx1+WVwfvJr+YhAuD7oDWnofFA0gNkSKx0fq
qdSO/0N3kVHGXXeGaIVAdKSZizFocxdOEKd8PN7SeOEWU54qtIqkKMn5erYKT59c
IXOtJUUi1NedcJnANXuAYfuQhoJ4ZjfCwU7tk/aWP6oZjQEM+k9oqEVULRXqZ3l7
3wros3HWy0ZSH7cJrE1DI84XVGhcU734AsJ58tOGUsXxlqj+n1k2TXYd3UbkONgl
N2ktAODOCwimC0Ws/aM3FKrvMyLMDSxpcK3KkaEVDT6366aLO7gkzjQHhgNVbfL1
noUu2X+F9Y27qe5HipafLG1Vv79go7mN4hCQDbARxU1EoCCM57rGsCsFY84/gUG5
jqWKhrcszfgTa13koNC7Hux3wdyFW2fwScxc/8Ojz8QB8tad6jbCcTUFkE3MTF+Q
5VX13Z6Jwj/hEQM1zGjODyZRZ514iuVuGj/EPhHV2tkYhWMo4rF1+NxyTYNO6l4n
VDDU36jKnmxgKgTyI79hvrlO/LGxlhDClZsGQkt4q67heM64NjzIInXKFtYZdS5j
gOOgWFC+gi8rgnPR93xP140K/q+erM+Gu//vw4/i1okw3D546gPXSrHw7jEsvxX2
W0sMeJ25hjIeA4GrhLpXCk9yV423AoYEG7wxLLzhm0QIBJrJ74jCBiDZa5oihPZt
cxbJ5uQz32rcuIOpBovzhFjIgE8IhEQtiB5wKtVHk+gFFOzsNSXsGgiboWbUbw9N
NuWHZl3asFn/BGEHkBJqNewHUHPQ+yYPXyDr5broZN2I+DWRGR2w98+zVXZXer6E
M6wEhZ49ceC9nkORgCfVkGj5rQTVnEHhx3ABVIAeQhW4ABhHAHf3V1u4N0VivA2/
gIiID89xqbzx3XyIVl51xcUXmXb1w8vRAWJhz97cnVUxAyN6zLxNqwaPX+2IrDrH
H1RvBX1Vu2si6yzqGr8SiVssKlFMYaxg/VxymQjeNxq7m2pl5RoyvqX3vFX5V+uj
gJ4ygF2saH50F3ZmDGO2I2w4imMnqn5pgRiiyxSJ3KV+Q47Iljk8AFaqpK1W9Hsb
5pOnk/YPIVJhnhSul/zefUVHhcghLJdfd+uwiz9OXPVTx+dTp2Onw78ehTf8g5qi
PwzEGONa6cg2co37DidERlJHLMpBtNEUnyryv5oyna5s7ySY8tszfloAWjbeUwnt
p5NDOBmgsoFKfnlg4PETPOUCV5khcG0XACwt/7UzGY5uv6OJfhH6RlDlKmWAQpmU
w1k+6l6KtAdrJzurcvIa+goJaBThIoY/3GXxBTmWj9hUOX0v7qDZLOpspsyScdle
qWGrInl2ek6GDErj3TRwphy6ZPTS2XxdjIqsopO9tJDVP3vjFLVnohF0SsPglns2
uY2QDQ7izO9Lx48GtlYjexpPXCVhzE7YrqnO2/+DFJkEPJlYitUzW7EVFAfYrGRk
fhrUczxKemwBtPxH6iZ0EnS1j1RwV+QWAbwak5Ygbdl2hy7OV+NmeYNHGDXNId54
AyflSzkhuYLFPqg6TQU75F11jI/9oja8XfZHo5GXQCXjZAgwAg0jzr0GKymHGvNg
8aCwvc9vvFPUg0w8G54MXmBW4AcNPa/t5tPemQ1FJTF2g/2uCx1EzNs8yN9Ss0Y8
5dM027qSsDgMTzxy1OFknWvBvXwXOZ0otTKTJg2Q2zcAG9sKWmO79V5Rst9DStm1
jZyk5gDCr1E4ltQ3lE8sDM4TVtyZeFPbfMHVfc5xpBRB7WUKR3G5RVErR/cmDPWY
n+aB/ArT9eToVOx3mpzTwRs3Bn2Tdn2gaouX/Ybwk8KNhYuANi/T/jyvbZ5U8baS
qPBqD9i2o1p4rdYBbICMORmniBzAIvPG1JobBGVRwk2B9UhYDL6hv3ElZWB38a3u
tPrSbf0EPcKlzXpl0dxa6XatLp5ShYw2n+RWbp5E2FFHQANk+L4Jo5njSb2jHyV4
b/epUvkluotK3ik9JnjkU6azHe6WLnczx995JeaULVXUVUy1Uqpau/1pT7u0dLs5
S1GNA9eNBKUSOmY/S4VDIKxmIe9chagBlNsN5ys9ehtjFnutbCqCPjrJYhvfayG0
OGTP9505vomHk31Wyolq7K6Pipo3fxP9VogLhyXTIsFUrY+XjYng5ucvicTqhVCb
XUuyiE7Ry69/vmZ16inRmSwI2/oSxqAr75SnxM3hyMjKd0pFSmHH9axoOg8G0A0V
nY1YrycXIdOZEdt9K6t9N02wlvXUAIj391BYUXVw7NvJqBRw6NjZz6bgqWUoBGxd
jt+wNfCqFTzVV9HFqjCGbZnwunL2jLq/ZjKpUq6JmHJl5i3v+zmC3Kv2Co3TwyEr
iTjOctMRmjEQvXoi39YQ5zZlGvjJDXZlK90Jfd7vQasi03XrFC+J5beHuf6sqL1P
S8X15cLUk+Pnzo3DWwb4U7HdNAFI2V1vpdIkaxT09cygvCN991T/CWMWM0CKb4Ap
i0F3ZqiOxWxP1XTv7b8O77Zy2KeQKcllwT3BWMYiLMjdrINNN3tcqouKdzi1E1NA
PjAbcsgy2gecKs/MczAOcvj9CzuZJUBfIVyWILPkoop7qpHmy2UDsguUjFU4osUQ
MLga+HVmSpju9uaKo7XT4SJ1aXEzHnaTf9Xwp0DNQ5qkOQg6FpxFBafx4f+4eJ/p
fPhj9qVsrKHOmDeUb1Tm45iF3Mdd7cFcsQpURQk5ntOKgrKbvK2NvS+O8SB382ru
u/AXZkMMnk7W1WuBXEePwvxVzHjuT9WbIf7JWV0ASaRRFd29vBMA9yYqr2zQZDQ2
jb1BT9Y00E0IV/XIlLtnwsup+nA48NY7gR+Om7iPsOObq5iIjrhfiEeu9hZcWyq9
NfKmuiWkziKfyHmFVWAkGoV0EXVyyUcJ4HDFSlmwmnAcOMPB4Vw4sZjimBCzlK3F
cwVZnsR1X0j2gqeOsKHUNcEXQVhoXM6J9z+JqGa+8IEjfqa5jM3J5INhoono0Fz5
DGmL2KcaZ0920tyBw9SJF4+7TM5WLDQGTlCrFO/j0D1INBuPlfRgoUkjuLkv2+EG
ik0gzXVptA8UmPby0xakX+5VX6G4H3DUN3v+DzeNwOt58dCbN1YaQHIkfuW0lARN
ZjANzd0xBcMLj0Aix9AQPDpw13NKssJbF0RAa0cZJEX6/qC8csVBMih3UNjUre/e
gsj3jIbte7+H85eGxL9Je4A/xSQwoNN3lHk3rGFX8ytJhCe9BrMaYpcH15LDFo1A
+VXYZTBxPmdc7cB8cB2O4Qyapy6ID0QRtBs+0vSvIgPzTrPyUsdLYEPTMc2fOIVQ
tPnXkgf+P7KXlqAmEjXZDu5N1pLRpY7dhrGUGv5UIwierBWSGkN9CyGx4LFanNlK
+NrIWmLn7otdQDP9KbvhkeGoyWDbm1Nk20R/SC27LhnG2VU5Jyo2UKHVwYH6mGDN
izPRkbk5uifareoQRyaAMu5QpNZHG83JP+nuHithzoJQ9sO0ofeTC7jss9QugYa6
+X4SwZ9rRQU8rq04OORJwA/O6G/gSkIIb4xq7UllM8Glkwx7K4W9SkL3sGTQw6gk
9QckwH0wKmOZ5juXDM6HG4dADuiCGILjCAGhbKLCbQwFu6rhD7AswrmPQgKKNJM5
S+pOggFpHuv/wEai+BzuKbL0L1W75pWu0EU6PZMJLwl/sspGD1oBo8hltBFmMdGY
nPb75F9WGKQPGCIBg4H0OWDc5mUUFcGbAEYkkgobewNfdHW5lvAM7S0hGwqeMeWi
x04T/2ftejUmRaaDXFogyiteLBsiPK6CYnIswZwdGkzwg5KziAz9VaBfKr0G/Zrt
f9GsUx7cOioL/mvt1n1u0pNu/7V4dSj4adHMnwVAc+yGQbdKnW0qOVtgC9BvjgF3
9qEqoWyzFUoTnKwtxHv9XmXHN9bcv0e1+9J4OnxUE023xYsymxJZK1av6khGN9zw
W+EpzIkmnVrdjArmZK17ToCxIXqOuUg7CCiDMIUJjGDyeyR3XCMEYH5XhlT4ZLAX
0EjvFIu2t51oTSNJgjY6gtdEcTIBdls3ANkbyNRhFK+GvdgwkK+on13HxgQZLdwz
gny0cZS+TEBm3C6C6zTldeGJ72iSRURsB3LFWJBwzEu65eCc56EPLT8udDvoxGMC
yCK0v/gSni1d16Ehk+GJ9DTzLygvZ999f8qK6imjpMF9t11ieak1DN7vpo0HEn0C
LpP/HD8RHFBVEf+jBjB3+Z0nD7WRuCHHJYvmZ36ODMYDavHdAIQVmG2Q9duUBrds
fFaCORmY2jJsKleXgSSilF0VpSqdVtDDtHe6L4rIDZciCFynuxGz6zvQXWc22CsO
c71zCAlPKbFUwsYbR6FqSAx48uQyPMm1hdENB91chNCJdGmy5L6HK1Dv3pLojtQq
PB9fDYHlLmR0MseSGpdFvgIDeWmbnbmGsThVCoKpkP6hujlEbiSbPJ3F0DJPP/7S
k8I8hPgpxJe1qQ6Nn4irikqT8eULomQRal0rMC1OjP3rzqLFssBuD7TF/ibXr4Gg
txyPlbpiRBfniwjkNrUVH5FGvQfR3G12/P9FRw5kc3Vi4rL9LomK44fJXXqh4Nnm
6AlbRjtEIbq7bEqbSHeZQuzW+F97JEYtXO7ibwTQvLitipcE1DsxUp0V+O75eGe/
evMaWF71WeMDC2qgd24C0xr03/wvatIhRbD956dMaeoS2/Fln2Sc/afPgnyjKb5R
nJs6G2XIhLOSU/mfJsXmng/yJ3c4x52qUJeLgeScDT2kPKgGKyB5acrK4Dt+Q5WF
kyvjwzcyy5+pzhphnsTNvl63K41jCeZhS0MvLrb0lqAAOFGux7VUm9vJOuEWUhuD
JHoxy3HbZ8nAH7YVWtIBaWueZFCf9UZh14W8rpCxLdEQWdcZmIwcnR4XJ2VpSXJx
v67S82KwTEkNq6i7hh9pemHS6Pb3aPnmPB1UcF6kjrcuHtAc+SSElzHg9b9CXbxT
VmL2HoDRz5erd8dN+t4plbq1xov34bw/alVtgFmdBkguBWkgDfMxp1nmZhkC3VCJ
RkrRY6pOEQWR6p4jLcFUn/JXifd/L6ctvxes7nluwiBjrRk0xuTpeC8jdvYuLKWo
qmOs8G1jdZ38j3j0g7EHWnAAW34hnd7q0F6MPr+R0Gix03xLzce0tYWmk2NB6uFA
DeKBJvJnBZ1a0OtwbSMvHwLOzvJ48YQ7yWy6dVdaJW/GjtAqPvJhU6pmOsuaeMnF
u1L8nn0Jrd/7VMtJxwVFDfi/H0H0tvHP+zJfc2AAc3fH3A7jmSVvptfB0OL+r6Es
MG411sEU0QAVt3ZpP8E6I2w4/1u3la6OSQxN+6Ji5ZA+Sqk/99oXfsHhCbhRix3V
OGsd8ey1bcOqqPnFR/saMGnC9lT+Wo7wRJjxb5na3KumNzz93B8hVSBeA+YDQlwa
Zs9n1/uHMIRf5x8WZwiReTOSyTiF+MePXVyF2OdQQnTuCZjnlcisXariENpnla5L
mtnbmaQNGfTan6sKN5nUTKGDCSGKX1jkEjf92MQI6mW2+BDvGqcUT8NailLRBndc
OYza933lDzfGa5zrD8meUNLHYGg/ZD7iJUJYfx/GqufwiK+IWNy5nyl4tdXzGrjl
eOuVJkQOWoY9o1XiEz9ZPM0IrVOBxyhsZjwoHPPqhnC6BCg/qub4iza4AhnNwW5W
7DXOPZ3moivm/6x1BsSwy4wfptSmHe4Jm8dtwIgvK0WVRpypaooojXhuSLcLtRP4
e8CgnfuyQBLe7bPMrQIXVteeK3ZGh3lj8dFNStmhSc06EI0/dMWIb7vKNW2WBG7u
PFRjRr/euSlYNlmwYvHURHLD0bkCzex1uds29baMyTZe50VXmjpRkA7DfZCMP8MR
q0XnmbZps6cDTQgDm/giMFkGzNDoNLfkbGLJeiCUJGjhnePyQbcl8in1dcaU/tdC
20EiEUQWolU8/LYYd5DMKJKEV3yEon1JPubNaKdnMJu34/ynOGrse3HoxgEtozhE
J+ic4K11qkCxLwOjAHt1hdEIV5FCbX6Z40ugdVB0VnSrJM8+wOkj37jRyfMuCkPo
K3gYA13Bvy7XbQqxsVZhG04ajvaLgNJw2WypRcK6CAZfeP8EtXC2mz8nOYhHYP2/
yTHZCyMkQFdkIJZWIfOYJkzCEVvlBEPr3UONoT0oBLXOvURq4qBRue+PqSz4ynyD
TA+AWKXg2rp9SA2rJsjd8iTaIoPCJHr1OLXwszjFT8A5ig3TXe23QgOHASsjQ1cj
kdtIRr3RHnAFPFUwk9Fh3wqBOh7TBG1lLe7aIpImjSuDMUGfmtf93ofolDLpzQQ3
d+1Ksdvaq3a7QuwoQS+hUBRTObuItWPYS3EdbiMeoTXkIsCYHoie7w8z87d/GUgB
a+gyWWW3KR3ztjNoyFMCobZvJZIJhFVe3EUqeMcriVx9jPXO1knpk5WmiyAy6vpk
AnYrxC05RJGQ34xXZVA22be/A/bh5nD/w6SWHAzl2SEpsvRnbt8W6i+okA6R8jPE
ysed0Y1rJCrFs9FfnR5nZKMYrd3zRaKpzWMc0A72hMDqsxpnhBWgc/O4g8Aik+kc
99Vo4AbWeNS9qOy7jkbmgkK5T2yYTMUKzy8awFmsPAhP8KRACgQRZnlUXrOLPV6R
n0e7sGfDYyBxRG57QvqoceycPLdfkPqumz9St8FrT6fBKyCHxu1Mq+4ZDC/n0sYX
f6polAgLwXGQzZNBtNR3ZPyiIamwNV6OaEG4BAJJE16gla7wPDzzf/wOy010vcON
bTMXWafkJXcHfShjdYyEguoyP7bHBY2CfgNrLxpfVkGtKt2/2HdmxMuWjaw6FZpw
s8Cxk4hbBeLotiFI165HgWdpsAnLTswTvaTFXOHijlkKVakfKyT4ZWLpVu/5yXxy
A8yIx4LihFLrbhy1L/UJqicuR8+NBMJFcFrXHc7TZyPwKCPW7yqmrwCKZMfyVu78
rEg74OP3sWUzBQsFdfg9YJyOujAm1J4t56+zFetjM7xFDSAQNfhbzFsXjIHf69ZL
NHyhr0SZjG9vGTM1Zjw+lO4mL1rQzSgVxxVjXeKBG5dm704IxwzaiPH7cb6VYACl
1l3ONOlgj4zz7ECK94bPZ2AbDMu18IA0345l13GHLidQKB5tK3KOeI3UWsE6viUh
/WHZnpo6Nh9Z1O/8q/XipE2ssM/MlVpqbGXJ3osV43L5pu524u2Onmk7vUlgkwbr
j8mTkTzDHQ4jeML4qWeLvc0V619nSif/ZsbrMU2sNFip0toPkccnAB7GBPCoq5bN
rVVp8hqFNM2azd6vhWnbrbzQ5uMBojioUw/enDspra57w2UcItnGo17lr22bNmmr
tOxRlm32EP/38PsTUkmHPs6bXvFKHbAQ1Gyi17IE7Vmcf6V3cUDj9eMltMXzRCfU
SzxKRuPoL58lnQEiphkeFx3wxpTRE71IKwWXrfMAcTD2m6WOt0SYuXmZrLA1adI3
N3R1rYTNNXpcYjO9n4WJ3ww2z8CcnHGFTHCSau+as6XC/dcHIE4EqUDbJ2ff2V7Q
ySlUz9GygzARvyRQs8bOk0+1ISom6eOVXdiPtBPoNSf1830sWvyCgeGaBkH3krjd
fWu9OfJcHKwLqstDQ6+06FbhfyL7YTwvaOmvZAF7vy2IWct7vjkYNtSrXeXQ0HiH
A+lOOUWSguMoPE1D4DbYSETkAT6zkDyq1aiMWQVfv/O+TYIw7+IzNRG6QnL/1sEA
WXw+pWbFBRK2FBehiKB2XJjxqlv6btfwxPtftEeULlGagYyEHN412FJzpPtDziOV
JJsQgHu6ZIjQEDEFBw6ZQWfMcLZlkyKE5rIo4fmPWhVheKwr9CkOgKBKBzuAhv/l
gIFACfrEtN+yj+cYKLiFX6G/nlJcsh3g/ylY1C79AKA21wms3UV5DOTGKquGLNAt
K4oYpKkO/gDNfKn5DgIzuym+8woF23RkIo4yClGRuAnrd0WoF18aF9rvSxPDUpH9
vk/uD97VxbwTZc8mh9XBgyAdLSP9BqY4HmYK+33ZZOPpfbo1xWId2AOECtC2wiX+
dkbrp8KYh2UitIBZMVn/JkLl+5k4FThyNC70jtzU+2geUIajnXQCk8sQNwClu/Ej
Yk+DeTaYfIHoK/3i/T87ittvgVIv4Fs496BowMkwGg5RZMX5hIawCJdSR0qoXer/
q24J513HTuECsSlxY5+xRDofrqtIa9fWbpW/ImyNZbLfeugff062aPOw9ggJxIBy
IGhyv0HjQeFaKG7BFgyCpud3CGSRGiCLYIiCbCH+UI0K2Esh33muDW9Td9t4UMQk
5H7zNfrAC4DKVcW/w0hHo1PCFJ+97FIkX3mYuqzAAAd3UXJfH5N3EFwIK5h9JslV
+XQG16J//wrxi8UfYkW4i9PThEfO/LHekBIqJL9Yrt6eWa/pelb87BfMR0zS7X6u
58JvuQ4aMGIZFkCkvDVGBXZKORZDQXTKtSCEK+VzWdpkXPM7VrL+CEw7te9PP8Mc
iR9qRBJNyBbZZj3IT2EhR2g33muwpfe8lA9a9D1UhOx9u1OeWwCG6LtJ5ppNmijz
AdyFVRxJ0nQLttiW1oEPDkWskXOgQcDZGFO2fI4qCScPdgvjbK15OHCAThpxbR3K
CTz6zngFVmk3YwKV1anpA5DkAm1pZhxELD6eRaeUbMvtWyZLgn29+33HgJVVyowQ
GgANfkIfRR+zEnA0QEoxCnF1p/nuAZWF3VWNbUkw8xJ/Vjo+edXIKheG7xJgUF3c
Lyu35bBkOXDB1N1QDLlJDBgfuKyfYfTiWGLv91qvuivCzzWFpbBz1PicvQh5RBQb
Jz/8U3rhHNAzsVw7JsIgw9mGQep4mzneGA5VoM+5GVmxRK3xbktVUyUuE2Q1fs1n
X+bHi31960Vs+yLoGKMuiLulj+GMicEx5WRXd6Ge9YXlg5uY3desx/xDe9bUApUL
PwKOm9yUTKWcbvSM3CXPis7WPNJYwd7Xus83X5m8KUc/4+iCZu7k7+/iXi9I59/R
ku6KqxpyoeKjFaAStkyZ0yxOap8/aqavHjSd/OQvTnB6Ibr+xisG2LnK1ebLuFo5
mmRaBOkHwtZ+P1rIfETmBt2mViF4qJ1TpB8vHTvPvZfQBfNsQLjabSmDSI6OW3cZ
byI75vD7Tvm46IKf0au9nLrXZnurIeNAZ/cbUkLJ1V5DgRjTfQrXg3mOF1k9L/Wz
kP0OrXg+Ygrc7+nYylg/n3aJnD09kdUTZKOHcMAU56DE2WvWKzvbKcYygs0YRQ/z
u1h/q/e1Zf1aC9zCKhKyR+XVtFpmAmk/SgsLariErVDVSdsJRlowru9jK49JbtYd
1hay8ZhihplGbwwKhvFfRUEl/plEXqbcUN5RFVMj/GSCXODmd20XufMaLZfznaXS
ebyjQEJlqevoPGjd2S8vrQd/qRBVnohg/Apzwm+rSJO/kKP0bH+yjtQZzxeonikd
dKYBDbbjmNaASeeLq1TyOGLnCOGSNTVN/8KlYNu+dCos1DgflL8wQf5+uj5CtE1l
ck77HSvnezWgezFo+Vh99y1dEFIwVtJYFDFXWwNUuRDdcjvYankvM6l8rVdOPjrr
g1cO9pOMkUg7yLxyGYSmE7Ij29F7vrzUKa8qq9iV+qJih5N+5gEw8X6+6xjq1YFN
Gwj5EW5jQyrCGMhxNKCW91srjYoB5gunUrIXb3Bxmj7zJlP5m88rfaRcDLfWIRZ/
D72PFwwqYY+5myO9xB+qtRWXSGRbvQweCMFe7uvrakK2rJF7hTqX4q47X8Om2q4i
n0MK6uV99eF7LvxaeHqLD9rd9S/FDuC3QXaXTEAqSEDYjcvbZo71w3DGTfTgZQs6
C2dGGQ9MwGfA+42mTzW5TTqhPClo3dYmvULajQ2yoT0DZHYPTlnRLz6g5zkyp7jq
wHjsO5VCy5uR79X7SWkMp9QtpuUIU+ACUrnBjQXj+5e9MAYTq5NYRmJbjQW/18mg
oK9sRNV/QXnSPWUh2q5R63rVQMGePctt9qUsXYv4+5VaFrA7CrEbnF/CfRgZBcYe
diFQcc1TDTcnY5HNnSe3ds/bcByzzqSxjTqnugL77erRyq9VQmga8wtNWni+7eXv
KwjXEBSEBCfAicPR1Em3SzsF7yBbYMuStCpeGRPO+a669inqQQL+HjRg5mj+pNmH
2pPYTA22bte1KuWMhWfCL/vkF0BrIYkt9pqK6VCkneeRJvqj4zfK4DG8UF4gpny3
0BiombXhrQlF1fCVTFPRbfHwg0dg5ygs/qGqhLkOJmHJHB3izJJH4t/G02OnIL3X
7TIm8DItF1cl7egBsm7HrDXwa+I+Fn7IXXUinxlzB5zM/9avFRxREg+4tFnZLmOj
G04XcS7dLgy4Ikh/qkgOg7TqZu66FX8+xxj/jzJnaC6T3Dvg9U3Nvos5EXNch34Y
PcdwlfhJZLjoPp6KQpGk2aKkB2PzGpyr752AtjBOLBHlwVOduJSsAkSmuANtUgoi
oRHvmrBpAzHqIGiort9jFuPJWkStmbNykiPnhZhkeMPT7FUh1bk5sBJToFI1/iIw
y1Tfr5/F2wkT8unHTqbAhNyULsLzbpIkCGwMACqo9qFLzaf9SmLNkUSvwEoZNPrm
VNVTpbTpnpBktMSfawe033NP/bFl1BiWnB25K9XZ4/wsuUQ4L2/ZibQNc45f3QTD
rsX6kFf3ZdAxGKsobkCbF4b4NBqxSe56Kpy01EKi+dzGWogpN61IsrMCROTlVprG
PL9P6DrndteAs4uQRSiYhUto7NjBxxSp7kb4lsqgXFs8BuZCTCowp2d489h7ROT1
AJvGCGgZQRn9eHQ1j/JyxgJzkqf57M+GGefMz/zica7lj+veB62INIFIzI5zTWje
/y5miouuQI77VnSdhcPgso6tnEwTDAPFXaD0gy4rxFI67y9PzRlSKWtdy/EVTRlt
Z+htlK0v9Zu6seEAv8eMvMM72PqTR86K8azm2qKX3uht0TDez7uS+8i8h7hv8nSa
B/EfeQWRtzWyMJ/EyfmD5VYSwN9T/Hhh8Hi886Y8vWUJX6ajxvVEpqonLdc8tHer
SiyYKlm+L5BjusKO1X3OoBsaFALIa6T6sZ8V4amLgU51BOsPAOgnmhdnAGVFnnAv
9ZplHk2mJ7/GcUJ+myBqNpLDi4SpH4XrDMQFW99dTu6HkRGnsXqI7XrAYRwzA5VV
sOFcSAVVni52UddF/Gq1KVvc8azoYTkW5JcwPJPaJdTpFz73LY/y496noYsUQB6q
iHrIiz8j99P8n88TEWtpYtecOWKX9TMMgXeXp058sX4xfbgUQMRieJoBXaonffgt
VQLtyOUysUwCUkGJZIaaV0Kbfr+pjqMZD2RNF3Xzt6NXGp3MB6sG3P6Tgvy3IEJv
9MQF8Ua2plpdtZ6bsAfhm6T2UL07cbDDn49dchdaenNWthfZXjM0+eXgoTHGSx3v
RlZHQfpWoLX/+ZYiQi2gHtf1zBIVca3F6vJEra4LB19hfipaCH+mZMfZCy+egm4V
vQY8Wn+sbTNwbQXVHXMpLunGjnDNj/BDBMgfVFTKnJx1SH4tvkToR72ORpkl1J2c
Jt0SX2dDs6UhSwQEV8qtyODNw/uDYJZJZLxI2W8m/pIZdj2diuEOg8k2FfITz03R
9uWEwfPQHsh1DwzFkSmGDQGBcTvIxrvF3o/iOi0x8NucGxvhdeR4GCVUZBmYqWcO
l2l5T4FcFwslIdONeVyFPiAjpkgmjU6zUmgkqI6UbT/gSVlUCDjyuQUFGtnQD3pn
NPUlmDNKD51kwAY6EbKFZnrugFYIlRgZJpoX9yOhg67RkfHE1rnMNZWCsSJrfu+Q
nV1zx6RquteRTBt0XUZNInj0du8yr4sRlaWHlfKnEOLLHBL4tEE00awM6q1wrF0V
hRyU7i6LRP9Dui7Q5MTObRIPNsogMWPJJkxoKyqAKU3FSxrmgMtA4dI1ARrfsCnk
CBTevoFpGvlt2Ge6byXCNLAmw4RBvoaq3hu6mGR1HpXqmJFB1BNZPFOZ2NB9IRfW
rG31y9UPngkkxnqp9EY2LnMbqE2oxXCN+2y5MKcpBL6C+4i5kcIlzEABZ8LyuZ0P
do9p7M0qYTC//jqOH5C/jW9wB3HdjyTlGFy0mEvjjeOn5JilAEwfJGt/qddftCjV
ATQq15tlnPD8QeVyeKPjP6xUGjxKZ9lBqYPcs5KS5GQqPd3rf8sZs6hTjZPi+QIf
JTPu7cdWoLTuQl0RNMOiT/7ymfZv5hBWPDLR8eDn5U+Aj/BHAbMNPu6vlpoNCaXR
SBOBVDsFA9QnhvqHvYmrgVVIbaqoZbA5XUZPpmCFqiWI0KEHd+oArBsUb+cMKBlL
EUCgxUCkv23v1OBW3PASVRfwP9Qne7zqPkcJv9KvdEU5PwVDZ77uPJT7xHgyVkmt
Cj4EebFRawb/dab6ILw6D/8fMT7bvuqGTOfbwW/CQLqtX8rpxZlnAC6Y2ikKrEr7
vWWWWn5ZGm6Chme+Uy6HwwGEiSMoBh5UN7W3TWkSUcU=
`pragma protect end_protected
