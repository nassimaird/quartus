��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�˅������d�xp� �5��B�{�	e��Hk�Z�徒��{��\�83,�p�)V2V"'������'v�{��A��L�J��ʖsk�eRGAO<M��a.p�b��@�@a�;Dep�r�p	1��"32G º��*ڦ���ƫ�r`�c�}_1������	H?���}� ol4,n����������\p�kх���F�y��f�T%���^5�����8
�2j��pVq��zK۴N��@� 0 �	��ev����m���z_ws�=����#͑��]�Ţ���FC$����
�4o��3[�Y3�v��� r�'��̷�l���S���W�v����E���1��_���Ѵ~���;�ﺴ(ܢ]9�\h-m蹞����3���Q�ó�?�A����Ƶ�̟(|����g��~�Q��6�tg��}Q>�CW��k�9����ΨˡI6I���OS5No��k*�D��p�(ޚ8�5���6����I�0�~����ǏFA�2�;ҩ7^&�'UNg7���ZE(�����
J�E��B�:w���'���W���;/�R��y�p����r��Q���Ĺ�х��9�v|e��E��(h�,k�NNk��xL9ӌe�9:-cJ� ,��[��.����r�A����eA�v�)����8j1�A�ƨg���o��������Ƨ[cP��^��r�Qfm&�ؿ����I@��3Ml����Ɗd/��gčZM��H|,*-�r|��bo{��@C��P�eV�c����C�u�μ0�3�,������N�X�WBC-���2St6�8� �7Uƃ��rX�p����4�P��V 涱�P�n��)\��*՚�S
��V����RO�����d�׾�����P�䈾��*�A� 3�b�S�|�>|0�X���w�g�g=/�CmL�~q��4|S"�p�Ń�%Dd��E���5��@}�n4��`���/�z4�5@���Y��R�����w�!�w׾�J����Qna�5X���\@��'Z��8Pj_1�$u;���d���Q��4���@N�<x��!�>>�P;NW�!���rm��!G�1M0I��/�Q�e��s�	�;'��d���e�U���:�AJP�2X��J��7%HWqZ�S�Bh�l�YX}�\���#�,|%`�:ڞ�g�S��P�c'�t�\SO�>�.E_�	3I�O�� \�]�-M*aL��7�h}����_�{8��\��}��݆�o����;��\��ք���=a0���o������k�y�\sC�	��Z奼��3�=����g�*0�BE�HN��#���	7��/	��_����uK��8�~q���kb����s�4ܽ_h�����\�xU-�R�2Ή�䱃�j��.=���+�f"�6�5knf��D�������,�=z��������	�ڒ@ȭ]�ܮi4��(8{���_F⦈Ѥ͢��u����u��y���,�	GwD�^}���v�M�N�!�L$?�9!W:��B$� y���
�r��f����������_z���+�jX���'�1^@cP=k�_��O>�&�86��4VV#�{��VJ����K*}ҙ�g�����B� ��9�n����Υ�-E��>��A��/(�ȻKm�[��nI��Q�1}�.+X^ed�Y7x�P$�RS�C�|ED~V��N��G`G8=h�#d8�3_���g�#��:x��Y��/N�޻�`��LYe�r�W[���xu�s{ �(c�jcAa��Isn�ir�[C��Ǟ�X�Th�`ڶ�k�7��:�����uw�ؑjR�f��Z�O�i<3�l���4K{(@�E�7���z�D��*A�
 !_��w��~�~'��qY�{y2��,�I���N��9�����Q	��%�)�+E�Tx{E��6��I��ԶP<��O�C"�0*|V���и�_y�_�'�N�����|0�p>��F���hņ��ŧb��,��>L�C�_Ҥ�e�k����w�%���϶�D~�f:�?m�Ca�r��◜��0�)�N;��Z�J}w s�R-c�D{�0{6���
_�}7MB\`��t	Q����;a��A�w^c�	iu/_��:�������8q'���0��, ��/�E-�7�\l��b̬��ql�"3��i8��[�No:$p�Cw���:d�J����t��	���HH:a0�K�-�4x;o쩼!�-�WZφA4fQ�"!_��k�U��\��x%����{�#m7���Eq���+�o���iВ�6 ��B��]p'���֒��@^-k�|�D�繽�m2$�������x�L�=X�qM���P����M$�4Bi^脿H�G��Ӱ3�!ťJ�/�tnL�;j�9��H��y�~
XU�i�S7�� �d��]��W��&�D@Qe�ZS�t�H�k����i�M����D��qa�wc��V�&�/D��+���`�i�����:�	XZ��І����l�U;��[>c�re
�;$͐�n��'_�Ģ�L$_��2kC����d���=n&�<(����d�n3�Ä��e�s���RF�DG����
�͋NĪV�SZ������ȋֺ��Y}~�˄����7�1�s���,6���?=�?b0�ʘ������5x&��(k�N!/���V���|��Q�R���4a;ȑ�ՀG�XD�UW�T4H_����@�N
���:ѷ���q���#H?/4���������;!
/@	�*�f�P��$]�J@a"�e����r���;�"�&�7m��etg�_�	�%�J �.;D�X~��h��[��D����uzx�m��N�{�ƻ���e`���}��S����k����1�rf�Rt�� ?��e�����M��T[T�#��-��<�ó<7�m���(�o>�MN5��L��,�$^&[�	����ഷ�^���t+tҽw���rq��T�U��.;'4G�[��
���t�l!��
Ե�R5��1!�iW^�kV��P�al����=Z�biB�����,�t�����Q�(6��S�RJ��-�^N�[��f�M򳴅:�H�c�DWG��ʒX���/OU�zDi��=gC���w����c�W�А�g�D�j�5Js���avZ+vǄ�&.���e�B�ҷ�H�%�����}ǲN�#^��hd��A:G�)l"�5c̪/ẅlgҜ���ܶ�6�T���0>��k��j�Ҙ�P-(���;(;�De�}�x�&1��^fRP�7;qx̓�;�
AQ���L	������)�F�IA�>�z�\�bE�3��U�O���:�\z�/~���&Yy�T����\��@X>γ(D�����rT�W���.��$ጒ��!���4�>� �F��2���G�P��D�@�P:���4���܅'�p�rs�����#�x3Pbe9[2@�<��$��߲a����~��qm@ݏ�8h��l�n_��*�D��e��pՆ�p�yiklTi�=��a���[_��yW��tEDXކ��	 O0կ z.v+��sL����?�^�\<��x�V�۝��G>�c8��]���4���E�!���;��70SR4�Ӓ4�]����v�Di��˭d�3�u�"� �����N���(h�]�'�7���T�Q�����/��������ǶGy���84t�4�H~{�f�MtO-|�g�;Z�d�H��(N��l�>�f�tم_^t����o&��&j�1����H5W��R��O���j0c��Ǆ{q�f��=�n���)V�V�;�Q��C8���S����V�637�p�i���/�$T#�2�xѐ����h�ye�o�Nt��G�`��d�Ӌ���Yn�J��I��g6$t/�9I���dMJ��Ξ!G>?�%�+3;�''�����3���H�Р6�t���?�H[��"J^�i���u>^;�5�;"�����|Rq~KZgG���!�z��/��w7�ь�-�����S@�/�)/&�7όE�K����%�|�E5�N��}�g#^�����T[�P�|Ȅb�.4T��6���`��bH��lH�>��I�1�\���]�E$r����Z
��/�c=|b�:~��cH-�kN<U�]�
�4����`!��>�L$`~&"��>g?��>Ǹsé�cJ҆��C
���/ik������'։bl/��PG~�\���Euh��حB|;��p�uM�2�|hl/�%E��-]|�Sc�`h�=�R0�g�s8Ͼ��aO��Ǹ8#��#2_��G��ܗKL��>��.��y�]��� �i�C�q����+�EqX�u�5��t��s�������&��l��|+��>�� ^I�E<@�ب�6^KQ��q!�3�P[WC���Ni�|���g�c�F�vpq��B�/��T�(�fZ�29®aU�!�%ؤ�]�%����_wEU?�vt���.�%�M,>D��Z͓l�O",s<�c|1�K�
�&[D����ҙ�.�����}dz�K�G2�*�"s��%Y���.`���|^Sמ���vQv�.�!��W�����ܵn�U����9k1|Ak�D���-M��y�V��"3�|U�A�y^l�&��i�`P�l-��̵r);`V�EW0��uڥw9��<�?��d�֝��45�7;�p�y9�F����D����nL1�`��6w���ks��n��_�k�����XS��
��1%o浥����D���n�x�蚽��IYI�(�I��J����z��,V�@���{�n^��-,^m�^	
�?&q�S�� ϟ�������h�����M�L&ܱ�G�1x��I�qQ��LY�"K$t-�#�����rRm���~J1������v��Zܜ���_��t��B�g(7I)�0��?���C������Kp��K$h)b��w����%��d�^T�ܥY���2�4r4W�J�XM��z������<J�4��Y��� �Y�����m>�X�J��J�+{x�[����A|Ao�;V�������A��,���zHK�!�/$'B��<~끒��1�N�S^3|{R����:{�4�ޥ����E�=��v櫡��5���~���%v[�v���U -��@�V���5;��(�t��,"���g�Z��_(�C�;]����Ӆ?e	��+ç�;�����~�.1&�U����.�t ��'`
�����rqs��:s�p�m�x>d����D����kr' \=�9v�kڎ��D���ř�n�MIP�Z-��ijS���	����xmL)ic����J�;�Ыf�h�|���ܹr>n�tC6ޚ�HۙS�b�|n�͈��mv~U��u
��-�<S�pH�䈲��ۚ�Ǻ*��@�}kek�Px�μ�|Ɣ|����*_�X�ѵ����#m'�є� v�CG�,���QBT�~8PYT뾂��)��(��<;�'�	B�b�j �� ������)t�f	>�u48�)Ri�F����'�ꩇ�S�L�`��,�F�U�����_:��=��ur���B'�\+^Tg�7�:"f|�	��6�cHp���Ӿ5�#�nd*�����L#!�P��4AP'�25�4b��L������1��x��g��*6 qA��"3���[\c���\�]��-*��̽����r�H�E���Ͽ������Sf� �^�÷�ujE��ͫ��Ƹ�����U�p#��M�=�:�+|
�\`�&5|=����UX_�^� �Ek�b�[��������<-��:
��< ��D#�?l�������� (�@��0?n뾴�ĝ��_�be�8����~�Qy푖���5�p�SH�:�����[�w�Y86��,��y~���ĻՃ1g�	��,j+�^>14%el����)af�+�@��*B6��u���s�$���m~X1`���߹��� �b������Y/��l�3����"�n�=P�p�vw���G��\];�;�����NR��<6P���T���^��5Ͱe��1K�-U�Ĩ��*��\����\�R>�7]" � �E�C�dVosA��_�M�Byzh����q��5�q���U'��9���Z���p!�Ns�
y�Fpo݇ei�Hsj3���\֞��E��.�`B7Ό[n���ʴ�F�zX�`ٔR�w�}�����i#q��F)��ڏ�^��f�Q3k1#v�[:�X�#��J��\(�/v��`�f�t���`��֣)l���kz��)� '\�k�I����P~��g����}-Q�@�(�w,�MS��J�e!�E��=��0�7Q�^W����j ���6�UHo��;;�h[��H@�LE��^t�-�9���I��Ul4�G��ғ�3��(�Z|���^��d��2M�0T�'<oTc+�]���@gx�ܷ�/V���w�eL�� Z�]�)���P���tLN��9� ��Yz=~-0o��;��>�;����o
^9g����kaC��)���Ol���ֲ
]�rg噻E�f<�����B�lP(E*�����;~(eg��=@�i�kx ��f���lR��)�A?_��Ҹ� ���T����
�S5�DL| �jg �H3�J�o`���rؒz�ͷF\FP�lF��g:�d���8�;�Y���B�Y>��ɉ���RM�)쯗7��F�ڗ�[D`x�vy�/���(pldm]r�`��q��iZ���h� ��tbɨ�2}�6!:���-4n	����O	Τ�A�㑶j���R���P��R��N�DR�_�����+�������RI�V8 c	�bv%�,�O�?�����#��B#+!�6�dЗBy3+~�Y�zO�K��1,�_芹ģ�6YQJFNd��6q,�g�P9��}%+�s�b �>G��߬Z���^#��#=Rֽ��:/^+
c�����}�XQ�T�V�� ��W�*��Ub�q�	�0���<!"q�OE��vI���{�d�q_0�Ġ�سU�b���_�����w�o5�G�>ɣ�ļ�����!�0`%#���Ｂ���q�6��0��e�H�ݤgH��J�n�9�T�0K8��O����-���6QP��MB����|l��8�DL���Z>�m�ǎ"��MN=_�3Gݟ;1�e]���H%���hd�c�RIa+�0�.�CIo��>���Xq�����;!�����#Ŧ��|�D����I�T�ơ'e�m-�*��I��T�	�+&�d4��/�썹��,E½��p��J�A:_<��2�b�cW��)Z�O!D�ˏP�2�l�:�¼��c�cR��_����m�sx�����A��ґQ�p�v�������ٖ"��,���ꍋ4��5P���֯Y!{���������F�O�<�7x(��SOʨ`�R5J�S�.�������P�/I�3e� �6����d�.X̥��9�f��Hu�� �L��KPVW����r�ޒ��e~95�+<eB���=��%���Y)`�]����ޝf�tWCک|�}�"g����M`0�x�1 B��1]XY�J/Y�%cM��M"~$!Aح�:���ZR����~����?�`Y��ą��:�Ǻ���}�K��Np�}�%k̽��3����G��4�a�"W巛�m�%���HV��a�۝���qBԷ�a���t6�v5&�ͼ��t%w50�����C3�7�ۜD�`2�����2s�����w3��}�e���x^�N��w�Y%×�$�F�S׭��is�~>�;�^����P�\s��
��f�F�����&�}^z��������������M*��Q]{|��گ��և�8>DY��#�̽\��o,'p��J������,d�U�vmQ�Ѳw�U<7g�b�z}�BR�K���ǈ-�B )L�5�ȱ�p�SXàW�9�㻔�zW�@%12�H�+a���\�b���t���W�\Ϳ���-�8���yϟ����&���	���9E�W��ɵ�P�2��0
��59j�nfue��U����V���2�5^�1���N�H�;�� b�6`�f�x6|٪�������D�$��_1T��o���'�\������(�Q#Bh��R�rfE��L�I��K���w�p���?=H.W�{��MҧG=8�kry{5sЍ�Q��MPL�ն����֨�ؽ3��~�G��4��,�+A��}ÌڻW�J5��aʅ/�~���/�Z��n��L�D)g��A��K�� �uҠ���j��7�E2en�tٲ�uw`@�сyw�N�i[TJ��=1%c�˔�>
y&n�n8���^]G��՛'<��{tC��Ѭk����w��U�ڻ��#JOb���q�4֓���	��
�C�����.�O��ǳ���b�Rh(5�E>7�,�B�g�Q�E2N��+5d�T��/̶����	�b"���2���V"��!ɔ0螢l왍�\�bL�ZW�z��J�g��7R��ܷEN��<��.F�.�u2��]�A���+i
���;��df���!�,��f+S�#+��'X-dr�Ǣ`1�m𽲣Y�����W���ϧ�(0t���8$�8�/�pQ���j4Rxc;�&�F��[y�����=�a���dF<�,Xp�m�g�d=pѼ�_<z���Z���>���t�F2.^qdD>Za�I�`\����[�}�M"��-�\uN
/m�1���Pj%�Ǧ&;�jǠ�`GuR-�I��dђq��lcu�6�3q���L�irdG�;�e�\Z�����w����dU��Ҹ��]:8�e���jq_� �K��39xJK����WR��Z�Q��ƜdQ]#��33�`=
���{!ԴJ�"�������qa���wyF٤T���s��J��	���>b�3��+�9�k�j�H;ji��0P�O�>; wpA�c�T������[%ɇ��ɓ������Rm5���es'�k�������3��q����Yp���k����I�*��S�<�����ں#��&��}ʷִ!Xv�_Ec�-@W�;'����Z��6�X�M�fa|iG0�1�^Y���j��MW���H��!U�ړ���9�#�Nif����l5��z�K=l=.��\*�>�sS�L��/��U}W��P�5
�Я����i�TUw��*	�3EC(�Qh�%��'�_�0�x�RX�jٷ�㘉厨c�4��{�]JD@?Y!�?��+�#h�WNkh`	�\���U�!����\a�n���W�g'�v����Ҿ�F1�E���K�{q�Hz���_VL=ݳ�ގpVO�*f��m�Ŀi!�4�zts\���/\9�MB!82��߁!���u]&	씤����ON�ع����Ïf�䦋�WB����9��.-�q.B�mC�d�M|9;�e���5���^�t�t��ǯ�U|�'~�@<UI��t�k��U�i:�HrЄ`a��vc/�^ �P�X��V��e�u�gc80��v7��v�*��n8���e�#i.�Q-�����'��lh0��CR��^��щ	q��+i+1dY3X�¼�9�q����*�?�Ş3����ܶ���nU�s��3�*���RNCL�M����
{���_Z��xP��B�ip�c��I�g�X�w5ˇ���\�D}��LPg&�CT�NR0��*i#���WQeuq���'��tj���J�e�S��7��w��gڨ��)�m?�9Ut�(�V6�u�vu3��>4�5fi��.��0�3��8>�B���d���w!�A<+Ժ����<�h0\��P��4^^��|ciP�N5�j5̩\����24���Ë,�U�զ�3�4O��r�����ՙ��Pg1���R���'r��{�O��@HͺА��x<nD�a(�G2��yC�#/�զ�ƻ��-������z��t�$Z�{o�0���;ޡU�F���Ư9�_&����"��tA�)Ƌ&�+b���w��꿔В�DS�۾�84J��?4�{.��(%	t�}|����N�PJ�>�%d1+IM�q�W�?�!Xc�Ҫ�W�9���O��N��	��G�re�{ܛF,��v��C��3t�u<�"�&+��)�x�Y�{���9�D��n�I���1_y��9��&sŰ\�y��7O�ISA�O���K!>�����?ht�β�����rT�jӧ��cV�w�m"�1L��#�צ8_,������૥q���j1�+�ٽv[����%��cC:��+�.Ԛ��=Q�U9>S�p>��qX��sأ�ɟw�J"'�h!M9RĪ|�,�!����ܘ�����u+�l�cH�h�$����M�q@Ҿ���')������|��i�p�O���4Æ���ơ4�QWҐ�r�࿍����A�x�䯄+�
��,ߌ;�1B��������D�%�s6m��)�[S����`�n���&��P���Fk4���oF��3�+Q��������,�C���ŢI�?Ea�b-&Ĥ��j�%�d&�a�Wc�U���g����O��S�h��&��S	�m����!( R���ނ�ߊ�SG*g�F�|���w��^L�ؐq���oH:g|�'�"���ӄ`�����F#ڂU��[@&��,���۴t��	��\��4��Κ�N뾹gr��V|�8ޅ[����H����З&�[k��䉎:��[��+��"�iK��F­��`�`CV/�|d7�dbv­�,doW����/������_�̳����D���=S<�g��[:�ܪ�i��l��BQ�R�(�G �g��/�]�7�2����V�gE������*$6�e+����\���Mw�5��K��Fi�������:7 ќk ���?̤�ɱ�NXO�5�8���T�� �c4����=A�����}j��Y���Wv���&���yć_�l��\��$a9�Vf�����
I��ō�J��Fn���"-ֻ_oo��Y�UNZ�g����J��mߑ��(�<���i��7��9�u! �%ߩ�#��?� �����%����7q����?N~����;6tRl�ś"C��F��,Ӿ��[�6���I�����"B���X�y��-�T�YMz��a����&��@TV�c�SH%����~oT\"+�RhDj��@�7���0��&�j~ՙ@۶��O?��hg�^u��N<&O����9�]�3�Z��IF�1K��%�q�zɟ�:]#�|ŏ�#+��f#��
�%�`\q��cu뼞"vi}s:Ʃ�]����b���3��L��v�X����u�u�ng�db�i�〝N:�,���Ȥ���T�X\n~�6�L��qKA�.:�V�kw[�)�ܶ�).���:e��}���:������{�ٸ�C��9�,�n�{=mR��m�_F�D�@ނ�d}�.�I*w�Q�rd��5�	y�jk{n#�)�z�nk�ˀo@��� �/͊��/��sD���Ƀ�$$_F:�
6y���5���{O���7v�Űu��Y%���Ύ�dt���rm�IH;:9�3I���i=�U4tUk�U�gz�M��TR�;�1�����*5���]N���W�z�Hr�������!È|���[� ��Ҟ�md��Fv���2W�}�/�Y��*���k�B'���ͅ.���������<o_�y�j�lH�GTE�������5�t%��>��Ҋ!�i����p�V�t��ζ1�_�;��£2�&�ni_4ɟ���#��x~3m�к�x��LY�GQx9�
B���n���tI�P3�[�o����LR�W���+�4<0wg^~��Ϝ!I%a- ��8��.b�yL�L�5�Bt�Hz}�J����M�k�a�Fu�.L�
�.�M��RpfWmɘ~��Vd�<�Ъh�A�
;
pŎ�4�6�ˀ���x{8܀��-G�	�X���`����ѩ�%��",�b��c��>���	�������5��].0�`y�x4U�F|'ݬ�-l�$���z���[>���[��@��O
�qI_j<%�G���O7�c'3��9�-�2?��鮐���~#���pw�0�/�s��8�l�NQ-��lc VO���W7�n�$�tR�z�X�<g��}��'>�B�}���]����5�-�hՏބ:{W��f�	Hв��s�7���>��M2U(��y���� h)b$�  #˷+��d���b-Yn�����u�����,Tg$,�%�
�7-�GH�N���m�o�9/y�qYk*?�����f=�$��~W�,Ծe�גi&�b���0���71�_�!��s�u���tKig�}�}�0�uhe>�3���H�QV�R&�%��ߊ{��mo?�~B��'�PT	�_x����;���2Qrj�/�Ć�%n�t.��7���
a�Rvv]�������*bv�#�������&'M?�z�n��F�w$)��l`�`������<��^�-���VQj�{^̇����&#L�F���zUx�{˛3V�v�{��)֐�I���0����T���^��,�Tc�))J�,86�	d��b��
J6�r�Ұ�������%�?z�I'��1J�f���I���\�or���\W�_�x㍊��u`��9ol�8�Ên��!��g�(1���.�g�[OYS���i�.$�R�/�g����0&E%���0���.�$�B�w����ס�m�a0�����.�v�%���~���f�@��D��J���FoT1ء{w���6d�_e+�+��%A���/��w���#�0�����{H�����V芜�[M�cޕbƇB$��Z:Y���������1��%H�2 �aX����@�wQ�?���VQ9�˦�C�ח�^��3��h~|n�_�hGi���<h��R�ށ|zG��ͩ�S��m|2�Jy���*u���B9Ԟ1�GzZ@T8�Gs�9md`.�Z�j��.�L����J����-D�5#z�LSp�{�0��o���רoϣ� �Ɓ������+s,G8�nL�R+��O��ٙ����QJ��`�����،d��Ef��5�/ԮF�k��%�E�!����8�?ڴ��!�.�PoI,�X�����Q�*'8�мa�m��#��D5Yhz��##� 8�%͹���#�sKI�,Gh��v��m�>ަW�~��J�D��0�xy�IQ�(�w�'K�jD���B,x~7��' 8z�0���@Z�y�r�z��ʵ {cQd�6#�%OfLڦ�ѝ*�,�Y�����ZqRzʟ���*���8Ͼ������;#����	Q���6�r��wP��׬JB�B��8 �:�l*p9�[h��0���j\\�)��|��PQL��w�o[��Xa^R@��W��Y�3�R�'�P��Ņ����U�V�=.�9�$"��m˥UĻZh��Q�}����ΐvI_�*�_�����nhBKB�;����GFÕcK	���_L�㿨��Q�]�I�e�gM�bҗ�Ƅ(L���Uq�5D�+�����C��_�I+~�$V�He����<"��@�Y���DP������VY�����`�&�*NN��7��_>��U��uV����N�"#��U듽��TW�:'��p].-����^�ARm�ĜL)�A���/�6/�+����%��lp�&m�'S�PDGo�a��@�nAvR<����0�'����zR�HD���Tю�G!1������j6$b[W&��.8�5I�9�Y��:����[�h$p����k�6��R�ģ�I3u�����Ic�i��1x@Ԃ�Nv�kQ��.ʞ���pQ�P���L���K e}Zm�8�S�C��,)^��H��|-���s��HuTP�UM)��K󷶑4& �� x=q�VoY��wY�l2q<H��uPgiu�h���p-����䵼,��N��ܞR�����6�َ%QR�/�0������] UX�w&o����Xz65't����nW/[�nV��f�	:��J-x2���2������=6�%x�Bc��s���;��;׍�?�eL3Ι?�f�O�:��&���m�ӎ|��������a3ց�"�����Q1a���0�@�u�J"m'�*���.cv6Ջ��~3�S�ǰͳh0�p+S�6��^��7T�7��փ�� �E���E
Lar.`/E��h;ƅ��(t	u�P�`A�vc��]���#���(`�-�$^�b��+�
��"������6&A������{���ȧ:O�R��.fGM���Ô��8M_˰?���ٯ�r��N0�޿ݳV]�8���#ױ'{�e�q[W5f��wi�$I��eT��z)5��$�G-xO�Pс&�cj�%������KS}��e�8&/���G/���� ĪP�F1�*��"����u��7�M�a�i'R ?j�H��S��M�)��|����W΍bf�+�8�S�L��^nm�����e�JCZR� �s�/�r���%R;�ȝk�`��\h�Pq��%�/��L#�OHo��A��k�m�W[�6̢�
.s|�/qF���{� �)�o]P�O>���]�a��-� n�u�hR�z�qTEє,L�ܽP"�(/�Wz#*��b�d����O�C���5�O�-��]#f�l����hHIM��,�}c^��L֘w|s��=�>i���=��a�߃k)��>_�!��T[v�Ć���FWsCH�h��d��jD��~GV�z�'�s�}�C��N�a[g��>	��w.�99�iI�:�eV�6���3�;�s������;9�/� �z;�j��0,�R�|<����=��r�(��-1��Z�Ys�2�wr��\Z����)�B	/�dF"� K�����?��R���°ZR�4�{��\!ɄY�{^1��C{&�m-(U�djۛ�dμ4$��Ep�;@#wh�J4�X�oa&�1E{��ޱ{f1��i�c�����Ks���@%LE��p,l���+e���W�FǞI�a�H�l�v�AG�E�D�ۺ�t�t�P�}��sD�C��螡ɍUȾ��ٙG�߉K?r=�E�%�WZp��D�j�M���6�|�X�1&6��@]u�,*r�E��Q�U��d/����k|ǉ[�p�%��i��,߃G,ui���cl����~%�qP�w�\�BC
u�G8�xBMLT�� �C(��q���2�G�~R�D�|���2�2A"ؼo��!H��о��D�)���� �k?"0�J>nv�z�Z��щ��3P2�O�N,Q^�@��E��N� 1ځ��e,$p���>�f���8H���Qu�,!���n���,��x9��%�"�i�S�F:X��c�*5[��ǔxe-�g$���yp6���(JpŃ�o��&R����8q]R���m�����@�&C�XMݯ�UV�,"�v�s�� mڝ��s��P��5�E2S��d�$�_�1A8�
o�d�½(Gk�wKkn�vz���+���2�!~:�s�Z���Uy ��	��'��
:���c��VI�-��[�7w�[�d8Yߏ��-7ժ���r���"���p\���m!S6�z�}��`���+c�ۄ�B�s�}#�)��@��9�5���i���AnȢ�֬�d/�׽���^��~J�6ugH���zk��7��*3IO�Ǫ� ���I�(`�ՠ�c�����2s��]���dn愜r3��8�ߤx�3 ������ǔ��I���UOZ���_gv�A���X���q�}q[����du �$���N.���(D_U7��'Ѧ�����6N2�0R�%,��mS��5Iz��
g:�����_�$A?�������O�}:�Py9��W��h��������e`"�����+M���7�v?����l1�h�l�+Y�G�LP(��D4A�l�Rg��V�J�C� ����T	��G�\g�l_5�)�b�6t�.a�{Ѫ�~ysw�!5�OJ�yM�v8���S=���o(����f�i�.���� ��kH�'G�������Hߊ� 6��Z٠\�"�(+�&�c�w��.��H�(u,�ȑr�R�R2����7�t56a ��O����R],�?tꓵ&D�\�������g*��f�k&
�ʓAl_����zs�Gh����&�%ӏ�<���ԥ3S����"�Kވ*H��}D��"��>���sH7���ρ"�$2�1�(�� ��~ |��_�!q���x�4��݅�T<��l` }%,�(dp| �.Qy(x2S���8D]�E˸��5'�ټ��/�cI٘��Q�g���-�
/hcR��¯�pN'�h�K�U���7fs���B�R7L8�����69�xp�칃[P`�	f���YH)���2��(�9�k�����J=��r��7fG�����a2�q�H��r���ϡy��֑�#���bOLE"�CnW�B��|�%���-�y�A��+��<�v�+�@�)�]v�-І�g�a�2
�9�������Z͝�l��ÓmA{��5��a�0� �P�L�'@��$~���XJ��r��f�X.z8.G<1��{E8aMj@��͞�5���bm$V�O��ÒB�P�G z��+ک����^4Ҁ������"�u�sV��m﬚��A8z��|��[��W��Q�@����$���3.�ϭ�L��߼��	��q�4,��֬�δB0�s�����*�s0�8�aw����-ĺ�1�˲�u��q$(,7�Mq2�$VuNT�!F ��+B ��2r6��D�1�HE��@
u�\�8p`�%�n#��|��B[;�0%�7�?�؄T���p⤪Хr�^�LC~G}I���@�n_��z��)�(�:v�j����2f��.�e5}��N?��I,��+a?�
�o�@�n�YV�x��~!�th����0 ����v�f���I=�A̊JyD���F,�T��G��	��B����%|�m�3�}ͧǪ/&:�5R�����䉅����u��9r��} ؾױ���ɀ�S �J[��c�(/�_o��4Yî�BT����漙�@������\@���Q� �q칸 �7K���G�o�rk�������FJ?�~	M$�nv��A�w�V"�<okΣb���[3��"(����c�����q��+��*|���qXW{���PZ�\���'���'��T�=,�f����#$��	��C�X����?�����7�٪����]o�8�e����+������IB�W�!�OSY�7��Z���{xH�Cڃ�����J.0N�P������z�D����ȗ��_�-|��܂���k���w%K\l	��<A�K�����~ϫ8�U���E��.�H��E˛�7�f$TQy%|��K9�B�><n''���@s����K��h��.�G͖7��_uAF�w�w����Xv��h��<��Q�!��E���
��o�q��^yq��?��ֳ��c!d4nP ��_��Q$�e�~
=���\��T�Euk8E�>^�lň7�'�'����Ղ�Yc3����;�,�G8t	��T���� ��вm�V�X��%.�۾EB�N�iZ��a�kU�a�}]�%�`�{{8��������rSe�����v�~��Sp��s��^�4�\F��P�(p!u���C}s�WRi�q�?�a�yy��e%F�"�],w�I|gS��}7��t��B~UY_����g��� 8M�pꔕ5�ہ�
�ws��ݓlMk,?�&/��G��X?���B�6@+��.n�$y��=�뤽�u�js$�(��G�~�*�Y�=����rþ��{!�h^
������)
����Ah���+]�F��#q����q<��U��47�Hک�.�]��C�M'*��΢��֘��5�B3C��b�N�H��1F���7�0��w�Bcۤ� ��v���<�vF[��ʿ4eK	S���еo���E�y�'4�eD?��A%�Q@܎v���'�p؈���)N׫�j����K����+_��5%sK=�1�1s����SAB]��>
R��z�kt]x!z���fu�ڐ�8_^;p�c#������ȸ�N���jB*�[!�v_7	����J���F���M��񇔎6�m�\���jK��H`���]���\��.��f��B���x�OHcc	ġ5wV��|�R� ��b��T�=�׼M}�����P`���4���be��7qE��j>��~��Pf��T{��0ځ98ƕ�9��h�.^�s��@�׷�}p�������`��\����8�� 9�ЦZ¥���%���ָ �R9D����~>��U�aѨ7�gc� ��|�{���z�@���6��w6��r�V�!Y#9�u�!�X(l�r��Ao��:�[
{�
�d�����91~�+s��R�`H��3˖J��jv�D9+�\�$���4������aUa���9�6Pu87ey�.h�+jj��Q$�������#��]K�G5��p��x0j��$ޑ�5�J�bj$������Q0z`��x��:Q}&�4���ʮN�"��*��qS�Wz���s��S�?���Q�㤏�BΌӯ���y{7~��E�E�����൤C�0�ث�3�c;��C�dP���	h�m��V]�I%#΁����<��%E�㭳�������j�j���g�P���9�0A��rlpcv[xb��1q�j������V !V�ۧ�nb�{k����Z1c2�/��?��c��PN�]�t�;b2I�����f�,�FC�p�=٧�B�p�*�T�'�1r-\7wn�B���P|�ӞAD�0�#<�H<no�'���n&	N�`> �d�M�3z}l���Vi�r:x�I����T�[!��G�q�{tX){���A��/�ڹ�͘�nT�ZX���U��2���lQbd�{� �Ȑg����E�����a$��,p��R N1|GarS���D�{�(��)rHa��,_A E�!byd�f�ګn�tٽ�yD���I@�C��m�������^k0O�&3��)�lJ����m�b�����r�2H�jL���ߧy��ԗT`��� ��.��Dhȍ:�����< Ƥԇ
�O������@	sl�S��f�����|�>��}�T�ݤ��;&\ڝ�&�SN�ܼ�����$��X��>�	�@�|'����9q��vDq]�H��#K+z���Fn���W�)q-�Q�r>8���N/�S��9!'}�G��;+Eĭ�����6w�B�2��h��G�����x�~�Rh��3�ˇs�Bw/��8����d����#�6�&^�Hٶؔ@sg�	�DM1�;�L����g
r=�5�'��Ii��V��=Tg���*� 1���4Z�W�9Xռ"�|�kd	���`��^�]�f 	�Fpǃ����)k
��*�{�z�1�3K�q�ܼ|٫��aľ����'�s�|x��v�ɹ��q�˖����!���Z#�-���D�o����G�وO�m��g�7G*~}�:��V:�EHt�D�[Œ'��uT����5y�j^OM"<Vt!k����p}=�v;�y�ƙ�
��4�w�`����'e8x�ua�y{g���xTVmԿz��{��\������^W 2E��iќ�a"{�<�&�G��jh�A�o�
�u�;)�K�iK,2w���l�������A�L����t��H�#T�TS{ۈyQ�i%�勾J�w`�8���*�q�'�1��� ����Z��;��f�"S�=t�fR���ْ�0�I� Խm+����a�&�O�S+�J�sB�S��u��l�� �*-�빱�YD����~�qhĬS5{�gƭ���Ҡ5Q'���M#υ�6M�V���y��l�0��p(�U9���L}��ۿ�=Fm���c麻S?DM��x������nc����~��ގD�v4�����Cz|��Cv���vP3,���������M��J�haNO�p!�C��Dߛ���f��z���0|�uQfxx����������~E+�xiW�R�2��#[��y�W*�V��E&�c���vi`��F��Q|�$k�;����_��c�
ۤ`4ެU�F@3�+�
,Uk������uˑ���,����s�lX�E]Uu��+9���"0?�W����ʞ�w@^�э��Q��#i��٦�}���޸�1�n���7(�������nK=S�����>	SD�tU%�x��j�r�@�z ⶡ��[�0��J<:��ٴ\�d~�SN=듐���ܹ��)fĬ~,q��E]C�l�YO�)�	��R�U/�z9@A��)W����v���{|�&;�M�A�3=�27���Q���w �*x[a�K��	7[�D��o��|W��s�T]fЭ%u�NS?�ݵ�&�:/�=�j,�Nys����K�AG���pJ�5�$n<�������N	���΄��z���w�(C!�E�*����</,HfI ������hG(���e�0XR/�/���6�q��!$�Dk��3,�	��+�������J�#ۓL��'���>ȈM��Ι�;��`���������Tx5&��ek�5�^�jo@�-����y�;�e����N�?�1��X<��8;�V7�[~�
�%n�?�Ա}X�h]�C<i�7�r���r�����[�2"^hsظ7�QF�����{�$��uS�./������|��c2-C&DP�*t7��&î��!>�f�e����M���|�C��p\��5���Fh|ՔLJ���L�k*a>4֘��!��g%� 3ߊY+;��Rf����
 Wl�����Xd".lsm`I2�⳴ؑ����A%V؀b�y���&�0�n���M�m�%p��+hN2��/�+/���K8�.�""�t�B���ι.1��������Zr�ļ!J��ۣ���L����[��7.�c�)K�x��%,)��t���Ç�$��T"3\zn=C�r~�%�`��!8H	Wev3+X�U��
�,��t��B:�L��J/4ғd0	g!��'\�3�ѓ�,�2R�Jñݘq���}�9/�#�Y�ƴ=���)9m ������,c��p�	D���	����N��lK�{Wa���U{���/�m	F�w^���7	S�G��#Y�Ҋ\���D�Dқ�
^|�<q՜Q�0�w6�H�Ir4D�=z5xxܱV`{�hM�]�ŴZ�� �.Κ�^1zq�:b��9�L�|Q�nњ
��4���X#R�^�7��bQ�m=ǆ�������}��
�4E/�1�����p���8��^)��92K6����RN��S�����u2U�h
��W�h�[��_��e~Rb$�����!��w%�����Vd�%�˘��,����u�۔	���I]�W�Az��dn?�&���<P�nPOE���',�̔f��ZD>�2�|��t`K��K��D�b2眍��@)�kSG8Se��N�u^��J�uZ-���"��o�F�6/�~#�O�7 �%���"�}�t2���Yx��8:������ӣy��4'1�E��R�����Q_���=���p�l&o�|��ڿ���:G�Q�d�I��H��W��)樲껁�Ň�-�e ���ef�1'KȌ�C�c��o��%)(�{\�E�;�X:1i>����T㈇uI}�i���7�˱�o�`Lw�k���(Ay4�Q-0nz։�{��N���=�H����kk���ϛٟ��V����� ��p�\lc���qǟg��Pǫ��%!��6�{ċ&m�a��=��p�2��l2ww)���M����<�(�P��!Щ������j�>8'u`/��$Vy�L��ު����k�0�!�D\��c��G��vqt9@J��3��U��6�gf+liI��O��� K��c����e�/�lD��Ye$�I�Q�,�����$4���0F,*."��6.;q���$�.�Õ��83�9Z*w3WN�h���ݭ@��N��J%��5��6�47H�pzM$���R��L{�ZP�dUf V����'3�`��2��dͷ1~,i�p�p��5���T(p�5z��P�'h7��m4��d;�MF,����`�3�^��k�ɑ���v��.�ҝ6��ĭ\����11����,M�}M,�dN���3/Mߧ<*�.o���PǱ�������6�����֦pP��$'���Og�`S�Ԍ�i�,$�L��|����R���X�)�>��[������4?H�I����^\2c��K�V��*L��-��3߽od9�����ɚ��4�4��ӎ��"��(�_����-cI��9M^��0�&�&�
�fڮ��]��C�wx
�?!3�8�m���F��n,�Z`��e)Hz���p��^%��XKp��B�u|�z���D'��T�H��������d��Z(�O��g'G���!�O(�aA�aHcƤue(%l���0�5+���E(��g<<��I)A@1�>z*.��d�5�ְ~Ip��A�-�}�ƮO��<G���z��'/Q�n1��" I��r]
:��z$/�Ѽ�_���BE�T4���1��*�md����h2���!j�P3d�MYe�hʊ���h�Z1G��\�9%%Mf 1j�:��oM�na?^�1�eS\��gc�d(�u��sJ�\HM��NDzHa�^V�R�o�7e"bV|ֱ����B	i�,�d:��L�	��s+ �V�_�}��2e�[�y�n�����E@½/̼��l��� =D�Ǡ�'�<Ɛ��EktlF���?mQc��M�wuB73�T�Ʉ����9� :/�������ǓY9[����
eS�mA�Py�
֘�`Uu̾/����N; �h��������qр����� T�������at%���4}���!r��eeD	ͷ��� �;�Pgp�f�=��O������O�$��!&Q���~.��L�s�����	��VY��Ddd��x��y"�r��<�-Rx��WcO���?Em��)A|�7qCyB��y>����+�z'��j�8�9 y�0�G��-�K6�aCU3>	�"# �9ab?�Z�B ���O+��1���byP3(S��n0���>~[��>)��"�|�f���9K��{��'� ݪd�����֍7�P��_���b����N����R�I��*3�*������OH$�,����&�-F�%���"'!�f��\�`~N\�ے��A�l᯻W'�o;��7���b���ݲ��BJ���5�<0�3���6)}�����S}'����&�~���\�<*����=ϱ�Lvo��pi/ן��i�!�o>�ي�0�8(x���'{��t��Fo��������NlƬu! ���"��2 {��x�	�W?��q�%�4�ۊ���X-����eI�.P�,�������`�sߛ*Q[����TG:grs���o>O�T�)5���*o"ڻC�Qou�6Ka��8r ��?�`^�[�w����������v�
��,��b~w�N�UR�v�~�?����Î^����ϳ(-6�mWDFWB��m�2uL���B�챵"�r���u�[V�_��p�*�CRZ��P��J��H��BD4x��@���+ ��t_�R.�&�G��}!`I���,�"�5KK$MɁr�1��43�V%Q��L��EO(�ъ�k!&�MG�Ŝ�R�.eWq[i��&qI**�/��E��LG�a���2��X��tds/?R���vԬ�S&�))_��Կ?77���S����H�0�:����ƇZ��m/]y���	��g &Q>ɱ2�17��V9�$4�蠘��5��u#c�	�R�%���w	�5Y�-=��tP�B"�a�$k��ɨ�X*��o�|y<��P���j��/rP�O�	������q�C��+�zl�d����ԩ�{��,����	5B�H=6Y����_�$ ���´zHu�7�lB]V�l����2\L�.��*�*��I䢔m��R2-��nC6[0�P�{�!�5鎭�bZ5��#�Ʒuz��� �H���X1tE�����YJN�=��A�voh�(@*VdRB��zYn��F��?yL��OV~�?R��&�W%?w8����#����}�܅gɍx��
��yN���k3�/�/���>�B@��SG 6�W٥0w����h�����4���<�r��'`��2".���O�c��3�Z	֓�Q�?M���R�����?]�Z�;oʘ�� f�fe=��C�67]�p-�C%c�����[�}�����)�������"q�q���ն��+�m�r�yu��M�+����-E����y�e�_Z�!ZK]Y��{�������F��"Tޟ�+H��Aѕ���u)��%��e�&���ϩ����c�i1O���M��8/Z$+s���"�lg����6S���{��S�K^:s�����y�$ӻ6=kKiL�_���:���
4[a�q	5��
�	��Y����b�Cǐ :���f�J�{6��2�}}a;�M&SS�~v�<IF�M�i�T���q�I��o°�f�P�t:|��9�Gؒ�8Q]�:��>�x�@{�1V�5��u[�ʇ�t:4�������n=q��17���`��W��x�r�f� ��mu�������'��U�=��Hs��,��N]�ܡnW��|����x�q�Q�?����щ�R�X�c��;@\k	-��������X:���s����ٯS��f�]�^���R�9�EQ �)?i�6�?"f�������L<	]䂾l�S#q�� ;M��(	� X~�/���<U1}@��E"�)���[l��/O�ꍖ|�l�K��?j�_�+����A����n�����VV0/�I�a��/�%��!�m���1��y����1����ݢ{�yF���4�.L>Q��Mtu'�^����m�+䱏H�}sl[3ܒ��{6 S�͙�����GY!�S���)y�eS�π3����	��ea��Q-H�j=5Ԧ��PA�a�_a�qS����C��jq�YX��C��W/��C�xZ�J��Ɔu1��'��/��J���2���djJmID���S��.����F��CS��s`LB|��[��h�}s�P���0g��L,I]�4撻,�`��k`���]�� �a�6�G$�T�����`�OD�a�m�X�%*c�`U����(��7�RT�!xu0?k,Z��f�;�b��z��׮L�2k��B�Tb�2D���04�����\X@٠_�/X$	w8��dYɪ������rz�����,hM��0|�&y:���_������Z��;��Mh�T+�	a��r~K9�����^�%\Y�w˳�w ��j����=M��Hgb:�[�c���A&��V�ܷ/@�Kc.���7s*��Z��S�ss�;%^�؍Sh���B����;w��G.Ph�٭ @>}/=��^��%�����|�]�a�^\�mOו��ተ�in�
�U�?����/��a��<�h�������_�����I� c�C���*������� 0�Y_jD.����݈����)��Ll�"h�$q�-4�(:��q֝'�`f��9k�yE�;y��qΤ֤V���D%5K �������~CRKJ3!`�v�|�pi=S�b����^�q�3�r��~�=��2Nȹ=�%4q��c��d~H3X��r�!m�"����"�+��(�7��pW,�zƸB�2��	�"W���������%��x!rjB�����4*���)����dC)���G疖t�]���.���Ņ�*�G��y^H�}>kv�Mw�<:��U:Z���ai�d��l�΢�N�M%��2�ɾ~%�5p�uk�n$����K����<�j�R8��C4����'�M��~:͡��{]].��}V�Z�U�s��e���Ji����E�t��1K�Z6V�1��M�/�V��@3�2�%H�)��{��mz��}���" � [�K��]��^!��TPx�W(^85U�Yup����nu���XP�S��My�s��k���$R���U�2��սrM�Q[ٝ��ʀT!�0H�}m;L�;J�OZS;'�����k4seq�����e��{lk�S~�8��%���%���4\L�+`(�Ar=�~��k,�'d�����"l�i"fo�:�߁�pV�}��H]>�\["�����7*�N����R�HV��\|��m�uj�i�n��ȏaL�E���}�� p!D��GmG������^�$_3&�#�R|:�R�f`I�N�e�:�\��JZN*b#q����S����}0��/3���iGv���d5u{7��۽H�Rxi_'����Sy���T:*K�K=�J�����F�x_��^�\	����g�r��4�a[�n�u),�U�Y��Ň*�Ij�(��͛I~��_Ⅼ�_\�������ɓ��II�<*ۃ�
%N��׳ @H�p�������GcL��Nm�pmؿ"L��S�3��Ӥ.K*�9��c�'��*��/WjgI1��w�(��GPݣ�nA�Q�B�@y�2Vg���BO������ib��T���h����=��\�I\m����nuWbq����Bo�d�Űa��qm�����/���R2.�ӊ^�Х>?a�;�&�/�օ��f��Wܶ{�N.���E͔�W*��������RTS"�X坋�����C*�.#b�l�����<��X�f��yyy� �w��J�:VB�����A"iv�U��ei�!�����P9�P�gk��l��gOC�u�bklP.7��_�ɗ��P�G��p��D�47�X�-T���KN�e����;�I˛��JO4�^�%��G��|#���ѲBR����կ�F2x/.f2�	�9p/b�	�����d�Me���kb?j�ȗ�z����x[��%9�P��`-�Qk����qǦ�M�Ȼ�چ�O�����8�Չ�|P]�ٚ����``��٪W�y�S����j�e�GK�@>|��M����4��DC�T�x��C-���A�ɵ�o�>��I��H�F}ŀ�|[v�X�n��s8�u��+5�S?������N�\#���;X���L]�ϪE�6�s�0]�H���!\�H�pRi�&"�������y1<���US%v�G���^��S��l(�X�3���m��c�(��P�IF7�Ax7��~�1�������\[�v8�_��(�n�imm�W%��t�j*�m�j��֖1S�����e��k:!�90:}z�k6]�V�i9t������T�;�&����_>B>Ò�b7����#F�W.�?m��%y�C�-aqyQݸ�ܐF�>�����ȃ����'��c�Ҧ��9��;�RI�x��@g�F�)\N����Q��۠�	"��w/7���[�3<�Hc��`xC��g����I��|)�Eݷ���l7"�Q���юY�+É�=�ԉ�5_����O��W�c�c�z4��hS%� �u�q��9��xS�����H�u���?ӀuN3��h��,x��p|��]&�r;�1�.�o�� ��
A$�pcH��L��k��g6���D�.l�m��o?B�i\� ��R��������<�� �&U�P�p�M�|�d�+��L��N�7���R\V�E�-��|a�Ԏ̬T�����h��~�����ݳ~����#���	ǳa�5� ��u�Q�,�)(�뮿�u�m��6H��v�㤄5�澠rqVRM���ؼ2��U(d�N��Bv-(�Z�PO�U�V�����S����+I��vy�[q�)�yqK�ƒFѯ��I�
�9w)#t"���h�2D�eK"����3��@�e�h�����K�M)�^7�H'A����s����eu�"`���>�"b�I���#tt�7�%�d�$c)co������1�̐IF�cp��3tғŊdv;bc�&���@Z�?D�%o5kF��>>=B �p	s� ]�u�+���%��ub�Pݍ�Z�7�͠����5Ԡ؎=`��I��H:��W���vIi��:R�6��𷅎� �H����h�֟|�Yң���2���Z�<:��T7�]��;�D�����+M�bz<��&t�'2	�|ˣi"5�"��K|�ы�����[F�֛O�9K��"�7�W**�r���r��>B�ߺ��Z�L�Ǫ�l#S�祃��ҏ�0�������l���*�Y�Xb��gr6qY��ӝJ3j����U_'��6)�,�n�uǃԢD�+����[�Y��I�[L�Wz����'>��9I�>�D�n1�-Om(Wb{��ݸj��\7O�M��RC	�g��;��
H HJ�{�
e^!�Ͼw���M�p�ݶ�@~7���s�����><D����!*\
�(���o�Ti���A�8�fu�?=fģbcx�i��}5�����e��
s�"�Nܿ
�_��:��OW�`��j����ڸ�b�5�6NK	�O;i����I���iZ��*Wee��Ģ~E9i��6�E��Q��	Cw�">�
��(�i�#�F��B@��jR�y�]���+[���AL?ώg}A���e)�{y��tw��l�$.�U;,EC�g{o?ƌ���-Jfv2��ń;�mR���m�Hs���rD���9r�k�H�\@�����H��T�L�/��"�Fcx�Ҷ�f�B��Cn*����u�1	˘3x>�Fha�&�t�M��6��<�Vq�X-pG+��;@��6�;`"Fs��Y�;�W�+�2e��.!���}�";"E��NQ��ɜ5f�C�p����D,��xT�K����G��
��\M����m�Fz��ue~?3¤X=#w��H�b�U��nd��1VGI�lu �Q㲖�t�S�Ο�p��d���@�#�>8jS�h`�Cq%?dm�k�P�1���+>��[5�@��p����r����/~Q��%NP[g�!P\$>}rP�E5�AB��O�H
���^9�@�	�i�a9^�H�P����w���}]%}�ߍJx�{�\p'�&r����j�t��Af,����)�q�hP��M��=C�Q�� ����5!����?���ӓ�O����,�P7TM���G	�{�Nc�����M>������JBkc��0�#1�֨��?�=Z%3���ǌ�xM�ஂ�&0,nR�`3Ӊ]Yk�O��L��.�+�VZ��K2)j}����r�@)ز���M��k��~6!�f�#uM&�@��U���hVA��IX^���V:_��M��"���2��4�p:#~�˘|�w��.f�+g��j�G���QeO'�Zؤ	�!2�̶��h<�BOne�h�,��ОQ9�߃�t�xnE�.d�c*A9�/7��f��Z��^�J�4�ږJa��$*9`W8�\XŃ�Dʶ2���M8��YN����?g�z*a�_U�a䉟����\���տ<;���e	��E��*ܡj{�ڦE������Xu���{�:+w8���b�����xP��X�GwOӵ~ms\'�8��3��em�#nhK+��,ƾ�ؠ��t/bb�������(&�3N��j$�/�Q&�K�����w��H8�){T�EW��W���xNx�8�q�6H��	�>������,�t�Vf3Q3bn�P!
�96�6�M}�Ag����h}���l0˳lnv�餔��|.�[�G�(�{��U�hʑ�>���� �8`�#���|]B��WiF����<~y��J�xF�F�O��f��-C���;�Y�% ���p�ր��|�F �m�~���}x��o��<,zD����G,�����MEm�5����k�J��z�v����#�H&�����˷�u!u7�r�͠���8����4��Ϫ�'��p�T�EG�r�k"e��X�E���'&�dҨb
X�c���	������S�T�^O�����
X�X��;�L���_6=K�� �g� H����p�+1��<�	П��5�m�JO" "�%d��h�e������3�수U"A��~:)���P���"�����p���k����N�G�1r�jK%�>��xlJ��̈́,��%�Kn���A����e]p|�j��ÏJ[����(���B(n�Y%(=��τ�6d�lc�j�{!cX�P���@'��.�����\
���/n���Y��m1+گ[lU��(��hJ<��j���GH����{������/uS��m���P,~윬g�h2�Lc�b?�B����H��"tZ��8�P�X_D��l'h_bK�\��t�n bBҿ����R~���82�t����G���1�����j���>ۭl58��H���̶͌e.���|��j�r=~k���mI�x�M�K���z[M�Z����,����z����� ���Jy?���^i[H1�҇2���Db.K%�t9�[�/;k����t�� �h���F��񒈴�+<'Ȩ��������Z�%?9)GNJJ���6"B)��~Ůț�}�X1X�]G�Jӎ|N@8\gW�/���fMt�e(5���N��w5����n�������~WR��n����'\�ܟ�r�vs��;q��X�ٞ^6�Fz1�D������\���n������i	����l���!	�ƪ�qz��u`���=h�"�)�<�L�+@�-{m�=��$  J�W���H5���KQ0rC���zg���Ѐ[O���r���~�G��#(:-Ԁ�ǺE��M��$��r�����~l���>�ɷ1�;��J��U��T}��p��Od*f]�^����ύ���m?�6%E=^[�-�a�<@D㢀V��ɟ�n^��:ީ��`V� �V�´�z�ټ��:�"���T	��Ԃp��E'O�	���}'���ΡA����qgK�l�F�Z��4�q����|| M4/��u9�Ծp� K�tU�q��Ys.آ ~�n�n��p
��������qE��M��ųL[Ō�ѸT�����d�0刍��rD���\�%�
�`Ν�|��y,C�L�(9�ho243���ծ\��"Lt��ҷ�z=־Tk��+{���A|I(��^�#Z��8���mq�����L���FR����K�rR1�K�I-A-� ���A#�Ʈ�j5�e$�܍צ
U/�[������.�Gz�9��dØ����rǴ/AY�5�QV;.~  �bG�i3^ݔ��s��w��mJ瀛���g��@F��0O:Y���.в�Z�����+K����&�XJ0OdZ7���\3x��;�h���au� ��'����c��uϭ	Х1�慖O7�*N ��>�Bw��h�1����sGYc0���Kd�N�sς����m��>��7_�ڭ��D�W�ì~��i���8�B[h[�j­��U�5�o��	e�\Qk��*��*�y$�8��}���)B7+��ٶ|��oig+j��Y��9V���3+m"�Wwy�bTan�����^
B����� Ϙ^P����m����Hڱ&�j���-���B�n�
�b�":|}�>B9h�p�����^��<�mu/GH�kB=F�Z���q0g&l}��C�8Wŏ��>���xki�5l�� h䵚ߏf�%D����p�z��+eI
ͧI
��}D���[�n{q@��=�����R�szy�O��\��A���A�se�����0$;�B[uH����:S�RU�������)���xbv�]�eX�HT�ԕVh�����d�.K�$[�RnQ�J����8'��C|�H=��{�Q�g��� {ʶ^�I6�p=�=>���y״2�g~%���k���Dk�q�:\lV;��g�4"w�:�~��6�gf�J^�Z�&Ma�y�J�9�� T�;mO�(���r�2P�4�#�sH���V�1}�(���h֕��l̑�x�Gn������Z��
�3���Y�q�ܖ;��iU�s�C���{R��3�W}�e��X-�R�����FP	�ѻ,
�@�;�x����P���c��5�^�j��߶�0�~&���ҕ_�wk��v�,���f�S�`�q`�ӜG����(���d���Y�t{�#��Ȼ=����ťJ��*A�@)'s�\+�D�p���/$w�-YL��1%���w�0�+=>K�>�t%CU�yHp��Z���!������K�@�Ӎ�"[!�X����پ?0�"��%�T͏{�f�+2�$�g�81�U�2������S|-�tk�r��bd3Xr�Y��A��o� �luO��<c9��;K�����na+�^V2�R>� '_B����j��kx�M�T[w`喫U�A���T�^��tް�&�4�M@ԍz�#�2�ݨ���?�3�g	�1�f�I�ݘ��Y�>Q��~��C��Wl����q�YGY�7��\-$÷���4f.����V&�hp���X��%�t��c&H����W�����d��V��k�s�u�+��+w�K�g�g�s�f3u��6ߺ�n���fy�X�����ej ��C�R���Ӵ'j�9/7kRd����c��賵���A���\0�k�q��|y���`�+v�A���R@��xc5�8&*�7��$���&d���\'~�_����_\694`1C�B�i����w�>	ͱ�����.	
n�m�,�A�l�BȮd�~XIO+�W��#ԟ^�����'~� ���;���[2��T5w��ĕ�o�{�,�_����fl��"v#��!��l�[�6�W��=�H�J���I���-��g{\(K`e������Y��,��Ѭ�;
ўwV(�.�o]�S����A�K�d� D=ju���Vd2�+�AE�+��"9��G|�����]KY[͂z裏�৯u�y�����vb9�ԭN�6̼��G+z>�T(.1]\K�
[��������^m���	_���