��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG�V�����3͠l!I>v��c������{�^J�ڸ���V��P���l���#���Z�FMf�P��k��u��.�W:�l�Ԩ�l\�fP��+����]y ������K0�DѱT���*p��o<]��M;r�J]2OKS<�2�'u�/�+f��y|m�E�\7̈�O� �ͼ��>��L8��b��[�8?tw���Pώ����>�~D�0�X��c��g{R�L��.}x{M�T����㡃$)ѱ��������;��b�M`�x��r��1���_ʲd�P?��kM��ڀK���1r���%b\�i��i>x?|ҕW��7��vŁA�f#�#����?ac%����wWc���`��?x���Pұʐ�o[0��i�b��%�b�@�,)|�I	�%@C��s��YY��~�u�'/�FS<�!��5l�B�#d�Wc2E$A�
�\��e��q|��	���=�����mi����Qz$7��-�d��[K�$�Gb@��@����S(w�"�Y0Q�IV-jB��6������~���p�����3l&)�5�������jOt�3����ƫR�&U�PZ���ү�~2�O<R?��=.��c����.E��+�8�ѕ|&��2��_��.1��H�4,�A~�|'��p�%x��.ʎ� �Sn"D��b��=	�ϻ��}�Z���}5�F�;��)80��� �luX������e `��3��@2�y���ȼ��BΓ�����R�B�')��J�x���ٖ��Ӆ���#�$�%#˵H&��u7��B� C_���Q�>z�&�Ѝ��Eǯ`;�-�v_,��*8sB�5��t
���D��q2z��R2zV1Y<�f<���6�iK�b�%�5on�0o�b�'�
K��<:[]WWhO�X|-�Bwm�'�Ul���!�iZܷ��GU������_�%.Jq/zvB�)�u���Tf��k)z��1�������jtV��[]��ޛ�{�&VK-�����Ƹ�<���}���
�ɓ��~�!@�qD��Qז�<&.Б^��mhp�����e$�*oi�]�s�X��	�7=����S�����!�*��F-�ɬ��ٶ��R��+91	���X)��~���o�9kR���c �*�-?[���1��_��R}g�������dFƲ�o\J�MH�}��ԉ����4�	��h"��ٝ�;��Ө��	�ꁰ��dX�to�J_��.�.%�r�`�$�{2�o���Q�Ю�QU��w�@s�.���V15�۫�f7\�BdT�	��S��Ȋ,Ϯ��'nz�_��+r�D�	���Ho|H�Y|D��}�9�Z�3���3	S�YP���{�v�>��1����v���Jн�ŮAP�;��l�0za;tE׌�|FD�v��i��b���@���
��N҄cp����*������5�M���C��='s�"�
#�Ћy�6�L;�LMmϨ�,���G08t(Z���Y�m���_JLrvE]�R�gt�B����J��Ij�x��᫶J�X����H9V�y⹁.�LX��E뱩w�l�uT�**�Y��G�a�(w��(T��o���?6 �*�ͽ�Ւ��dA?5p���0����B~�����Vr	�i�q-{�E��y�� O#T6MA�҇������j�'�;��U�����S�u'%-+E�"f7E3`�ΏP�o�i��B���m	�֨�Q���v�(�K2��4+� v�k��;'�A�]�*!��\��̻$��w��Ē�S�G��dY��)c�!xx���^���cFd���j�:�[�?�lZckMm���ޔ-l� pf�;a���4x�q(��c�yۣ�FR�R������G]��=�3��X�wH��OnB�M-G���d�_��{����1�OD3!�fc����}=�]���fW�����u�@^�+B�b��<s�ꓐ@[��ۅ�N�G*�������M���`�Eν�t	��f�a}��sP��W�*t�{Jvc�`˻DW�gOb0C��	.�H|}iF_�(�Ϙ�G� ��Q����u�9��e����f��Q��� 2%pJ�8R�"�,9FR�f�����<�3hՊ:I�Π$�O8G����y�'�*Go�z�rU��I�U��#̺:$@� �L�h�}�}f��`�G4�`7�x���v��X�,
l�s����L�Z�uO�0$����ŀo��$&34T���#L2����׸I��X�	�t��rFۇ@n;�����9=�x<j7��i'`�"�"7�q�qaŀ�,,�d�Q���7G9��Cr�������k�	J9mFR&�A/���&�������$T_�)���ٞ���_��� ��$<��&����}ӃB�L�����TK����;�~�J�Ђ[��c�Ǔ�ڶ�&�*�0�cD�,�ұ�z�pl�ITy݅���S=}����W���Λą�HT�b�C�I#�L%��2$C/�'��F�<N;j�&٫g�"��C�h�D�����~��%��Y�+���������Ǻ���3�TVư�pQ�Mz�R�lG�	�M`�[}-�Y�d4Q�'$"�k��Y�}���X?�7J�z���;�!�e.w��.y'���O�L��߈7JC�*�ޑ���H,2C������Z�.��&��O�XP��=mi���K��<]9=��-���c&�&�2���l������`�Pu�\�/�*v�����bAzz55,/��O����HW ��|0���?���3�����~�cWҭ�Mcd	X_{,s��K���*����C1�d���|��@1��S�#!�!8���i Fr��"�O�����)\��c 7YI>������s�A�P���D#�S��9�`mj8�l�rن��(Ƈɴ�C����.�7�
���öS��.i7���-uc�oȋy��U�����6�-���h���$h�$y�.���I"�c��Y\�Fp��;�%�G���;[tz����B<W����2��J��a�y����*8䔒8��߹U)�H�'�IsX˥�w��?"]x�0����֙{�r�)���*>��UF8�~����:^�J±�o��Y��Q�1p<R�V���Y+ⓨjv3�?����fn��ו
I����*:s ��}0ؘ����Ϊ�[����W�7Ť�QC�����l�݈�~g��ҷ��"lF��e]�t��f�oY3EAX�0�-/��C̵�V��Ԍ�qUd��
i����)��*p��q�-���)1~:�&���[Q!=��}�h�V���� �QK���nǸ�aK��)�_*!d� �ˡ��Ǒ&�	yZ^�a�|��/���^�}܉=�2Pltcg�;+��\E�B�z7f	x���V�.�#���lot�Z�o{'��,7+�h��B�]Xv�ͫ7���^�{ذ����ɞ���\���X��#u�J����D�~(X�č�	�=�H{c�����GEG?�L�์�u� �P	�򪈧��6_�o���#ڟ�����|~����N}J�^B�c��pD��tIE<E��Z�f���&�dˌ_U8�y���E����A���?Z9x��S���Z��B���1;ٗ$?���<��~H̝z��ldk�]�-�R���^� �r�LP4F�d��77��S8[n.(G2�O
�
	G��#l���|!��3���]SZ��Rk�S$��[�Η��6U��1@oϧ��]*�eX��j:e�3�>�Ŗ_˒��OZ�b��i$�>�Z�j���yզy}\%���L�X�խ6>�
v6L�B���9+��LC��"�Ȃ�ǅՁw��s��x���Թ�c��s���5�C�ηx��~߈@�)/���Q_l1���� �s�TZ����t�HH��Y��F~�s	8?��v��;z����s���#��.Я��I����H6��B�(8���2ߤx(%�\���9L��su�Q��q��a{l<�4a:;�%�&Wno,_w.��%��'k�&ҫ�r�͇��?"�h36�����HZ���9�b��1-9�e%f����ǚI1�����c��@�.�Urӿ�3�4��r�;��e.�WM��x(����O$�0%���2!t��ڰ��:i� ���x��0��|�oP���D�Lp��m�� �hDt֡b��7}��º��x��0�[,��,5s~�o�˚�H��{��;�~�{�ש����?
(ym*�/���X�S0�M��8�9/�2�đB���j����O���6CFb	+�ȁ��� j&7��09:��>�Ț��X������BB"K<�ɨ�3F�k;�f97bBcU�B�GJ����������o+�=s[��i��i��m/fV��G�r�&i}�}p�]��3�[װ��K`�矀t� ��M�,[r?>ʾAg�B��FT�,�U�JHV	p=rH���_�7	
��z2����W��bt�>i��Ӫ�D���p:� %�C����'�q�\T��]|%r}D����=�|n��Ȇ*=E��c>Jq����L��@��|d��Ч�(�?˦����Ɉ��A�{� ��ġ~�o�3[���b�N��$�7 �\�U��0#��*��L�s"R"3��^�c�k�`�	�.�ոJ�����Lr]�q<�s����I�; ǒ�����&X��a�f1R0f-A�\<U��7���u�o��^m�2���cD�V�wG�)3��d'�g�V�S���
yQ�]
�Eh�(GT�f���XO
)i�*��";p��4B��H�
���!"�2��zAW^VV��+ײ2�����OwJl���&�@/�
��xO�{��������Ѿ�Xk8����}��f�;�B�f-;�e�e���&��y����+tLS6�u���қS_^6C�#y���HF��KB�T M˞�y۷��tu�5��/���F(��6��Y�POy#lS���t�G������pHM��J"I�e��9r���I�91&�/	�����YC�'8�3Ҁ�F�K�`J�.��-��N��v�Oe��9�m����zW�.�f�wq��<f8����5'!�iH����װZ8ک䍖