// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
bNuX3sx5dfzWrh2DRhepHxAaQbPo2Oosk4oSEqYbl//rkahWpJbVYUGA33J+Vtw7GHcz3IBlxqd9
syZZAaXHhkBdmvargqVe+w3usBCrhs+K86DBBocqK2/LJtrA9r+/SgFUilRwZMV1RReLQ4bMg493
z0MRveify4lqEoaYWcanW0Uo4WuhHqKKUWwipF8jvtHb3OQkvzhymcsPlYKRlsTseL0Db43OygVg
Fq8uvKhZ+o19+Jdxz+oA2JDafmcF/syMuxX54Vzx4duKLMRvUALRhMJ0MPBQLf6b/IGsx/RhEIk/
cVVjUVsiv4lLXXwL6rEWdyLVUX1Hqq82ehcNhw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 33136)
HGpjilmY8diTl77Nm3L+KItn+/01rNq5UtZWfSPiOLPBfO03y/PFZ1kpbPO2XMUBpseq1TUkJkd/
qnH6GJHOsagpVAjggOXib031oMGRh9CRmcsvyZot5QGRX+cp1se+yGbRl+QAYsuHlooOR6E4yM2q
zHX4OIEYPqESTJu79vYM6QPBQaNwAW/fnvKEr0d10nSqIedj84h25JNocXLaZC3uUAlJLtsW+/xX
3KD5HhBT3b/Tju5q55qtA2kV1H7DO+GOnpf2gaY/ygNg+KwmJ8eRRscRA74qQK9T2LKHDfT9YFB0
LrVcG2N2JLsK7a28j92FNtL433gAHg1+R3CY3KnOZS0juxbYhn9SLr3X4BThjdayexozihMl6bPu
Wz1KehioEKBQdB3xgKzP/oFhSEKSkloPZqAk2A/1nt/Eiwsiz0OVJX/oyCkRWLZNrt3eiZRuAhzu
j8IMGFEPSF3hSpxmJ6tWA2z0AXl4ZFcO+G7oAbzk5vAZNFM9egB2WNFALhX+5gbOvrnLRMsejOGn
UE6L6Qtx0Q7sTl3c5n7N6occR79W1P5O20umVaHfLG2e6XeRYOEpS7+A55Wf4PpfYJEVyazZRa4I
hRfI0VrRA5XdvD7YtgVkRpkxY3+ZilKB6GrMrlZV/mm8MNqw75bH7c/jXZwABS3ZSwLqgnhibSiW
KWnsM0jby270w72ln01hVsKjc9ms0m7D2vofs2/L2XzTJswRDj6cP4ImwoBaH9gB2Yr+z5Rb34LL
0d8/3ltcaD5sjwpNmyDo7jgyE6LkPLGWsfe4BNYqnCKLf4IXgin/oSW7795B9IukmFXQG7xA/i/+
HWiUnNQtM+AqTTUxiL07eAhPYmW4n9DnJpORbdcaW6UZ0VNlYUEw0S29wZEAvmOA6i7P88axxXP6
fdCR2aFOOVOibxWO9wkxyw6EPHRMFvpFU1bMXYNsUomkw13dWx0TLrySdX6elxNjq7NwnheTWf0e
a9cPxcK/fcsLUQkHyuKnMmuPrzJhSi+zSo89eWWlYnRZFYde/LxVBkMc7ULVTbhHxe6mpJdUZsqW
zJzKQ9BMZkjv8NyCqiRzcUaOu4hL2wRW+o+AungXU7Sd5z/TyRvTwuqxC7ekpHng1q+tP5eYsBX+
AMCsRKyAFFd1pYXzx3GLx8tAY91G0aqrhOhpwRjHp5O3fkRHbGJ88FrID6DtknxDmIuWQ8W3cLgx
FudEhoUOCY5KkBEanVHUf3ioEk4Cdr/KOtsO2IfocMW2JdV02ORJfaNUJTP2itH34c7xUKvPG/iT
Z67Q7ZTiaIWDCOsrzKetEE8Fwr6gfx8HescwjuIlSrV1Lgvy5r44ED957Pa17DkJKoJD94moaoRs
xsO32kYYkdGikqub1E1A5KoihMNjobFICMG4Xt8P+I5I1PvymhandzFlRXV4xEkCOD4qqE3wk1ll
aAMWIfwegRREz3g/8p5RrQJv1kJypiaePELuIgsORcPyEOxUdE4hwRkrLSnCicfdSRw6feg2+6U1
+wfPP8czuSFiKs1+VJLu8OPCNLb7eGNzWmukxeVgFRgFsA3GVWH8wA9H1jo+J5bHFTN9T65Li4gX
Sepk/KLZhQwWX2RhQ81S4qQUx7A4j+h744SnM7LeC2ckJnBbiNEWVsBezuIRAq0anSqIMi+I6TGF
kjTy99su7N/oTyiMZ1qSz59hzGpFIseKXK2o6Jd+ry+/UEMN6EZN8ERqdVcG0R8iAEcaOKs8++NR
tO5ccpvfQc8KHxfnzqmlzuJg4+awdErJCswQpsReRHc4BMxLG/uB2vMfTZ5Fevo/lRw24q4sYtP3
7+IhxsHEF1EVvQjEj2ndcJnOD5u/jEH7oHKwV3JsfCeUHwkXhzoQoDkOyCg6JXNaDQ2j0GgtaWss
IuUiFi56U751dWRZgoBmVtwL7/w8uK0LddqikpsGIkmxMEMJ9BlXR37wkJAeMn25FbPEEaezpha+
5oO9zdbhQttO2IVWmQ9tZSGLxCcVi9Q3OJzmSW+OUqbbCKlt+2xh/t+Va0ZhDLORxLe1lGNpMWLn
K0ZTA9ypNZZb9GKuNvIGpbFqEtMzYt2psCrAt35NaLNSnNlY/I0bscaZ9kiQ4uFgEAW6u2KFXu/L
ie8gKUtUgA5cuPikOCWr0GnUcAKrPmcy2JvqrmGchKrupYkgeeCtMhhq88APXAqVfEMUCHb4Q3g6
KBBkBYJTywMqb+RtoWcsbGk/FKHD1KTw+91wEN6XLAPkYpLpzmzsiyjnowaKhIWJ/Zflo4dIDAZm
E4f9X6gvrUUbgTThzoKiFGl6AZ0eP7v/niuvokSoeEwCux/giDeNuDCIP+otvom1VISKFCYzepmb
Ns+PiyScBWRWM++8votE+EFhWDR0x7Hy8kMVKDZpquGMOs5r3UxYDsV77wzAOa4qwfQGe7tMCv7b
31wGjY9GScVJ36K7BjTzwupNwLlnLmGIprCn263szg1DWkS5dVB94FYhQRJ98spY9M8Y4BOF595n
P1KzRcyAbZy1oeafq5iHWOZy1/A92Xyb0nNG3orJuc+ewU1bbda2/hXz/CPuPu7p4i1fSO4VYyoi
39NK0RPz+D3zRSnA/b8BJ9TtoLASsvhHR4l1f55jMVo972eH3JUDPId65XmvjYWXWiyywv09VXDY
lFZGeHAJt7fa9MTEZlnlwoRPNSn7xmI9CHSS3J0Dv27BCOt8labzZ6Q6mlQyMLcUP5bAgw/0+Cqr
yAVuQNzLHrPi16qkHcRymcbRxI8Bw4KmI00vPRTJZv706rd+rfad3498YrKQyYpE89UpEVtQqHgm
jTfubJyizDj07lIzNHPuSjIXy9fMyXpHH8DBbE1YotLV/u3Hd06Go9ka2M8rWcAI6JcXZuyUjcRP
NgkUqThZFK4xQOqLqdzwa1YuYX8nx0ig5AxiCK+2KW2hU5jlkSN1YaERrb1ZsHFbCDhWBfRMBc3A
vFYT72MoLfBGFGePVSMy7qZhN4dzJ1nFsY3YER7zLoysjAhCU+RmjheAh/M64faa71ypWOgfHVUW
JLnwlt1oym6OA1Gd6TZx7bhPY6vEhZladmjdT+CiMGH+WgBP88e055fEo067lxaBU0pZFWO6wva4
fZ9ka098VrW5D6cPLtmRj8mE+EHAVsiPpFcbZVxzMjWfSz1D2S68PQkJGG9pDQMg0P0lNGuFcgZZ
rjF5iLbFvRqYoNSBn5BQqOiFll0vOyrsh39afikhGxlFHzzQ5ELn3ItRRzeQHI4GFj5Xy2P5UH1c
QSd+LqwXNlMOvuO91jLIArn61r5yTyh/D4P3qYe/QuKRGb36hOaKkfUKtpn8dxxHSoAp5cnU4E5w
oa2HVl3sbseOWw19W56Wv6lgHVJXdtdxD5XTLAH30z53ZVLdzvDSsaypCv8y92sG29wYq/cAJalV
CScZ7K4lYwSABh7sZwR+BpwuyPklCVXUtnvPjzEB7irFYxcgehCFKk4N3Hq6H79ks0bG6qzJiTCO
zlAy1F/YiReQMOVqcN2DDAVdIrso0sRDusPQYNaEQyUum89bGplmfQet/aTbqAYSQO6S6hj+jwFZ
5ox+Ae/URtfSQnNF2zrxQCAFa+JwLKkEBLUubvbtXMBCdf9Ej2QAkCs8RzayW/pE5Uvt4D538I2r
VSA5obAdD/BNnzh82XbuWuce+eAB8ZxcxzhooiE5HXN4gNbW1Iqxldaj42/5EQsCpT6U6xSS5db6
8RdWomQo/BaQ+b4YPylJnvPV8eQixuxEmAMYPCyb+nKHde5nHmqybm/d2I82bZ53Ghj++y8NuFqu
9KfFrQ7W+nLY4BFM7GXcD+496vmjwr3csrVf9+sHPqfJpzRXgB8azscGJ4P1ph+p6qA/3sfvWtIl
6X4AmdJyqGLpb1spPPRKFyysMMZHQ0KvY5dPc++K37XTZyws2hOmLUdiRzHigmMVRxNLM0hjv1Wx
ozcCUKo3yfJVBTOs9bw6jUlXQi62vKf7cTFUEaFCuIq3M8HAcKTpNc17uoxRj+gRbXLojehSob6n
UIoXDl361lahzqjzdvw+TYHtEjCS1CmBezeSbsQ5NoIbaS3wqwU3UqiifoUVmo8Lp9ALkHaU8ZIS
vEcU+KG6t9ARBqMLHbAsh7CqxVgmTEl4dURqxj3M3vgo42TjvZnnoa9/YKm9ILA6PFXjyN5LSFBd
NFmYhJ7H9me1GttjWWexRFd8hKKhXwDHVRM2ZauRiECZzyxT+Uim2zTGDpQ8AfIOlkrqLQjEqGTf
XVfsfvLqSPU2i0/f9YRiDDBArOeWjtdzs0F0GF5vT+NY2LYKl3+G6YKFkReb52bgVIL7f32SyFIi
ZcVonKrw9QKMWGAFzYg7vT7ltoNBjxDVjOnzfdUYupmoolSdM9R7STvYYrIHphDRGlvmASm5UNHQ
MhuDAce39IgiwWF5z5w0qsLPUGxKrTDe1QjI1sbC+h78ikQxy/Wygo/tVBBGBfVeme4PNfCP8yvX
EuNDr5/cNHbTrMC5RL/G7JLe46HToPNhrbq9/XrPBBvp1oB7nlWiXcxeFTGOQNtzUDz9lCaJm0++
IY0qFdtX/opNRV4XfNK0eADwdtLorKiX6IghDsLDJz1LSK6dmuNqKD8E1CVhEDnQeuPCgwnWk5I2
y0ASp2a3TPIEpCW31luqRnra/zBogBPXUW73vUul4iYE31oDvQOtUqOql51eLsNAxwBrM1U8dpGa
t6ojIXEG5qR600m9JZ2pv15+7mp5rW1oNkJIgL68vhH11blm7O4bQpql+WkiLgC7z3P/xprMOIwu
0JPzMT9wz8Zqyv79RnKrctIy2m2yfoaIZo4DRxZeoszPVnG9II/vqH+iGNSpHXxP/wi/QRCZ2ZVV
Nu+hPIWwNqgUUIsAdm/pw1UAmLlKzMNmue6+bB0JE1UH2Vo5n/TgmBecnSEp87/j/4zAtqEqOUBK
8Ey29hJAY0UvEkZqSu4OS6w+UmAS8yf3nPk2hzXZwXAqGSSSEA9DlwKTvL+NzqmDhbXhxOprLH9n
vpQb9DZPo/7rDgtFIG3ez+95mJh9CWr4fmFL5qMjxyyaTziVIigPNQ1KtfArWLRKX6imPjBGJRc1
Ubw7Qxj2t4mnwnVUKVby9ZdToD1Fo4CxD6uiX6QmYOgAXQcPxgaydg8YUSqDNOd//xvCu55UtSgB
iVmwlhwE+6mcKjZDOML0sy1tJFzI6FU1pqYZ5rmGTSSQYnnsimfBBPupingXAzc1QepoYmhfGH0G
GNvtP8K616k06AsFc+NqOUgYgQ2jumvxZtnZt9760VU0mkld/JQZX+81TCv1Az8LRfdXXsAGYf+8
uppvdj0Wj9NH0optp7Z/Hc/0aGaTsKZvhOJ7wiydl7Fo5anK9bCBd20zppD+vFbF7GFkFM2W/sRM
z7pLX50Jt8zBv6ZzxsiIQ2HzLOIFHuHVgUfgGfWJ2BSKTTeVXnKtdfW0rnunRo8OAjZxQWB/LKXH
JxM9krxhMaYL1+LQAu+yz3qvhtcZlN0yfPkSLsVfJDq9B7d3bB+0ZXHFNNSzxirAsuw+FF3r0924
QlvT6XuCTwotMgzKhgLiebwOtV4ViVckIooEmQ7vQ1Z9/gN46tEDTcp/qBLtw55GR7mU86mMsul9
rscHwuImA603w3GPm60mTMSsHBBnOWmjjYpH9hcwVgUcT3BNc41BNnXawljPHQlvB6k0aymsbpX6
toBnf+qcHgr7efOmMC3VqBm9bSU7C7ew8QOX7SS0M9h+1qq/R1TBdPp1LE4nF2eKAOTsZfTheTJj
ng/V5kRcRaEPdxqbwjwWuiZ7vLGlO2K7sUth73Ti31APFO3iKGVz+JsJRFxoFt0FFnmmM2KQgT2D
s8Hg7NYF9u2aIZeKea7/U/0qUE+cGzlEcILVibGj0WPW0FPKz18fc3HsPTAE2zHwV8CxaQhoTTKE
kujTZxLEk9OplyFGv8lv9r1L+E7F6VPNM6E9MgqfXx+atbwTmoPxFJiXS6R6m6KbEWBPje1T4HmX
AEj8uDgYDQZRqurxr+wXq+ntg3KaI1txqJdFyM4su/v3wyygIImGovQf1RCwqsdJO0VmBaTuD3oQ
KnhEmb3MaYXPIVvBZUDiPSpSYyDns47BPhklaHPWbGCd3kNgqC2X3GRQTd2kom/knCsR/7zM22yu
1tdM+jQo4QubNfIfXA0f6uAlIxswaifUMgyKPfQEe/a5V9WuG5AToA4VaOrvVWSnDarV995vAB9f
fUYt4Lod1Dh0lljDG7q4CxrwIhsjOO7lLVWO/DwLlXOncavchWqFTPDp8L0H0z4ddlRzi5S2nI+J
9VUJcXF38n0gtla8GleWdeqE1OLLLrDYnH8gda085dsq2wy2LgRhI3lAz4ZDpYQlkurIMf7lXNNL
Hua4CJM8lOT2Hs4HVkNYYf/Xbvryzt9Th2hwU2WM1bsvx+0MjnLECTJ4U+LE4swcG08TymQ77Cfo
WCws2/GRE55mvIapP9NSzyM7pKuPajw9MT8U8pt0NIm8Vbro3qU/D3PXXgJ5XgkgggxZvVQKSYMU
ZVTbS/jDpEUU5xH0kqavORgYIetB/8qqFPxGqQ1wrpUe3cOj40NRa+yj2AePiLgRwZKyA6jombUr
HYOpO2kgLUYceX7JnlsM6HkmU0YhBL9M31lqNwJ2Rilk89RYOfazHf4w77mKbWLlt9avI3nin6gQ
CRbLWVnlwLf/uFcsDydlYQHjDR54+nRi0t4qcxYQwkzyut38LUsSfHveWWYrd/+p8VxpxQ/8CW+i
wAaBVhmvQxVHnwjfp/osXyYjwAAfCgfsgPGRzdxFLu8XKUT56hX2TxcmgojJMk2MXQNZEYf5NTJL
sRDetZNL+JPebW4r1S7GYDUe/dg3Nd7OESzfl4WzA8Pe/7bArytt4YJWH7h5+w/bjWfjN3F5caMK
IJ0UEZcX2EZQsgG9dMIHljXsnX8Lt03Ht4uVogUlIfuM4o7DSrAZS7xwVfGgb6aFvXH58QaX+b3y
dMyAiRha799qkphIQeu5lRqd8R+prO2OR8DY7ApQJKzrViyAFiikM/GNMapZ2eDGhab+pNDGUxX4
M2nTeXenIvNWfMfbTjm3DNQT9Oa2oz4xzthOExYmwNhrgDJQ/h2+Y1CRNrISpWcmfw15pliGbamM
+15Ub2k9YIAkU/DuXodEJf/UPmo4JVpLTxz+e5tSLEKyy8gyOB1O0kJBZoY/uFAX6+jl7tx9SEPX
/e2aU2Q4Aso1utMCKiAQmbFtJmKiJ+paEN7MYSduiYyqUcI4E2lTcePahv4skSryZs3YkgtGFzme
aXaLql+AQi7O0Mh6df3WR1YrOecKJRW4TD0hu58lOVAp4dNJq8GEnEw5VkXGjvXWC7kxwmTfvvJ0
qicxOJbuWqEEz9kSzahnWNATt0pMiqDlbgeU6NdujtkgQfOJ9PLzXi8UPmIud2VuIs3nn29hsfs5
qQKckRI6aXjxAulseJjOOUrG+r8fVCOWAinkh4O5SghpHhq/v4f+Z/CN+RDNPdANMW0W+xL6cBD+
hcMvZ8ywMWXqUfcNZbsriNHbkBxSbRDV0wfIpLbTpsgS9AEGnbKL/k1gQhFPpc7J1UPAywRVwtLE
PKUuUD8UDDdipxXbttl+IoN96IrBWdkwIy94Kj0vd97HXwxkUc5I6GUIoxNAQZnJ37ySwGM/sS1l
WNEeDhTuWB7ykZVC5LLRYT1wPoUcdxFiY/ARphtsYX5cDqxMqGxwl5Y9LVbORr8hw5tYzjVMZScK
5Gk7FqicuP+9fJkXbyLPqpKXf6+SlrJCsTOL/94LiT9ebBlhQA4A5n1oxr7N2RfKkfe9xPQ9nfkd
Oggd8SB6jxrDEy/S/JntIgb8jlt78krs6ezpC85qojK6Rv3ArYMD1VcUWtmDYsVuJNgWeszzQFqo
1DaN66J4oeN/NWAaCpv5GPzbjELB3uq3sLjY1Eip6d9nH5/vVGTlbJyklEF1x9+58UvQUDe1BVPf
0c3A6+eEGGOdSQrPYtnRPCpkwJ633thk+CtEgXAoHnkyhNy8EY5dRGgfkVAifA9yVu/lsa+2iLfq
sdD0+HMtCHmUZiMgTaiB0gg1ChAdk0Qnsx5rad45anB+xhweNaAwCcWvWmzh1HkT5voCwSvDEzgf
AglQygfkeHmCvOpfFOAIeD/EetEaNzz52V1K3FBENIu3AyMNdA9CytehGJ3Gh8maqmuwZVYc713p
cijOmWzM3lo9ZA0KOGjHihUzMyMYKltlUbKa1GIdBTQAAhCXbWE43o1II7ND0k3uDsJImlr5MpvH
5l+WBC04v9FqtofZIbe18jlCgFECH9Bq4Xm5MLMk5XVW7Er3oS5l41ar2eZh2gydSI0ETbNXpYPX
ViH/owjA+sVeC7zSISMevl6inakJkdFTQ7AiX7knA3lNcKrk/L8Pta3yigJhkcSiwMaIWRQGvRK1
xkEwskqKrP8AKkMwu8lqs9RJ4URr1SZQsLn4bOe3CbJwUz/tYue4Y/oQ+wGIWmyQgLZ2jN0gbClP
JikR/uQx4a6KHWrBQc8AXnDodaX8TM8ptfSqx4U37m6k9zRBsJo0Z7SdGaKxj88YZhuVtDJYk0s0
JbhHG5WrdXyMliy8P1xrm0fBaMVWNz401SAKyHNphqq0+7VLYh4f8tDXfdI/PKEJ1fefNS79/56B
othIzsUIX1VC3tkTUmpGiuBIZAtKKmqRcBPICUlBtMtgYk3d6Bv4gMQGIxK1+aoVJ3YrNoYDQDuV
rN2sapLFPHJUTvZK4HIwqZ8rezcmD5cpN9sZsk8thanCK9lI27KJdNcnjBNCLaoM+vEefj+6NIcn
/IZokuc+nAJsAHQYm+3rIN7g1gbAlGAWrWvC8SvHDDk133UOTmRX8US1OnSArLoZLH/FuJKupD9j
DdnA1l63VhA/IPafD5wtoVnJR1V9YQSfxsf/gqGuYHpeSFFOWIWCvI/Sq1HIfxoE/F2weC4NGivv
sZ80u67BqpSQJBhoWyO7w1cRbUVn7k6UFdiyp+L4Xrpu6r03Gm9RQioDfCC8LpCY3QK9WdnvxwzS
H8/HcJYS9H+0s/TKs6lNfeAloU1wJJCzMVpD5z2z4XRDeU0dhxt617Fp97z6kLSx5/CAOecq9KSs
NRl7aj+IU6fqAajjcBQH/wyv8YTW1FwHLUA5feCyNqDnsMQMED3fDw9lOIhFiBzyETOrVF16oHH/
BNKDJyeSB0LNfEJFZHFVazOAeXfV5z2ckpqGc/jO9aOb8c+joUaEZo6YUYnKTzWCGaMjWRMLcNR2
BZgHCpL6a+wjxF/GlbRuRXBTGFErjWhkGZQkE7YrtekeJjV1d/CUG6ugjqOtsPvXiFQ8F8YdPZs8
XDnBrTpvE+wBqO5Y2hlF4l//amIbUGeucKJHO/h73fmfotE054P5MWUoqNC/lbB0wRiki+nM+FWa
E+l2jgrOzXUm3HYRaIvjRnOR2/PSRPDgOxOaVlXAH4iD/R2ErHtqw2+sJqgBUlTBdHCXONx1bKPx
3SgOB0YDoEomiWDwDivr1G6swiHGSVAlqwp5lc2prEV0RwNaifbY1JsipGvqRt06z2s6g81ly07X
6KFZoOnskIvFiHzPiIGrjeJYwXAV2T8xRtDcLJMxnocCmdaUexpoy78aO/oax3lrcKSC9sYgzTvc
ixwNQ/ak0F0CaEFfAE3W3smlvsAZjaITyMJHOAIquh1qCuFOHio4Dr5HwP/pUPHTNGToQ7NleNLp
DYomrNMMzFvOP5wwdy5SqkKhEzcTWScv7IiOyixjo4s0e0rhe47hxATmP8QaoIhjSXBl7pbFESQ4
YVTSetzmRKi7ENli07KoDARvWD9AyQVhsIXwkwPQvq4MoxIp3Kwu5WlLMSXwnVmj/tpCkF5H/BQb
l20/6UBPDkPvaDK3p/foqNHh52po9unczSPkdZ6NrSiSdM5WuAruv9ltUnCjwhPFi7T4AutlEpE6
dhqwnIJ3vBoW0GmDbKt5utExj839EMWBqZb2RXybeTlUk6j2BZFAkAdHp/ZHPOK3Mizs3APJsFj4
nRgrJwj9c9CgYUEC6njCqQ8NgOaR3NXIQ4O2/A+tHDaXtZRsTYNRudqoCC8oBc9/tgJ2O00Maq4n
P2QRNWjgBTNcFFmCxwxC9Aiv3qsmCERZgfKhadWmfAd5tAoy3VlCP2TKtIgnQuTu3ZoCDVyG8z+Y
Y/71LUOdL3iYu09+Xeh8KlBcp7PDouWB9z+jwA4Jzt4UsaJXBl4e7p2GJkow67JOQsURvuwZr8yp
au2NBaqEw8GheEPoc8a9+4VBbnbgYhXcn6sx8mGP2ZPRn+32Me1Fk4AQHzAAmnALYUIjOCqXOV94
HrsLD/8sqHN7ERsBWH+P9BhSP8ITvjWAxR/LK6WudaOAe9QL/35EZcdyxRYnTWLmv8ZnXEtvIOnL
c4GOuDkx7Uh1dlqlC3tuR3LMVnLqpicDSUCOhK+zipogtRsCD3ba+4N8a2SVGWqwuS5uX7RNacnq
nM5GblDVWS5eQ792zbW2WqgPnwxTXISZfi77BmC5i3Tz4klQJYN70oc3FMym9mhnMcK9Y/eqwA4M
u/ePR9KJdtMnc66aGwLVJxKs2wCXwyPu6bO0yAfmgixhcKohlg+6rDxC3jWqEOrzByC8p/sWtT3c
MebsGPULbMQsx/VVHZo3CgNb6caHCoO3tZXayb3ZC66+ueIod3ZOu1L8UYBhSmq1w9Fjg9Xyivdh
VVsJmiqVBFhzRp4CH1i9qjcNzU8fO2QeQQ+d8W9DxgRFUyK31Q7bcwuJ8NN/ksix8ft/V4v6i67Q
yTCv3qk+9Dlr6OoxRHbPHEPt2Kcm0uteYIeiEd4SzguBE2DSnHAGemm8A9TVbXPAZIvZZSB0Q37m
MFifQaYke8YXgi00W1ka2G7Svff7zffm5xrFkUiY+/cQCvS7yDy0Si59FPee94HA9fiDkYHgtEbZ
Fa0K28tRUnhB6PaBfFKrqYWqpWIrfE5tHYTUf0IxOzOBqvq6Gu7hThl87wOOjANia/5I4i0JXIuo
p+OMjQ/rwhe1PR/9g6uLS5iikE1bUYEhqkVwwyfM3oWfPpRg1I7KWOrGi03ynecpJCSCBUUdaqi+
aZeKjzqSUo6u+IB7bBnzomkcOxa8u7WpTJEa5oKyTlDLQrlLDQYfKgcB8m4XGl4gOdVoAheZ6fzx
kLn0Wdy6sKRP1O0PAuyqKEzaVjSUZu5nPDrqUIsQTYkijjuvqmu7TMJcwDGN/M8rf9zzWERMUeoQ
JaPCHWP2LUayxV7LWWWPWB7fI7kxTXRDsX0eYa7gIfCHf6yH04nmBfdsM8NNrS3RMEreLKj5M3O2
+wj7Xfds0UiHHw2Oz/Ysf7qlj37AATivYRMo65qZHIVL+AqIbpG4arCMuzazRizi43295XXA+Lhc
caK+CpabfbEXFkqLwcChFplMZIlk96ztK3QV4rlIrlH2+FbXnMcXE3MFljlkduMvEP8esUhe1fbQ
hI6PbUnhvUSeDc0Ow+xZsWP/f3sG4EnM1GV40ivgBds6Nt+nQGY6xzppW6qbBrp0Uf2joaX5kfeN
UW3xPOWzYx/y6sl7T3V14/uu+Z9NcRR9a4ytJcNb+DWNf2yx3ES1d9FI5OkwM5gOHljs4KDjGEBP
1vfwF5jm40E8ot8gZO4h0W8dZtwLcEXykpL8hUpFXTeFeOrWMacqWzrHu9Y5KU/BI2VXSafufYRv
oNaxJMZnUU3nBgNmPHW3GTrcDPUR+5FAmBZtGMzRxgNX3NxjLeHXMNXIs5L36+Cxg5EXrlW3bc5U
7t9Slp1oCwp4ZBVODitLDLkfgd3EdtfroFuh2oDDRj6kPK+5SW0PceoaIqBQdXYJNA0fhP64OksC
919V5hh2j8UF6s2u6NH+45do8EIx4/p897E/VUa78SflLaKw4P+d9B+1VnywoQJKvabhWj5497Jw
4li/NqV1alL9skazwEWAIcIEu4pXfRqHzxuwBbd0HXBKzei6sHyMON3ambV7X9zfB5idonWje73y
Rot/qEQu53LyKaDAJdhQk+DiE48+RYAs6l75NyHn2QFcq5SP9AaTeDTbo9VXKbjiMIEtbDNzqIht
C3rhgEYn1X629Lq6H/nXn3X/fb+EmFReN6DgpheeNLGOORbbUgKQZtmtsgFIlLilZWQvoKTU4pEh
N/+O8g/Ame04QnDWYD64VC0NoAI48mmN7Rn2w8BKhZyJBK53O1IghSsrsmYAl3tHzlyl+KqBSHKL
Z/VYL5QsXqsmYvFjy1Ihun6YF4AAHZI+XfQjlUTxF3tZQbWWEwk3SlRENVZXuZLU3ZP3OE5ZdfGp
nyD6GtPtFV1iwvKPioc43ycyHB3gJJgb4Ub2Ol8FnWbWdvooS126r3IfKFxsJo7svhU/GtQaOqyE
L6mRv/HFCb/++XYkFqh+EOCvjrXofBaye0jzdUhc1vkOnx79V9k9HDowy3Pe7TdKkAxUAxKezgfx
EHlbGYf1pza998rrRsyaC9SDyXmim0W1C0cXNZp15alFPMM04XDj0OjqBAX4iFiz5C91BfsaMOYC
2AHdl+zdWhXU7e0ScM5s+ZU5umhX0abQ2V0BCyfp2R9SbIoVQr64oBel9x00xVE/cp8KzVZE/55D
dODOKau2VVDdzFE+R8X0KnItPmTD6vCVG/TPEkiA46KRYEx0z0QIPpSMvPyHUFHPh5UNa0gEMa8E
zBDY0CGxR2fi2LWSZrKvsKFjuTW7EnSEamHWenijFuLe4lEpQqvzLLShj75kBrh04Q8wh9Ky6ozU
5LhlnHtHClSQEyLQA8QfAyah0RNWYRmzAuf24pv/zKpM9gS3hzjMJjQ2gcjttRGmtYlzml+8IgZi
BVkYjMJqqSt9YWLZExVKjZIoaG3CkSwPuDNLVFe0sipUTlkVvYvE/eM/OKBjrVWSpTo1Nj0S3k5+
MOo+57VW2C+eBsCpHkB0PQlaZ0jqlfp9ApuX11LlX8+9xeOJjc+t3zgynpZXTP+3OvIDK4Nmcii5
QKMuPBbmdh9O17auK6camC6MZg+n8k8jmIKruo6+PvUvJt6+54nFNj59eiDz0K8dtlmqMen7755s
ObgdxRm5f8JuNeTlTeaAp9amgN0S1To6OD+8CyQgq/nGgDYGIn6GJvOOeYAhsGr/oQZ7swDkcVVv
RZi0hEOBztlctqDE4YCdLAONQFF+p0SE8+7le73NiKL8e/EFR8DYcI+INCyPg/Q1lFmIk812VgBc
m4JZdgo8vevvdZtIlnt2AoI8RjqGmXWkTPkRYvBBFXdJASawN7H9KeCJgr8OQ+oXQ4/lBm3jHQCR
UmlIs3JeVFkL2ECKYCL7qc5rSvG8UzyW2N/GniP6CgVfUDJl0Lc/DzuYE/3EL2FRdMMyHPRl6vAr
AsfsQFSav1BGfnXwPlRjDke159J2H/3n8wOvqlIzuNeZGC3vPtHSilLvWlTdvcqS86ojNXb+HGRa
JXHO97VnC1hNf48lPYbemzwcugUqHR5SS8Kd3rhVTVSpNgMOyDZ6GGPlG1fmNX/teqIIFPkAGQnX
SXoGg3OeO/MXf/t4JikjyZYrSQHyfQI5EVRDW0SlEKP0Q7Zn9u9rnqPO9bWsFngUnRhK+1JV1Ys4
ydWs7PelP4eriu2Jk3uCWoc2pyF9fGq6XGHYLPsMGA5Xmrhb3vcS6RH8Cu3kDP9k3uTj0OS88OQF
YmoY2XzfwhYOvkrqu7c9mUz5fngPwKz6A1aqVGZjzkf77Zd0KolHbCoSpe2KFh71ugTnyHOwkRQL
aKLl95Vkjj2z7vJcO6+OYhkncSPVZfdc1mBbxVXVtj12byo6aZL1izv7ewmkt/LEJflETqJDxATI
BL8dC55/wU77h41XsehuRoSldrGxHqRqLw9I7V2CJbfL7YwRMv86TXOr9dyg2VIJbiiyekeksCV7
j02y0HUXfwxtihhWjOhkFGWH80V7abeyVsz4tjKk9QYWEy5C2N1SIqEaGwzjkHEanRbqdggxNuLw
AIRLYpsRu44YWCHAgaW+uetf3DSgJFtFWOfNRNIxLGrGLn290CG2hKnnc9fIUVXPc4IcfX+UTNd3
60o2R8l8q/82tAzk3/ZzwiMWY9VGvEjA4p4zG6213jqStIjBa5AG2QRLNg1MxxbrhXXpRX7JDEQ0
eKTg20OVOccJjwDlhh75GKtZD1l+OEMpxyuxIctGGDZP7jPP4NgcvPvG0pjvzZWSRDsfp1lakqSN
8wT78QYFB9jaIyZwTxxRv0Dgq/S9JJIy+DSxgjNufXlHWKDYQ2SXINRnm4TMtDgWqW/YQ5Igl1VY
2gP2shskZ2WMIpWT0yUM57DSG5K+r0nWrK8DrZmy8GiwEqBw7vFZPlNIQilFAbvKJ1BKzpOeqkDM
J+yQZ+wSgxa5KqG8zLfN99z4ASGkQYz1B1bzkUotT/fbcNNnpo5Wi+nq1r/xot223aGPjP3v13XK
dhafXjsZwbwoUSnbNHDacjX8fkgGIEiEvglIktpVt3esu8bgtYMXSFOzMzr0WW5Osr4NSC24XBh6
SZaZg70AdcWXtuhYzpEWj7XTU207wF/B0LIJy/wvfYk7EpooySd1QFZG3/uNw60ZdUpkPpdtxuzU
wbNtbKDqWVE5znZouKhvPOdSKyMypaxrmMbualdpUJ/35uoUrYtatMOaWQFK2o5x7kwEBQdo0FHt
xWFI6JNQP2XScRQ2FAa8R5qSj1sgCVHYUkQzJAmbQHtXlLn1xloozEmkU3sb67H4IUuVlEY6l9eE
NKNw26j7ubVXe03u1yBRCm/Q/Xa00pA1CDGWnWiNXSewBniUaiN4a9CXVk0O01g0wE1WTlpDjK07
aY5NfFInhOQFEGcBTR1oX/ZoDK3fuqpLOwa0PaQ4KUZYGAWkR3DydLPean7urNl1cvIKXE0L20sO
k2NsYifpw8V38ier459Lqvl41ZWKG885oMmAdzDjRjrqKjm5WVZa56vctHqUEcg2+aZEukiB3ct0
V4e4VvMShSVVAoG0ff212YYe5AJiVd7FuRY3tujRpS66gBWmF5p22AQyiEY8GUmnm4AYuq7JvavG
BImiyXoRXD2pqp6Bi9wqRSBru6vE87PQg9GDnUU2jD6wsKV4X5txO4lfVbAGz7jVpA8kGfMiznDB
S+rmBQ+H10CErK4LaP06apYRKp5l7UVkyasQcfO4Fs2ORZKZAbRVHxFpWwhjMXZIzR4K59zbAFn1
5OlKDjuN5wJlPF8t5lCPS3ToEeCiYQg1TpknKVJqGiznAaH2j+d+zoZvHyuHypVf2Z9fZzE4pqad
ZXFVFVW2+tR39PPtEIB4DDxDqk5+yCJrWqZO9YDaQBBRpPPWOZkXqxU7wo9VeooLZZZwdy5Kywzp
ewqum4eVeK73aZO8GvAoEPd7JsERqLM43VCQ7Ir52QUA3TycEMUa1JClUl/jJPOwYFjkZO7wSjjO
aPJqBz2Mr6FJXosiGhwu491QVaMFTuyDsPh3PzoC/OW9cHaQn15UAOyuV1drovvRqyZ7nxW24Fq4
E5O5boIAjm4P/dMpkHyBLKMujrNEoHXeNJ6tGwrVRUqezkW+d6nB9ZhA3lCDybDaWqOgjpU7mFK8
XGmvjXSEUVQkgXc7+uyCwitzxnIguc4np9KMBUib7GqFAZRyCM9ltNuU+mA/mNtBp0HJ8/IEe/uT
Q218aZ/LOtBImQu3msw7SWNM5Yp66+QcFY7klC/F285XOuCR/AarMZQbTJ/qHck23fOqLpyofY8b
oMQcl4T6Ht8NLdYgT2qbCjG3qK03kaaoR0xQYVmUWFm2d9zKIDX8cXDQfkFobCM1LvaNjg7gZtw0
IoPlLtSmb6Ljzenc4FYK4arUezKc/j9NeGEvCnq5RjFW11crE4WwrmPdS71DXMh8eRjDkbaBs0sF
DEgPtT0H6HKFgAzDPEegI/1Q34b8yoSDBEXnlonSjA2wTr5/v2tn1ePjLdLeqYc+h66RzWogfeK4
5olXDPSzLd5zZVEb0no7IwmwyoIcWz42GslLWAzjQLW9kV8kchlznu4NqfAwCNyV4MX866By5VAA
uOK5ECpjEnIWIMXeuDk5LfxKRaahT27bkKx86C3io3ZnMgR/xB60FAdjqeG/ZqGgKawJqAiOq4Xt
kJUTrda0GW3V4pgO/S6onvVIeR3WGX7HMlo0yPpxx2xyi1D0A9plG5ZhSw/GxpZyfpf9oJYW2pyS
ng1VNE5sJSFtvYaezqygFHzvqgOouREut3xI7v2LA4O02xkAy/IXHGkPblszFqHikEYTmFByJvOk
+rOIut8JxjGNnIVjB22GUvCeaqqrMjqgIBWrapc4I4+pd5pZuLauEPzEC6sNVZVqt690UL6d0DwA
+XWJIMST9Z8bfoGMQqGFimJP6FwsvgZYg94jNHAAwUxsXFbsEPnTn7Spv7Q7+qjTCFeab8pvaxNh
v8B0VA7jnKzhZVD4Q8dlSo5CGfnxM8IsFPuO1nBeua5mAPSWyL43upSfJ4xz3zd5/bkLHcyLqT2D
GJ57PDDxEXvBHVzX1a3ff0KnlLtnZPF3TGLVLk9Ld2zAmTeRH+ZxNa5RnOHg2c0zgr+ZxH5bHXQc
y9Jn5mpy84F7U1y72tig+oc4+ZvKKHJzubpmskMmBehozjMtAViOUgzeWVoxRQoQM+qdGLaKxz5e
/6n7JxTHs60UTwoByc6I/Cssnt4S7Tx6Y6J25BSqqYDvx4lHZt2d81v2zATEJo48KGLjo4Qgt0Dk
5NbhQJIueKbT+vpWfdhofUVCwHmVEOcsZ3Ldv4B8KWmkw4FkSfPS52F2LDNj+w5oUdStV4BM5m0Y
EAknV3s7I3hop5P7SSYPw2OmCEw/s+OcX7aQy1Qg/iIwAjRYlaqEGKgky5rMD9+mTlPqUdr2oL/S
IXOs1zB/HdmyLRFcDWS5hiTuvDo5i9rs8ctsL3Vp8JOV/EEOuVkfzdrB4TV9lm5775UIVflZM2Er
EXJU0vIE+36f2hAB1VQHJymYA2aRZl6tPh3I+02dojT1/PUsaJptjS0L0Px2Tv5Y8jGaMz5YTR/e
KorqYL35Q0lAb8f+cSZG7wE+FOoQFJCP1LCW1/hc6aXcnjttkLkqSX4MPno2xFNuSd/BxKq60gkN
G8TGPGV5hshr8a32T8uAc8cPLOfcd0sgZIxOfBq0RSP1OrK0laFVbz6wCVGEJ14OOvhjax+TXP6B
eI2cfVSpULK9GlhjQl9c5XAeaRFzS7EMorUfDM18682k1xut7fR9ToHiNESATI+VsesUeF71iFly
6r4dP1k2xkeTKGphhy9qx/jApcMIXTqKBMgdb94WbeM3X4X3X4+hFRxKn9jEkIw16cTMxwaambrF
LS7aOxWf/aFqtQ1EIHAS6SoPxDQa8Y9nVba+9ApPJS6tbBjUekSQcdwOw6kx5npwuyOVaTSLYZu/
X7+yG7DvY91B0cIqupWS3rzijCIu76dXPSf08ttyyJGrHV3Il5tLqj7/JXSki4tGLWf4Q+fRtI07
0zKTYc6+YS5/AfjBF4pQoU5NvcsEJdtD4B/o4RPl4c3A7NCxkx0TthNTRZxSDJm/OWEOeFpSmJUl
rA/XoWd03EiZwA2FwJGHmRZum5Ap/FGbly2aqF6J8YB7QBEcOBw3M9aIjTV6n5YkHjhTkF4IVufW
CPup3H2hwetc6+XB0hXhwRghIt26F3Be108W1s0Xz5CSSlp4rJt2a7GxurndQlVqkXzXbTn8xbDI
ezUWEWVhO0588ufx4k2DTDHaevriUDWLiQg0fB57k51ANQvkf5KKFhummWl0B1I96rneGmo33Smx
71YMOk1PUnAyL21+SpQ6MkSa+LpvvAmQDg4HLnqnrUklHG3DRwZP12YanY94c1ons+24DGF4I4sR
DgJNU+8ykzyhe8KB6B7ETTCZWUx85M36SDej4yZXZx60CKZOFK9Mgg2hE/0go/YGeANBDY3e+QWn
/VUgj21ctEZqOGWkabmPSzMlRDWkv3sp7P3+1XGTioBmBV79xdmnl4bevl07ou8AiKpIFjhldc9F
QXiTVZGyFo9alw4JKM1iV15OFXC0W0Qa1BP7FB+zxnGbrWNUy4gfewcokjrE+J52wzVNL0uyb9SS
OmB10qPezVZi7WceFPwUERwqJF1ugsaUSN6gEQ/OnNYC02LLPwhoAj60WphRYp/Kwtv5ddfjvWdu
wgihr1GcCl+V1IgRTgyepxOus2HwvyYC+QER4ryxj5zkmxBhKFzT5q7rFFUDPEdf/q8aSlMK8gMS
HwQKASzFx/h+2XLPxpqVrxRXU88WcSvEfas1N4ZgTsLEZlz6kNBQ4a5+CkyOIGWL4A/bAjAeoBe+
p/4pSKQ3r3KTmXQKbV8svBVe3JwZF9dle0EcmaYzfk0G7epQzhEPtieMGsyJO6pc+Mxflk2i7Fj0
lZ2aB43bepGTxkHIm0G5W8pG/+wbKpYO3V/8bodj63TXNqmIMCnqStL+ycaN56BPjbtAW32Nc90O
GaUyE9wysH6fkPFfaWQl+t7KEs7pu9LtjkXgQVmNWTvYQ2esB7KhAvgTxm3lN/SuInL7xhn4VJbK
6fl60i1q3wwcL/s3aHiRsrGHVa6pfTpFINAFIPKMjtmDh6an6qN1n2St4ncemQZhReFnffg8POuP
ar1qrxy7J3ndalmgcWkhQMa5g1tUTRb2WJslrbjr74BIZEv3SdVDOd4qbz3cRkqeqvDCh4VqD5NI
0/a2eF3GBuYyhRKR2Hs+L2Kw7HrMSUpd4jtLMz1ihbu7qxkTZSNXgijzDOebgBZ629YSHw4La7zU
Z0loZC8yHmBpvAbCClrIWNI531WieJIWLEvM/JOZz/aahm35UhdPu4ejkGjEkQy+3zc/oeMnaOGr
aM6cqV34p9DoNsO3vZASVOkUrMXk2FvMtcp9hE/8O5pqC3mEC73elp7s4t86NPaCx39+zhME85h9
BdR7vzGMYaVmkBonK3QWfO9ddcv8UYQKP/5accURRyrqr2tOOxSe1PpwblrEzAInuyAelNWjG+I1
6jNOTfOIe5dlGbF4TElY6uRRHoJzD4jci4gKAHGIeutDLSGNxc6Mdqfu9B+8qq56HPpwCUwa8lxC
e7ln8Fo+C7/SlcuvyyfjxkELvAXMW3sR0HxGGnSs3igMcRqlsuNfbtxf8cGTtJ+kVc5rwipMgvdZ
e4K+P1CcrjTo1DF6U2Azp482gNMpWTp+Ps2kumOhlyEQbLR3pd2QUpyZDcmK/AE92/h/XojJaZcz
gBXFxKcN/XaNin9OuKm+N6UG60YItx3+P/uQ6ayuGomFq2yHWXjGHb74Dom46kk/Kwmyuun14mPC
2dOmZMrJF61bkY4OYStU1m9DQ9pUJyPQrm5UAcigz8odXPcmCeZqznmldQ/+dzepiOvUpe7q1U3H
tkC9BC/lJ+9DLfPlif6sNZRba62qx/ajdHOPlzhYETHpqRD75Q2Z30GCdPBpDxwTz1xZku9/F9Hn
0g8jF2NsqNN+KR/5Olu29XpNvpFaTbac08t0idcvTSQSuDNwqG2Zz+mOOy9ERW3VbU1U6YTETwRD
YIXUhVkmLWDZRABkgPBbqi1ihPhvvkNLdKQqFUdhlEodWo+XKs4EQAS1R2YIilcxrYLOjAnxpV7Y
0empNgRESQdyUTz5pvpDIFTCVrZalCr4mLX5f9ej8DpCl9GQDGMKZ3zogFHe9z/rhXih2CTNyG40
5Dum+yI+SIL9zyV0ITd0rzU5trPaUL0OIVZVD2ATHrDRVRcq0oGo2VNbltycwOdiCZK88+31NsOa
0pVjf/JgmPk6VPLYkxqUTgrS1/iB3VmYe5gqLpNmPAkiKHKS0R7ON+rJSI6B2szk7ped6LyYt6MZ
6LsaQOe2tY0xTQAMNohYJOhEwULUZDyt2RKb9AIMa4HGrERu5QLFiMykfGYrKm1yZh+pZKZXfaoK
devLgmxmD0y4iXORxkq0hIbr37kguucc+bG1AI+6EpFWAYVon0qBPWVq08HxVOciKA5VVSR2PBst
xS5gvb+mnSAy/vZ4BZt297rtuWaRZ7E8Y1y/+Ks9fcsw0y/SSUZ3eCX/OnFoSLBd8g3SOVYCbxq1
7KnO4iY52rLgxckdpkKuQvIC4oVWdjPysV8Lw1zqJci7t4eTGIT7MCM7hBw7TusCGTubJb1Qo66I
BSzBp+J6aE4IN0So6Tht4HLdbgD8am77LKi7e/XjXoR+F9B0BPWkqGEYmSwnVqiHBODGm6eOxNu0
31PPLot7uIkpRlVAgeLX3692lw8PmFCd0qAOR/ifmPGra7+RtwBjIsTO++HTwHxJBd1zexVmdr6u
kguOcvEl/VQta0+aP1FNZPJ7FPTQMf9qoODk82F2CH7tUzc0TsuKNc0YKiKyTPKBoNE+iRDnIdaX
u3Cqpw/ayqDNByNOdW6manLdRX/72XpVxfI+CTh/vuZbu3jC8MZWOFxi1HOTvImHZhAdTBDt0tFS
/9lO+PEMKMBwV9/RvdxwbJBtHk/qUPK6d6TIR7eUYvkIfcClyU99aSnBDfbB5o5pwlWf5qQ7WkGO
6eCzGUA60d+4NSU1pZxsSDIjqmUxVMePZtwtn3o8atavWO492Qliv2rr8bqX/l4sSH5ytex9C3f3
GXkIUe5eQZflluNyS3kG/nO8BKPGyoNDXsXKl3+/yTQ753xO7k4raV8R/HmpofJuNwO7SHdm9I4C
sr1CmummU+1aWzHQ0Vh3zCxvDYXPm/lYl4jQ/6TSjrd9FlHihuO4F/VNjATG+hUhx0LqjhP+xdmP
/qKy8HoO8K1yoncLkgzbC7DDBdNp/CDEYlfkqgcNIRkiETK4sncXqq3XqUYCscWt+xR0i7nJKrYm
76ASOMIRIGbpyuy1u90faEbZYSr2PcsTXAfV13DIcqFsYeneB3YerBLYU4xZKvGRXrd8tp5QyXLq
5YGA5mu4TG2lLBWUZedgsyyYlxrEeb5u2trknTii9mp8vF6VywCEW/XDnJC+rwc3B+81qwV4H0n+
GsixXpc7z8GgNA2K9xPX2M/MdN02uhAWApuC1pibkFp9t0kqo8tj5ThYJ0Bwlz6PQB3+ilUyoZeN
raHWMulY55J34KBZ0na3pzpu5a0YBfZuO2xurh3U9BpXBE4ye4dZeVWcCR4cuharO6LfOaaM7ahM
75JxcMPnvmPQ8QqMxCEwXedGhXfVMtg7GE0wCCzP85wXawqsyv6fBgkr/yna5QkP/96I2OcprThw
tU+C7hXZp6qDL6P8ahmn+R+pYXgv866D5dNAI6rvdrlcK40IUzVwzqYK7darUkJynbIggD0fR/jb
O7A3UxNmnr2aI3m8TVhBQauPduTvlDP2oL28KjT7N9CLJBhN5QgFn/fRF91RfkIA/JFD4VehIb14
sIjugJVDjhOFfMJkJehiGiS2lFv1iXkzE04NtYra8noBVpcLYniudkjbGyQpUj65z3CvFDKk57Cx
mSzluajDXMizqHSwzoT58PAmVlARkobWALWp3S5PzY0mmP7XYsj3WuHIT9nj0kLyL9ZxEPAklKWf
/G6ETfE6MlBM1t0NOfLxT6C3xwh41i0ApGaF+X5/1Vm79xLwXqINjfqapeDBmW1Y7DVsvAjA/HKl
qOBM7Nreur7SnrBYFbDaw9gYNwc+mWDwYLs2Cd/DnwoK9aiy6MOGzqvR+EkDVLtT/wa+BXcBH+zR
09fMMuFuFna58TGFZVuXxWbathIM1lewVzXVzz8O0FlgkAfyD4WnqRce1v4+wz1FA5XyuAgpp1Ga
RU3gVYcO9UAXbzqwByfGM2Cb5D03vsUvB05w5vrae2WRdFs+/D1CCdr6snj8t/OTXGgdKS0OJePd
mkB8/AlkYfzXMwsgsCpcFKAf3YI8EtwTaEQ7XvCGgmGunHx2WrPMLVGSnwB6Cq4ID0V0CaVozUtY
5SZNneY3rOVebeSo7PlwSB2VIldriruF1bs0BRCcEUWzUBHhtOIHFjjAJULMdVfBIOfVmRS0ToTU
iwRGhkDHkbwsOqrpwt53duPAPkMj1CFG1u3lof76bF9DIQuetWsUR+jiZFp+uQYDn607CxVPcTIa
VgPIPsLwIYVW8H0nrRZppBB0sjVQFQQLHD5GHFceFLEHm/wnq4MD4iGjI0LnV8Yyj5wFni4FNhmy
zq6skG+H5R1Yyf9htpCT34t2r7/y7rY5YAr7XJcmhmb0tdV0Npjb3KNzXQDhXr7bOggpJe3YKH9s
qjVWYclwHkvm4OvtFioL0pgKDIIUE29I/trW3i6sq8W194JnWTNDlKVEWZoOI+fZ4SgX7VIREx2z
GmwRvBqQdlwIgrz0CcGlxz6czijxJmvDFEA+AWmSbpCll4nVZFVCdFVtjNxQzTzY9XMipOFs+HCV
uX1HOcfRDygBUDpiKggg65Wmsf+TAuN0TKu5pgILn/dp01MWDP3DHDrLdgpHIU9uveL3LmZPMFCD
bpLRFudYOTPrCCwv2Og1riMXzkGSR2QT4wggfsucTsrcHCMQtCYPTZ/sF10JPvi4oHIKgcP18bqb
HoPS+de8ZK/rWUJo3alyALvFWqZGcAQK9JxGNByVVL/zb3NzKMXMdWoFENxbe4uJ2LzGORXf9/bU
7ps3gM5kiZGTSfcm5YbnzRnrQhVGSyZl04U1bmLX9t9F/BjJI7CxfJxDn/Pww6IW9loYk+2n9RJb
pmP7Wd30iao8sLYKHNv5oxMzuT3PT84Ektob+V925oaDOoF8wRc490wiqc/Qc3QD0rpOPtoOq7Kk
8SR7C9cHVkMYJNx9K/+qFLrM7RZV5qgk9nVDPyyoLdDtKcVG1zIpjwRIK2JN/FF8haTucMEtekYa
x4VR0FytpHVPKUL8AbAOrFszGhS/eyg9LZpfCPOmKN6sa1lWlT1M7AxSTQ4mpM7KjRy9akFN4zjM
spl0sw3XPK5KbyN8T13idzbHu1QhxdvNtJlpnKHcupRy1ggeQcvTTZq76RPPfJHbl9mWGimZsyjK
3Xk6uogxaOvHAAbwwutblIAN1irlRWj2AnuZkvpvpFCYLX1A3/MTcjOh3Ymz0PBA4vNJLzMExAkj
BBWAYmc88o9EiTmRLKSZhfwbQ2bb6UNq0T3/gMSHh6I203waEQtNqXab4ypBfj3jsRD4GYWt0jef
phTY0xMGqBmagTyH7xCtQb0zb6eGijgtXDy5WxLUK779k6gdVl6DfL3LhSRBWJc8/eCm9V2f5iOh
UTB6KLEEYr9G7Bvmq7C4AaZyEF8FFyGBe5KKKqes6uXhBc2Bxi75T3lhHfxqZ/bLd66M7DvSVVRM
YTFjD5f7gbrWDOem76xPhsiXuF7O4q5I8VjNur9fcHUojeuDhCHzxlk4QxWLEuR9robxyEp41cgs
MWjsoVqRgeTZZh+iIV2xH+rk6pGZH3GwBTbq5UShadG5MBmEN3mSN2YtO9o89IcIRh2n8dRPKdgF
EkS+QMVKJU/lChy1FokMkSuh0g8Hvlh03hiKIpuAyFPhJp5Iy2M0eLHa9WLUmJuyEdjjsnc/cOpZ
GdTYMAgZra89yTSutmc/LIMAegEljOO753vrdAQ8+Ryvm0ufK1s8/nkE3Gy4bvg0bE1TsWNemlzY
jGHiKTE/2YTGdYuUScjtN93VdrWvn7gISE4ZV2VwWEbJdXJQ0a2vV0PUoYp2VIUMmf6Wf5Rh8Vbv
+fXcMVBYHxu+5qvDNfnbhZWGK+4VHbYNvGr+7cjAD6EvtaUXLTfknbz+lhLeLDzrmsUvH+tnGOKM
fvMVIxL7PCtbAKeZ6UfOisHL09oaVAjEuDiGefcy9BzkR6atgnQC1dwbQqLGttDAGNyZ/jL4A+0G
ED+7qMudAFsPPKVZbQeWpsh95r8kQwqePQKdELhnS3TZTfQ9mPdDYIHUJBermLRdpHVURMMEQEWo
X/iBXfh3NYLktCV0J3wqkJJOZ8cX/2WYOXfU+ynuGp2scK0rwicfm7oYhu0Fd5+QBfrSOKwDwpMk
TUT9KKzSFdm5LIDqc+7CC44uF7E2Wp5KeuEtMgUl9MUykTbW19/I/fDTmGLp/C3lSvAT/x+9NMme
4Uj2tGwmQICuuwCH/mhz0WWxJ/YrzxfKeLB2z6rSagZWZu50OKIBpcidrVl+py9IcHMgHeJvveI+
bUwzw9T67eTcZ8cCBEcXUedLxfI1KunEpzYN9N8KkTjaFPmhxBv6XbbH47wDThDaJpIMr1xN2+wa
BbFPfi6I1nEdvd8Efhz+bMka3JqIJTlJzLw4yo5JGz53llT5UFJF6QQ5Yg0vIbam3UXQOPYCQ2LJ
Gy2PzHrW4Rirson4vWQNytSCRMqw0vHm5sXGzmrDQmpEH2KLvrLbI/XugZVrFBZ2vgbFsP6z8Yg+
MMYELM4PzwmK+g4dNWoY2DVRZdiZEnSHF6NmVHHkMzKFImZomY9d++seAF3WyiAfiS4lgPve36ZX
4sapunAdF7eVy66RMU8jwM30PAecyRzRh7dq4lxUTc7kWWSIZ7KrQoVncZHhL6YraR1iUBAqBhsy
G9YPtQZJei4aqpvbo2ZHQxEvd8AP1WjNqj51zg/pTx3LBviAxjFBktXZf9u3o9b71/c9YV7uenfc
c9nu9uLqoXgJbpmEiz8s1jbCWF1Wzh378X7fAeagWqtYbmqoDB1boJAusg2nZd8wU54pRPQl9dAP
/O32NbsayrtChyHUJflSoUTAtBR9mtniy/b9p0jGeR6b6RY9WNtRRyw4kPCKKzsG+93ASy82lPwU
H3//oZZo1WAG/cTHqDoUKWv98R54sbZ6oSrYFBAH1OjHHtoaj3MxQwK5jgvX3qPquWA+wXEooV2s
il0FAe1eKV3y3rcJ91KJ1ou01n/C2ZWNeT8FtgdKuEdlPpIh8HqPqjApd1/4RHUN7N2dttM9mnCw
dv84peSRpa/WnGO968RwNbvhLWQVN3FkYRZ1KjF9n5QgIj9+i85iRgQV2DEuw34KZBvfrYSNNGxu
SW2c4ivK8uLC2L3MVzT/Y7Fn4/hI0MqVDrBGblt73nY3EZGsFcn3W5oQSOZkRBwxXGy6itaj7SyT
ok8h6Jz21ku3PDoByjjFJbL2PeJ0sz4EnRd68PlRMOxz7BqH4zRTTE3nV/db7tx7Y+wmMhjVB6px
Fj32mJ0GEXHYphKcyl/DbhugKa59LwB3BetKh4gEWOhDhAl3kaN4NLgRd65z7ePPPLeMNUW5Vjvp
VMd2+SsX9uhoG/5qcqphHAd9/HcdkQ//ep1kvlr5zWoTG7RPRKf1FE5CMUH1a61k+EUecMM0QYgm
7y84nsX0n+tKk7rr786baSSPweuWI+zJ7fIdHzlA/9+RjkDI+jvifnX555nQIM8P9V76RSThZwO2
P+49m7NiPa+vgbpBuuqYmEFuImlccA5geFn4gHeZPTnMYPJ1WR6YW8zn4gGsJsBdyi7L2l817wB4
L+Hab/G1N2LaF1HeMLgLk4Nl3Pls9ukKWEIBVzODso4c35aMVhNY0UhEefZfTlcbANI5Qm3eh0fC
BFLCRiQk6eRDdlozzHkCyaDwJdsGuAaD2bVOq2tY6Fgy1EKet0LxR8YD304RadjnH52w9551xuzM
MizHOK/BennLoanofQDbHNaiAskb+/ahmuSevwfNXyc4ke7ml1TtSphN0GftOOIswHVDAjM2nPgi
SaxnR59AENzNaS9f7/d2/zMGVY+huT7pdkyDuzVWVndkLf2WVHj/z3fA67aVCrXTVw6Pe2R6/A4i
c2u7USduMY9CwCjx0inoiRvSE2N3Ako5yBArJDCLXbE7kB+4bqUFGEyONZe23y8VDIXbM/0NN0el
FPcukhQcFMjkdA2hyh7rLEvx0uLkO2Tn1CkMUGFFoRthu5bssjs4DWsvP9ZGLAXTUjIks4FDc6fc
Z1ELIORSQMUXePtQQIJjMUPwK+131PPRmPmQfHjJnXPoELKNntxQ/DAzeQnjtuXkhzoHD8B/NcCq
DQ7eVCM9K64eXZt/o/KuN2p8qmbpP2FTPY3w16X8v1AA5N/0HFVsNoC62whdhwFVODCsBiECjqZ8
zBZmV3JOnL4zDpA/VVFmnoqFh4sQFQHUPb7Ty8DuTBhcYSa0Jx3kQDr/lMqEDXfeVGvr0yWMOvU5
ElE/qKwgVh+zcaPDiI+6xEdvMLR/XvXmzzJGaKTAN/+CKH+SwdmcqT2pSSb+Macc75NXQ+j83MXZ
yzdaVlMl2CVsp8AUWSiNkqhvqSoyZjsy1l/y0veJ+zuTjfRhgk+a8oGtxMdiQPYSCcoY5Z6CAWbn
VGNPeId72TBZK75ec8UxOkr7WleXfDck/3MMZ3bsVHLMJuo2Yfru6tPw7NOrj//58auRdNlLxdno
XfVQ0iVQG8zCimtg1u9+KIxit69NASw01n8OO3YBwmJ7wgKqj/xG7jsl7sJMjF+pgh8FXk5yqke1
698btNl3Le6L6FGVogxMIR7iHz+duhNem0463++20mUvf8Jp17Oh6Y9czCA8bmqWjJjKTlZscxm1
M08lgX7dcnvSDsLHjEKtgO0U3Ut6hiRJYW0rYeSe4J3tpHSLFLEqKhZ2lUIhoHNl6uTi+6dZ55ua
fKLiAefWwTxrtzyE7G1A4ZF0WvhqXHjA5Y0ALQPufW1VGCwZTtmkmJ5Go0CCvDXiQyGD6vsjLZSN
V7hK5nCPJ3S6nii4JN6khtsAnryAlrr2pNkRYkUcYyG5DR6RCzAaX6+FAdnzrZYK3RF+cS0z66DL
WhpfILQGlsksWmbxU145IeDpNFXixMs2nVUdl8cgiVq4KOmO5rK6t9waOQtAK+CSm3Yk1UvbgGFL
wB6Ecmo68w9fl5OD98nEnVO4XEaUWsOvT6peWQW8EFLMTBLKXs0DN7KQk7Yjs0IaogJX0l0qlKJb
xNuMznggXPy5yAIynqIKwacMQvuLIik7FJS5A3ArTdaHwiqMAZfi8rdt/0/Q737bkZR+ANDPtR7Y
k8vkPx7TmWr7U4uS/zjOhoJbLBUGPHExkv61W8IwULD2Q9+gAZ0ugaupc0q/VTso6oddY/gICBrw
sh0VLBN6fa+9z99BYVrVmvUqK7Heze7fTzqtK8xYaA8NTbxcbz6IDAM8oS/EmOE+VNE9G0YJHQLp
sTuYXzWaB+j43LXAWVUf90bzLAloluhp7H5zODuwPefMtehxVz8V+BCL7fESsOIAaBdOuiiIfOGC
KhDnDvWHMoCJdLbDRhRpfNCglL9z367A2e/o9y/XS6OIAJpSwn+Ghp5rwJjP2cPp+aCbDBS5qvVj
i0PTmLAVhz4+C+/uiJoUho1Q85KFTx5+60OXhyaw4TbB/ViJ3d5K7cA7hPWwbdQEz2XJOK3Ir+LT
d5d0sgphGBBtLRwN1VidQdKcp/weZ3vQ1d+gGTMom/Kd0yBWEQAJJFMhJrdsM4jnThenME5SbphW
Si+EuoWlFJLnPtlcyAIoPOo+GxTWUEpvaj89IgMycU3kyc/zzEls4VAxN58ALRvGUSpcRvUn8oIN
IPKKn09vD01Ab6iqPN5QjZyBIMjqhMU+JSKk3ZUtGkiYDwoAVmlLosbrtQ7tMKMc39TZIAkMzFB/
hbjRNgDGeyL9d0YLtbX5cD1pSWaMA+eqqmT1M0okgqbI71P4towW/aTj7epC1hI0QyWbh2LV+kAO
LWL5Ymzec3gdx2HhDyI5BPa35FioZfy7mav8GJv04gAqnJUtpvNdhskU2qd/PZHqf2nrH2NuEVsy
TFjeyyc82SbXxsi4Cl85pSoQ4RwaKMBDJffOosUg2TTJvfhR929jqHMhhHoDgZo5fGeCg4LrtAAJ
DA0/JOTn2gN7XolVUCO+sw4vKz1C+cM/l7MpEk5D1ixQQVYPvhG5OHMYaCluRqAp4eQF5boXib2F
J8qyMT1PL8VeJU6NarcKQRUNej8qrycbw7l5IZYiMyaLWQ+ODmIsf4eczYWNvaqllDKb2CMd06RT
Z7ZDYCUJ/LoZ6AzYw+cIXVgeQugwQmqsGu0lidZlPmJ4LXsdBc9UUtKPvdMxEPuDXUPp36NmLfrL
5ZH04/VJw2YWLo1qo00KR+oZgEefFXELbcAiocN/h3tuGYzCOltvkuA2pCy4dhUzKtBbYuVAO+et
flFLz93t3g9MDldYt9C0fR7fYuaR3TlBDF0ULe7Io+CQq3tjsz2Z8i56iCXXtP2XJwGJbPARzEe1
3HK0GETO8jiEetfRZ2EZNOJHNyiBeqyEJ0NPOpF9nPYAstP265w0/ZldpRPQcTWH56uXeCwANiLs
buooSkrywiVVw//XlHRFOtZQuJLf7kbDk+Q2TQRZ/H4hlh2t5X3LCF6rSamDj4ZfgUOD9h6YvzVs
74w1OKQbdbM2DwDGYvkS+idDE/PwTmYnuqx2UOsOZqL/Yw7ctUJ7HcnM5kdyPKwNURf6pnVWIfzu
ZZBO3mb4Np5JtQPmLX+0vzKBeTa2AcVHjmk+fw16L29UgTpamJ4RM6vutZrqK9mEyyfeAMXxv59r
IyWpiWpfjgwnNYUb+UPiUpLICfgv+xM0AjbQw5RCy6h20f4S7IyH+0AC7NTqeUVyrjNAE5yeulf/
THk/Hb+7THgK1tsayGI3G/n03A04PhiWPJQ5NhjAXNBdgrU5+9CzbBJ+CKiA9dYplxCtwNZ4mJyg
Hz5E9P8HmSmuFybvHmIXQ2N2ZAImA3iD92AilUn+zsKWtkUoxZEznx1di1qGuDpt1ZE72MOJIe5v
/2UhP+zMcSixto/WB5WH7IOidYTkyYEU6cP3qr0wRV7IChSHMt/3QI1sNpxcJicPoon1loChokHx
WbjUvfdRz4299BVVpNxKGDQJdIyIGHZ/dU+2/qvUKhDOE8R59nsMtgb/R15zJrnywV1mfhANxxZI
/vjQlRQ+jW1HTKq6wAFdLBF+8F1s3MEHb9TaaIFHrIz+1ClPYOAwahunoeHhmatcnEhMa45/uqeK
HuWJA1KjndM6OHG054QfcW3GX6KqmLvvLPCetCad802N3OLsSSnA5odgRJHLtSPulMlYLLHOPQvd
+c8/0+WtgU5S7PqrPAwAoDHCY3tRV/KrrCxN3uV4ke5VTI2QvOvVt0q7fJfqEXpIKuG4BnSUr4MG
QQNWYhziagNN+R+pFEYukkZD8UzsnnviYwMP6C5NFK3Sh59DD929C6Ff8+9j8eRzXMDgLPLLfDo8
4yxCA1qngdPlqDBFVlreLLjN60svwKt0QHJdeQhZrkIV3djfWm4zpYpUyO+z3T5mMNWzpBwZCx7A
b3bzHkda3zbNRhTXikX1s4agIrUREq3DAk6dK93IB5oiZcUwxwtSV8WuZohvWRodXZn2fiV3lhNI
12UEj6+MS0MfHWB7sGOzo4nYEyKpR++pHvxIkw5fCVCxBWDtNWWitNiHxiHYd5Dfwty4YFIgK93n
5KYtH5doTjOvBtQYZnNtRdqBhGITkTPCFEKInVFMIls7jvfslnXtUzBP1wAaH/8xbIhC+vS3pgSC
A6VBY51IjwR5xvriW1bSuwr3FzPd7tXgXoBdB2q/QhNaNcsvM6zYsrcwEocT4IM7dmSGhaNrkHbc
E8FtlOWJq3w2jX4DKvTdH8bo7kOkoQMnmY4fzgeQogFTG0MNIMWs/UeVut+q7BoDsafDuw8Gv7so
0KyE0YihHv/PkUk7UirD0iv8hECUl5oNVu9hQBCp1cGJnpuTX+bIVYVUZ6MUadijpmHcfiJMs04u
zuqo531pogN+O/H7gCy6k3R5LDKdVPKrpbj2EEcH3O1/mk50aGXJK1OplBSA68fzaJIHhW5a7ewq
Qvj0omjykZ3eBS4cWxNpMgFo4Tdnpa1QPCcQRJsE9pLrMhb0/1f3ftqvSpWdE9j882Bg2Zk9oP4c
qtVS+yKLWoRT0jG5Uo7BEum6fmNLZvzcz2uvZStXtGX4WoJNn+ECRcyq8p7UmJsNk95lurqNiuIO
PDf31SQGJj2znX6idWOnVjrYhA/ag8XBCuUnmWEAYNDPVt9/k5NQqAzRoYYa5euVtMW5p5C+OuFG
Y8pmXxnLzo5WRq/Sjf/PFoPliapwFIpq9GLHU/ANuc0dYOm1sjiQ9Vsrd3ju5U9kkLDlRKMbxCoY
CmiTKUWA8kScBVqqfXK2/p2Rn76x3xRPTFt9cPIymBDDbqHCw7RweAo3N1KKLs8pb4Az2AlAzUUC
fSspJtzFcQR+/THL2wmST2ofpq9JWXcitph1ppKhKrtQj50Vb0H4iByu0oRFTbOfOcFIia/DsKzA
eHbanmkF24V3CO8pa9TCJMhwRS5P78aKH8xSSS7MYCEjE6VVH7xmX8fqVpRpqSpl4qx/xjjQ5MyH
xhn19HsZD+PIYa1FNZ1t2qYdczkPHWJjNJoA4yqGRdSR6JolRiu1qp+kpbjoo/0XIRkR/KAGla9T
QKEy/pnroJMk9D3GtEyyihplic1bzUnrfjWA8fOjmtHVe+QCKTMVFt12x6MXY8DIvAQ1jZOesAw2
gnlsc8B2wzWs1mST+/WGa6ZHOlKuL0gM0WyoeWfcacPI25RaSIw1fBJzjYUXWzUE9VGBueXEph8x
XYDCQJjQs2+f7PMvM5f1P9MMFsEUtI6Qc97VJKtxhZhZY1jT5KwcwoV+JoxA84DVeo7vW59v5Oud
u5virhp2NgrHukblO71eKE/L9ZSCsVuoC4dUbsPgksFyH+0ulyQ1T4I42fz6SnS4XxXHPCqoRUfD
jargqFw4itOWiAfX2zrpdN4CO80TIs56WOlASQMJ4rQM927/DUqzxQJmlceaV0gMMJ8O6HfUi4yD
92dgq1XfIVrNiPCjWLV8+V1sKFavPeV0xOTEcANB5TKM08I+LJ3yGEid9mpvgxosnQZKPJld4Nlr
Ndncqd9s8y29upq4bCgWOd5sg3Pnf7bQm/TAf6NfrRgdsejEGtuhZh+jMpyZ9NA12Mc6OztxnTaW
/1ZSjxPa1IkNAoSfDwc3K5Kafjm6GD/1g3ClVTeTZeUW52ifOeoiVokenwJEyY0Ndq7SMsuLe+aS
Z/P216Hep2qozGKVYMywWQQfwpxM5v0yQ0B8IP8I8mxBijK5z26whCQnQWAGypN8xMQYSrwfl0D2
IPel1kAfoScWRzMdDNYbCcq/z9lzDvwyB+yF58vCz2nY8TT9tH2AVu2qhfnk4A/+HX4AkkXOs7QY
PV61SNLG/LTnIs425LanGmIM2YmYw4hqdyeqycIHLkBOcYLCpXCWU1L7ceIEJ1X5xM1CXzhlDEc5
vngElh4asrJvOXaLpalN1kKa/kj56V19xK1tj9HX0FqebA9zakX1ckgqPMZOJTQGhCIWrt1mbLdr
nz8+g3uCxzkhGkQqoWZKhW+4GCaldHhvr+gQWhKnZYpCYgqhYyfQ0YTDPBjtmhjLpuHuEsOWdX6A
hFNWn7dDz0DqJBa0GtHjpWTMElutDL0ssrmaMfFoaVuEAVNgQ05D1u9cO/fGgoQDiv8gNp2bPPez
3U3BuZi68dTbCzI9UaQPoVeFCfqOnamrgTdCfhwnOHhB7Jm/PavtFzk+N+8sfZmi42QqsboTaWV+
jmvvm8rTLs0fr6hhY1rcmFQynV21Mzwt5Ose5qwl9s+SgQ7UnRKmAl7QsqOcQ/2v1/V2yTCAzurm
68ylKHbdnPddd5csUAkLDv8ROMwjqsBat8WN7vR4FvtFfv60BgfsNz50gDDu53A7Jv9qAUqHY1mk
+vkwRbxjTX3+V9qA/C+ZRkSvrxakteaxXXGcqDY9J9CwNeoBGm0WFDMnHNcpKdrk1K4ugeS5xOb9
8b6tkQ9Pd8xhOqGJDhXb17SBHP7H7Nc4ZmIW36urpWi+Qf6P1iEfu2ZtDXc8zBbQXgETDNzvrzTa
bkOfo0w3q0J+hk2SWYrMckhxXFE9AndPpGPgA0OlxmTCKgzPO2RlRotFNFrt/lOOT2jyUFoVPq/O
HtHOWp1dvYo/SddqisfiN22hCoswtq9UXO9eZ4Jo3xSclte9fj5Vkb+NfPzpiN+/pdbTTP91LSTj
rLcOtW0oGV+r4In5mg/KzYqpWwxsVwWUxhYG0Sw3GCd8lWB6+uBiapsMQ2/kL0uvoxBcmES07B5w
Ylgp1INnrOCK59s6IFgN27kkgcX9gL9Ai3AxBhx+M+wOQOOr41BDukfR8YpAZ5bO2SmmbwGZAR9f
Vwipw1ud5lUFgY7o1270k3pK34ktC2mL3i+Au8OCi5D51/NogHoJ1iDFHlCzM1C0/55hVXezRlyi
8lfewuS40GUCoILEsuwyFALiBCMwSaVogIa4e1/cfFvw+WMIE3Gpuuk4vWi7gClK8hYAKQ77s9ZG
HE+N19bM3mFwc+zRDZTmch3fPcKmIyfYgcSdLTkYSeNrl8DdjuBTnk8qFPjj7LVNKvvKwyu1xR3y
Alcxk4ARSAFFXlMciXF/hxewNF74TYyLS0uk25WEa7ox8VOmd9frMPhSLEnYESJibn23pfp8FORI
pKxx9A958cFI118csr02Xbaunsg7yxxslsNJkDq4g9a0RNMoliQWxScuzZEXpsvsAILCZKsmUUDj
0U5firTRg9hTmMvXEiOwr5vLBP+Jqz341lnwzYaPL4O650cp1aEGOLfGeIli3fPela5doSyMc+L2
S6E0z0fXQp5BJBs7I2dc1SDNClw2FrX8LWJwnivghyO3lzSdr4qBIXvtCEk8LT0qataon41ONHzN
VvSDvQCFiKkG3havzg78111fdlNhgLyILScSerLWE6KXyOGXQ+mpwkHDoZyUlHm6+v6dvv7e6J0d
RZ+HJ7N602eizAFBhASB/yopI3demJCAazQIUJiqNlIS/+Tb9Ci25E5UwbFeCwpY4G1aYrrQvYm1
AdWaBTbpxnt7XuVhqjIUItJAemzr9J3IgYh6AMY9Iw9CHV/pIBMo8+vY2Jpl00R3tnijFGrdLoKl
UNAaBWMwumFHwLe282EBB0e47Kz64/dTX6vqIYwOTSSvjdr63VB0CAlTAlN9YaKP+x3qVrt7/3TS
mEti7gQzw+OV6MVRtZxU5VbM+WUWZqyjDKffjKVndHwJmTDsnXynLXO6sDl77NEIuJoSgKrERR+E
clhT1s1RUbKsiP1XZCf2ssyyI2zp2YiXGHTFFxKKvoPUvT9305AmqVu/VoMs8oBmKnyAfkR7YlHT
dvjUTb7Ijc9A5b257JnoHm0o1YWIbOwNcscCKKeAKE0b/Umg8wXHDiJKJgJOZFxA0o95zluriyiW
xnFNufyGURHhHeBa+rwAOTpcblZ+Xy9/rjBvj29B4KRbYlb3aQQXM1U6UeSGzDNpT3yG0Xpt0i9Z
w2Ce15kUh7fIyH7cZAM72uTIhw6SHstYAM3paZh1jYUn40gZyO517IsXsswPHP1XrDn6TCLzszei
1FeY049Mr9G+QtnmcoMml6y+puW33J+8IOteVwVxi5BjsZvgTo9kGV2DzWxLqvSjB/da50k2/Y1K
OAzf0FxyAWbie42U0qrxYE+b3g98fP9IQtJgOtICMPAKAhbbdgSEalXnfUjU06nA8SuLBq1c92BG
LnHQgriIpWkyFQNXUMBqA7fdAot4gjov7NfvqKxH8i9cjE9MOU9tatFyfqAj/sLkWDDS4u2AhusJ
OyJsbKgKnU+ooJ+v/TqAcpEz+1RNQyIQ9f4BiWwEIFkiJW4zSGDhpjY/zIWgy+NFHOApx0SZ//wP
b8/SwmkUYgqD8kGbwIyUHXvfhrzeNtdBspvHVekikdzqXdnced5KfPFD/6oi8i2jwqLoejPcyzpb
FLkcOz9olDXege0JzMEfTGpgzQEsme+HQPsDBEKSoeq+LIvlJXQf2tyz5LUB26EmbmsE/qpY4alJ
TioRGR/hRfx2QzkrqLjCDfdmCtuKhhmN86QBIM/NhU4nyQ5NiFQd7yRCZ52+IfKuQkx5T1uVf0ye
Vr4NRQ34YcJFdGSPvzfjNfc/FwDoXegarNHSEwhjsg+EC6nO2XTN8zBIm4/3ECVPF8O7eGXBUns3
/S+2RS3Mdzfn8tCfgFtlsR0HhSGQrm/zNFGgeCXsjVq/Yhq4+A13jDYfFxxNBBv5awpwRLJiCEyL
TrLVAB7T6kXh8uiSUjmDGqpx4BIs8LsW74N6TECqEcHbqI0x5HTXA0z+4jWlkVjlfi6W1aED5JXL
nP6X8kM8TpRHYWZiRu5zzfLDpvRNufxqD6jlM6kIx1OOqi4weuRwSWsCQybu1cpCXE6ObGSI408j
+DZgoMMPQ6g5qNGHOGUigiYc8uV4u00lrMJLBnlPoFCZw3RcnlRcoMx/NthSzZhBUdmn02E1xGA5
YM0n6iHvDeYBbm/quMh37WENptdMdGhtZcWsZ/bI5Bqi25lJ2w1nvBXQDv9kB1K9VSKYEbs+ptKv
96r7qvpHtTln17XhToUPRwzJIHRkyVUyR3ZlYou6+p5GerI3lMICPOUD/BKLhQcyv+HSoRRpv91v
GJpahqshQemEYqLqYXKaPprsz3RA/8ecnKTb/erqCgNS9ls2YnYF36btpn3dVX3Q6k2VuTK8Kjlu
ApRZrG3GLwe56BgQriTNfnFAOpSp7Gc8V5dfG1Eglr1cqjjJbD1Ah8DjYfUjfyOwggLoyqwSXqzj
F8TZvjUJ/q1wvfBD9N0762/m0Zve1kpqGOAoNWDKdiA37FXG+WCalfx6vyKBcgZngwUWli2bh8Xd
MZesoQZcBMyze1B1tl00Bsay1JJyDCHVfKgiCd95ENkgnxGpAWbDR6Bjpei3OZrBlgIygYyJKsdp
cd5Dn7w5jnTCLLscaWN6lj8XFueKNX1TlWToTx3UFZs8gPO9S6xsLnG7SKXLJzlHk+JdmT0S8hRP
3VWlJRS3Bhts2WFRbQuoes80FTam2serS1lQBdf7oClZu+/SHDIh7Nwhe/uZEM72Oc2BthjDoF5G
SAAtJLuG7sbwzSutjgWTYxEQ+EY32lrzIjSacLHmTFn2oyFE9W85knpUIWla3TlVCPdGgk6j2/wO
KBJPo/gK9sYKR3ZopadRxYfAbXL03DFfM9lsHBKLmdAy8/VqKJZ1s6lTZIPh6gfFAUYF6mZOHVYa
rlaTivf+3WjSAS7SClUNEA3OyMe7MUH8ujGZt3XF8M3t0gP5X7pw7nbqfzpwKprbjGC1wxr+I9Q4
8PLfjcetUCekW9cNAdHcpFZaCIbtf2imp3RWlDSE9w7qSnVPP/ZXwdFwzYL4sdg16mtW64VOT6y4
OATz5x1Uxm4FMXvmhUglQhTxLXQhf5hdq0V+dVzog+NQxPIMt5XVliTHN53dkgqCE/1/RX0+pNgk
GLpJ4M22AAW/Sf8hMdxrMW/W0jCcecJkGBA/t4msQhEN1ea3BM72bFuEkeGDgdSpUsvkpjHky7ys
WC2TgPTvyVknrf50OPkYF5OQuJckh52SFreoUk4qYnsjxFHrXcR9p65sljyYpK2cxTVZSEv+IT0K
5XVRgGjRoKQvBXstUzajDrdWfANPHa3EWKkWZJxCkfNfEH6zx/gtbosJIYjTJnJHybmlaWw6M5wN
4dfZggejzp3Uq53OpZwTtQXXAdqVwUsFnX3AuCBlLZzRVqArNt1nPFwYfCP3/s5Qggp5FTrHzvVK
bCC0qC9wak6ZQ5QSEyuK2/krCtBlt+SSg0sV9b2+xiQjMWQ6wyCnV30163YJFfry1WQo2QCn68bl
Ms6rzU7wvS9MUjv+Eg0J/bqTYGFeb+KPJSnloyUefSH7oJxId6bOncxNDLn5/HWu1nDGSwHjZzaH
RS0p02flfJjw5NCcTg0Ybzx+ixZQ6EDGeLfvzCuK5FVXox8vuuQoBt7TjgiGUGNoriD/ElLBbXMd
sZ+YlxnOR6AARcOAj6fzUHAyy1bokj02AFBt1ZY6z2UUnC6s7QMpKIChLPO/s0TniQ1EYfgRUc34
4bWCc0sFoD00RAV5meDC4ZivYBCa1Q1gxgIpcmpaoTYVuG2FoQ4lvlDozZX4ltPrVuMaVOKW/Sc6
Tribo4GAmStNzLQz5N/tSAm8hLNl6qBEk99EAcEWv5NfNKdWUtv3hJYl5kbko0Yqk0zX5yCW9kcn
kO6SKsFJstFY6PsbAFMxtYxISHEZ9Nhf5OkXK//IEHObVHeJ9FlyXEPM7svVHpfRHqi9QcgHQ7ca
Z9VUEtTXaA9R7sjYHPxfWZCT3POlZyJDvm6IAOfOtRB/G1rMaQndERoGSJkZTT5ck85iDWNzWyrF
p5QgaprTh/e/9s200/e1D3G7ZPswBa0wClUewbB24VV6GK39uGMTXa+xr8PQyggPOStbmFhJu6GN
ntm8Ey0D5R/KiL42nNBF3uvg041Dp+S1SHzNUfS9wedMdcKkdbco9oAcnq5MrXZ8vR70cPU2Hgy6
oz9hFa4VYwOcQSTaECJHaAaJmOHjUwzZA3TVwpSQk9gx+tSu3x6WOCfG5EMGvkyUfIqnocUsFP2L
3mCTPTAeTeYKrV2mjKAOywIa8Lsi0MKmiXdmWpVP2ZLgnaWku4CLdxpNkvXsjPYqMmAap+NBBl+V
uxtvUstn9ZLwNvIEySx81iTQUkK/dLn8G2yWSxBmNAPEb4p6vLoMndQPbWJsnLcrTQ3kFhMJROod
XGGJG4rUJ55EJncpEgGdX+hgESErj1b3iht/Qe9QwPDbl/lKiAet3XOr8F2b3hxOxnjFqNNZcP/2
yfOEHEWPa8hP51v+HN8ufbE4ICbPTMQi+UlZBpXVlw1f8ROh1f/CXJzFc124V3WqQIVprtry454T
p5ndOktuPlFb4O88+EKv1oDhb3vEYFway8296digpdf1ri0xaQCIRK0PRIQkSHpu0LoeRooQe+fh
DvACY1zLOSuOyu+Q30igDdv5IIQDtgZDfnUqZNmmPt+8HBpP0pkBSxtr/qNOUl6c+/FIbXB32VGb
skfKbUAO9r2/XkjzvGlranaftv0mnqksYYbhD1GWoeT41ZIwe7PAZaWmaKQ9+BmV8SxQZ4pITQ/F
LUP1NsTSC+1/cdKKtHeCtND6NfHLnmbmv6svtOuA1GbzO8HPVXIcunjHi9qSlCg0froU9kkJoOoI
ZA+fpp6WGKBP7ahGjB4xxVz+im6+Z17zKivhRhjGkRxLbblB90z30Csfdu/Wd+F2bVVfE5K0ulBF
g8CrsvkkmOXwbG6MiaPFsHd2l2c/LKrwBuyPhbb5jVes1YvVITS8N5nwqN3lC+Oz6TxBoK2w6XC5
Ad4Nk4wQCwBSybRZtLDIxOUlKpvDU84rZxAnbfXzMfepEtx9KBiVa/Qrh2dZmHiB279lufH1aJrf
fI2XMXLpNoJrWSKZulAde2OG+BRovmHEOwnJop0TqCwdAbyDCeHSQhrotL0/v/OZZRZ0ba1NUwfe
8HX3Nu/AQfdp9IKMngoJum7NVQ5cwQaS9Q6pODVJsga7bfPzzlUXemWITjxk9Ed5yG1g/YpboZBB
cY5l+qURQUE7v8tD7yIfNDTW9zwrOZW2YSznjFY1mJ+FrWTCo7xOAbMjxrn9RZ1l/tKBXl1GZUA3
UKlg9VWsVPusVnc+rykxxDF5PWnn35cXmHGSroAhEP4Nxz8Aqc6AM6q+B1V/Hz+YmQn2j7JCMfZX
1PTkZ67+jJaQ9nVt0q9IF4BtsqseJXtAvBUYzWYcsLwu5odOLM9siRicw+ayC8ZMiRRoYJFgDq8s
BvVUoKssp2HFd+HwW6+RC1f3EVqB2F2x4LbcVRnzVLC+5vjr7+QUKFYiqRMhzSNag2nN029Ev3RR
a2d5w+/Qft3f8BK9HApXSpAaGd212szqCtK3mTh2J16RmQjGoTHwIvw7sBKl09d18Bq0Pb1SSfSm
kXeECsEFd4/I3JO6Rxp35Vsa7BHjoeBfDm8eBPDxRuzLbyldCXD6t+Zxh6zAyD7XeELkhTJ2BOKX
kO1yUoWGu1f/q5tgOMkpuJoTRrFsdA0XUnLxg+8NSbuewjNhwADCh0J4vroKJXh+Ri4P8F+hvtkb
QxqrUNlp6YBkRwXmRAsusuHP5297rGrQfaYb5lFHnshRl5cv4+6M3SNIHSaICn2choIFaNxPqlaV
h4rkI56fmsLbXGqSexRE2jQbX2HymZkFA0fZXDE3k+bWW3/086L3xdrqXs9aJlazymVnugs87TaE
3gUZceDt3UMLmSt7AFgx/0hiNofuqCY0QwyS8pym7OKmXfFyolowwx2QmlG27/dndKNJE6s9GI40
vGv8zY42QYjNt+WBV0KejvxlUdfsHzUpVM4BY0HJwOfQhHtoVEnzJtRF4tZgBnL7mN555hZf6x1d
eEbk0aZQ2g3wkRGo4QGsmFw7r5qB/JwrY7YuowGu8xIlxhUeThPx7C+ymGjqNiyJ+laKoBZKkngO
HJvkEarNuZpYZlvLy7e6+qn9ybHJMe8U7aCOTc/5fKc/G0cj/VpXMdHgvBzAIFMTOd34AEax1byV
vO4rfcDBFLzso4kKC73u2yZX3RYSc3mFdFMtZCSEefoPL9LUqCItwIwidt0ac0TEEuM2ZKm+Gj3V
2Ubk0/SKe/VGyMHYEgDraQ32L3koScp7/U/v86j3mufcG7NXCH05Uhg91Nu3TGU7J53243OifZEo
6NuHM/p6a4/QlbDtAIRjsP6asmBmawHREi3TynnJoIDJWuj6MGCQh9xpxJhN0ynrzROmOqAfqDUC
QdkA0kpaQshnu7eHteHmn6T4bdtHOdwM+Tpb9w3RNbt7a/5n+CsDTa0SEwuMz+RAR7MBviwNn2rs
OEnqtZibIFgeIAbrDrlii4tydE+ZKSsbs9Vp4pHU3WSUFZI1WyL2yne/8+6MCgNxMvzDEc2CrztV
k2kv+BJ5mT5E2iqptLnrWIW5QyIsUHsmnORvo23WFlIwV1vHy8IJ3JfhawSFDlC6iA8nF/u7WRrE
hkjc8UF95sOBQcqrOZpjvUsSelDnYTLTbBOSwx/9cB2fC7SO2N2swSyAAqoDTEXjqhNrEhLInYoq
sW1LZEJMkQ4EwUEth43TZV+RM+MBLxucFLtpdLFuXcsL2bf6mjVp6GVCWEoP/4V3BHFM0U+tiaBT
hic5+ilcm7leJwnUdUdId1ycuIPc2u0O8PFzJ+3Tg3a0a05ZcoS6u0+N+2EvMlpJR2w+Bs7MwSTf
D1h3kLJXP2FV7LEkcCcO5bSqo30EoYk/VYbOV561QdPD1od8R35/IGAVqR1DfEUrAvAYViEhIT1I
xyQdgy4XA6mBugfWM+B040sYHnuxEqYOyW3rh+Ql2GdfaBa0uA8FY+R55HO0k+rL0ulmyqtgFNH1
shcl+uiQZoCnbHStYZgzl7q16V36SoHStiagDNWyWV+h0f/+TdB87uRKk9lmIIRAYVu3nOQ+1V/0
AYnFGFjcpXKFv54pqQAD7nNNjkLw1/JOQlUJyLivf5ofa2PutU70UXOy6F8B/XNJd+5cjkTqSvsb
sU/KZri7szZK8QMlTGlGFqVFm0nxnWHg5ApdpHHMPYBy4y5JzfnK6a/thi/yGe0ZyYdTLkKBB4SW
uZDGPqDGhy4G6hu4AMTtq8lxzY1loNu5OMbnTOfJ5wYKOtGz/mRSFlzhD3m2scR3fIC/4LtI1sA1
KjRokyspLLvubSdLqFdqNhosQ7vJaTeJ+TSKDyGpsWXz9rJGdvbxVbLEzzxY+tH7J7j9jYJ1KXSV
ENUwWFbsTxJfNmxoDjUotM0PpdxrufWaGeqTx0B1aepRnkRmNbCjvKisRhYAkMAc9eMPY36JW/nn
oSaktoGlOIjjzHJWBlXe3wiBBmvw5ERsobc/q9MCxnh3c6sGO3K9R7/6fHPWepkvBLZFps4QZBBV
XIFIQAjAyp10APxt7i243e7QSLyuiVFqeV1aJ1FU0ZWqZczT1l0LtsCEXJ1O2VoaCFNZM2Vc1DcV
dV3jr/NnbrL0CQHKBXjosH+SJbxPtGZRRs8aZQ4WvkTyvfyQZezsMu+1q32z47Cz0FfKSu6XJAIK
9xAIAdbVfgyHfRr5Y0k6YaJlwkTXE7LYffqMPwrcT3EUdJu3PTk+ij+td//fflXxmmsr6x3MK/+S
Jumy6RCfhsQt72sUcPngIlQjwWGxI+yDZDlSitlDLsjSaQHfmfISCrxdIQHlrBRaMpas4/Lrb7Sx
6a2xiyUSgY+8NxReV4OkLFFaqOsYVmj2aekp5oZlNCVB8H7bgt09rIpi7ltRnS0No9VgoqA6fHZY
15H46Pmc3ZEzILfohQwv3B3x3jSSXCnvGbCwXor05JSaJNtfY8JZD9C8c4T8FY6d4OdETEsru2qR
v2RC/Zd3pDfBF6H2mWnz/ywmdhs75qEy81SxOPrkzyO3uAXTZD5kepDHqbpHKiaxZGO2mrgOwWAg
DpbOIEryAyjqrPX3wP1V+aUjCu1lMEyApsp1PxnrxbgZrwdoVnjhABdaNWbepHxdRO27xBcYpHXo
9bIpFBfao39qzZtCTJSJpAXDdRhFXsJ1eAMOVspuQfEecoz+gMEYvjluPYEI2FMkkNJDW/Nd9vcg
laguYqwznLtJeXwwwP3Tg0bW8EnxPBinZu6Cn4hLFfNWliX1e5P9zZcihgQa8C/kvSmne9iZpEQV
LwBfaE0n1jA41oZpXnEDR/aYuoru/XdOkyNdLPKqIgddMLOwd2xt6ZtkJuu53cx+skDw+wdHckDC
pefVB4GckF+uD6nhLYTLGJgJuqM8X3mXkqBUqr2j60Zlpzz/8l95+IB74h6g1nV5U10zlM7t3F7a
MjaOfMiVaoTzXzpL0812Ko9augNStiz0SpLMpuea92o1HfNNtR6ZLvSWeQN/a6aWG1HH1C1BQcwW
svWa9jiTZfdsB6bbfXXQsQL84dpt9c7dUJEkMFEys20CRxfFzNZOcyR4j6MYLUSN9NDayMpvWgVf
gkMZ4IV3Zk/HzmMtySO6nAUuGdPkwLgoxk5d59eM7mFPA2E9H8JgTdNNcnCrk3xgKmEMrqpiLo6d
E2cbwp7YE44UZ9VFdeYmrIKDsvdUM+8tbb/aqVF434Iy8+HJz24p7/FvCcqfy1A0ORU1Vz4fE5Yw
LgY4xGKNBlNon+E4gPkj1Q7Dq4XDuA46A5WNDTGAp4yiBwIwN4Sl39MonIgLJ1GMGzpvBWzbV284
6CSU3XKHsV5Sau17/ynYSNhVc6XO7cJEMrK1QpiGz0wd90avJ+HxXUxj+Wf/iNKPrG79/0pf7p8k
lSJxCrF9juAqEcRhvBml51+YAj8GzoNInMCiAHRjygs1SkbYqrJOGSka3ZkAXOO6q1umnM8ghu1M
oxyewqeDK7NfZiTG5aydpYbr4wamSziKxGCGtLQU3AAtNlRZDLBY9Eq6QcBXqBGTv2xzY0k4yypn
lYMi9xlbGZfmnHBufdF5AhiKOhVMa1ds12gJWdrDDR1LFXlOt8we9WY3TYDtL2QC+Po57MSVnSYb
mClEnyv6w5Qawp/TnFVSRQD0zA5PbtOfAwSFQiBcYazkXChOo9eTZjIlp4Pen9hGUDeghBlpo/t3
2lrby2I7Qj7foRZQngt826owiDS/w2aQlCOog/H0RO9PglOlnGL5ld9uv5Bi01+PRqQXHl9GvJu7
Bcrv/KtWqcmJLA3tapbva6u+eCr8caoZz+1A8PgQUak5z2R6ukkpg4bqmmsPwstGg/Rw7QLa5bqZ
Q/Iu0JcG0dDfhZ/jsLEihhl47yKOrAvHODWKJ/jZ8ePZSdimEoUIx9J8V+pcq1bN9qMCzty/XVVj
WWmWWdQdT75I4SVkLGhPeR5lAjak3SLO5kYWi3tU6hqDZao0edC46ryJTQixwvcwpw38nOlPKaSP
C3/WveqciDKhdvQxUM8ZH7hzfi7Y/PvHCCCpgcnKsyU+1+GJjCfZbGW5HpBp3BxmEbh9FWSccEX6
5gd61+YxUUucgbaO7NIq+R7rYY4r4CpuQKdNckv6bO+DIMB4AkdfFKibYtPv1j5wSXLhGKDofAJf
oq5YCpkXDhTw364RJhqEs2DqehWTxoUHEKkgtzSaT0SCMopGMig8ty8msb+CkIun29zgOUZ9MddZ
JswLkyU6psNwCerjKVZRQnkhad2SlbkvFxNQvv7i6Kw4DTs9KtGjmoVu5wv0O8TZm1u8X0mTbF1d
pRA4bFK0QTuBWFZXM3lQATZInQQUl8JlQAzqf/YXqs0P7bMil4CcS89C3wm9aASp9bJ26Wq7OaF3
M5C6SBOxgJNhyZUx5Z5I+XBoFH44EKZxtWV6NSDRZ72SCNkgf2mnlS2ISsLDheoxF7hZSf/Ty7wY
8DZp46x3q0+vMxJ0uHkihf2mCK3apvVnZPh55ldYsqWABR+5SHzuWmh3FqV5KYWHpcnWC9EtMCpK
jBovuIFGY7b7kkNI6BYVKuv7Gq06AM1j7C5QcTvqdY2TVeso1a6SgXhXyVyqRQMMaehRWYLbmSNh
0H4My1dwauB9XsapucjB5au2FJsmAqNgqW3Vdg6o9uvillNuZkMMm3dYDVVG1dcOkUQqN6iWtNdK
1lEVhpoq+NoMf0IgQdNFqNQMmNTOqztBQqkRhHjUHUGhYYRHMR/uAOkhUPXa6CU8Sg57/G71Oxrj
tNsaN+nylB0HDu7RfNUeVJjn1uLAJptwc8C4ILqENIwSDtx2d0NhS/ruHYyIIRpFI6PDMfoUJLA4
ed3bh4Yx+h0C5MIwe/dR8VOz/LJQas6pXhpRqgOYKnOCyH/MLPifl/2cjX2WFI5jtom8WC28ypdZ
8dNE0a6fihqJomuyptV91JlXjC5I8VZDyD7oTKA2YgsO/VqoabmGS6EidXfU4aaFDvXUnCo3JGNH
gECRXP8GwfcGoG1eBvxwhWQtO0Qk1fA1RULyLmfAQO4Zu2aZIxsrO9LbJA013un4OdTnnmWFNSdw
BgZCuQX8qdEjFBpncbUr2G6+HxpxfWD49yjSBwdODyQ+HD86v15lvmXNX3cy2fPpINt5ZppG/0ij
wBzgTqst7HrfyyqybsY+a+Alq95xZC0k2zF5XISFkb3UN5aTg9NEQeAxenBl6JOFS7HAjovtB4hc
G6y4QZRoPEqcCmSMRihgiyD0XUA4sRvrUBC6F/wHeT5aAWIQDRsakSZV221mqJCFZrTXS50M2KXJ
Z08n4U+hZikPMeHQD3wwaY6NdH/KTqlwJSgI0lLDUPj4yygvzFKSoAiEfBsO/CjKho0/zQwBrH5h
wgxKabacETULFg99X7+8TmY9VpheY9BCmugfII09qAppIGSweOyH/rz5HhIpa0xHfEdv8TFvwCr6
b9MqwQikLaSqqlYnykccenxG9Yc61E+TpEAmuuSYEO74g4gYW+bDC0EM5NbSqec2GG/Avi07mhyy
ywxeSr5eTo/6wmSnfs0JXaN82DAvNYC2au7bHcc935L9CLLoHMmT6nbee2+45xQ+UB/HNfSD3R2F
sd/buCA/R+jkoGTjcJNfxC/MA2eoSwaIPfbieujur9SJjjXlbuQsriQFd6RqUtGaiHJ84oLeiajW
lEho2QuEu7rZpFHTzWkUVjCqShhreN6KcizWZLXVYN81fN8a/0aIU06empIpc3T1TqsRYHe2gQ24
pn69U/sSwDmEbRbUHf2dPvNqqCUN8ACSUY3PYcM7/YVwpwggLxix30eF23khLYFtzIMVKMBsbfUq
6QPWgYTfZb3ijaNV22ggLKvMfysaMKkj3LTesYLjORVBXKwa/Z3B/Y/WREI0iHwE78lCXTC3zoQ9
sxmeVdz0W00EaU1oxhEEOOfPGEe4eOD6y1noZAevwHJgMnaczrmRH2ovnFm3ZaJ3AW4vN094lWUl
Oa6SuBdyZRTx+tcro8GypCB0ii6yS60i8gjKb3FQ62spQ2RxDsBuYtMcA6dS2tVGtGreR9UcsFBQ
dRUjJcQbdD35Wr5wwVVhe6WFjpRQpxjts6iKp7JUsH1JB0C8Okt29lmudPxrmckw2vm7l0PEjtOG
Tsbss24n3kVTwVgFdL81ZyiqYbAHtOEfk1y9yDWUUwCWu9vLz6hyU2D7aL4f41qPU7zL4Er33Z/K
8CjSKQGdAXvbRY0vGqhH2eH3Zn7mqnu3zVBX3enrI3f2kouRBEaOFSzUwo1KurobQP4cslYITbbE
3DhsaxPjHpPuKPIZZ1g0IFTTHgMPu++ZDr+CZmS41xBbdareWF6F0jzLagLK2O1F9A9/brO9DLkl
yMxWzpnu7Pl5R/oS1EyHaDJscNSLUB/e2vKZcGGwab43rcIYhgFOgmjHAdj9CTCYhQWNpUW+fImM
Lwkz4uuYQaha0RZopyIjbwg/0D/4wuj67lIvNcRliq5aLDL3nzkhz1I0PeU18Ox53SDnE4VC1A+L
0g1QkwOffASqB06TTQHSJlPKYw==
`pragma protect end_protected
