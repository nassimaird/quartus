`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TEsSPWYTNUUSrjJjVtRBp2TCED+li7v5aSrS8kNxD8JBF87ckX35gNDjZ4TIF9H5
Uc+3+bc7zWQ0gFKwd4e2LqNRA8HQizOq3heRYYyItajPKDTvmsLl3qz3VxqDH9OE
TzpHRp8XP1UGoiW38Qmle9ytOLslMn0me0hJPPuMQyE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7200)
KbNuAdv/zE/nAPOAP6afj0alvhcMO6ykQ0aMi4qTiioxhg3jl/itd7BGfHXTIH6S
0e6B/DLr5YASAGkda1DWs60DthCeDjgVg08sP626fybzwN7zd+Zcl6kJDPN8lU/r
taZ67mta4nA5ozd758zwCiF4Ms+rKq2qj1JP2wWDQzPAwM5v3o6AYQh9mcnfA+lS
CqJmeT9jKT6lTaDuaN18LFatPPxx/1YrVj76qYvXF8Yh16CHkKE6dXf094Ua/1Iq
fNrYJCEug8ZThCDdRJLLCbOK/Ob7aIFDm0Dx8myrM2yisXW3SdUYksgiby94hjXG
byUJ2fIjdTc1Ep4ZFJ+0NBEJyF8Rgt9LOdYKvQj4AmCzFZqNjOEhhpYZhKwJUCKv
B72st5/fTtCuu45cZ6TbXsG0uo6Y4WP8gYC/aUmABieUPCgpZTMP8VCTZdDxdHU5
qRCxCBw0ARxf4++oGQVqgjNQd4XwE6+fmexTmuEVl0pftXdV0SWcit8oVcnCPkGn
fYig22eoJoVsrLv7Ec/Y2C1Uifqsi1IXEAJ99Lugz1IuXel7DFe8Tm3IC8X6tdRS
f2aITOpNXqa+ijCV/hXnpKqdZ+CSm3VOB8c1k7IVC/6tqIO7ssmeq6o0+foSAGCx
Pewzaqtf6tlNRJnvgr8RQzX4XhDzyPj9/JYAYy4q5iTPnE/Jr9DBVHL5eHPWHVL5
IxlPCUJb+XV5clMXjMeM5QsOZyAViQlpTIhz0xnvNmtbPakIlBxSfCc/0Nx3rZHs
YN2ST+KaMUKMV3xjw5Bcwx4opQhcCRsEaLld6NlqkZXwH30z14zMRLHKsMiqkwrz
1POJVbx2Fphu+oBFSOKnbSn6MX/MrT6vptOXg0qQSbbf7xauJUOS0leVcYOqFNdr
F5d0yawH4H+ylxa4FrKOqgx/eareUNTSdxb5suYQK4/0rShOitkLphdE8YQow31u
NDcAOtx45tg0YCXndwHMYUab+onh4rNTWFPrCisRnB6wR8goupYRi9544lW82Owt
C4PQmnnQTUqqoozjAuSHahGpgintyVJktMLMozPcJB6UMm+b7HmNomer7hr43ZHJ
qHbeFV8qtRDo+oop/aa+3Yt/t1gxZti6wJKf1wuTYaZA6hOcKJ7CBebmVnf1g14e
XbD4tNX2nbxsB91m5SWsn8sXqtFeIKNjM9vVxp8SR+drxeeb3I2xKyfFb9RqjmNy
1JoRPcQcXiZaHtJB212LgbUzUKhspUPfwuNLZLj9PAJlyMuD2OYR+lxuwUeyA6X+
X0Nrs//9Ld7zG/LfYGof2O0+Kg0/2A7nLhs94pIzp/t5szQIXOKYZkouUk0jnUcG
lIXORa8DDWUmnQbi1Fch0yDLX6AGmH1we9tNLaCTtKyxXX4FVtXHL9r/mfPMTTDQ
WVkFjpKO3cgL3qLu7Y5oOKHuhFFpBvDJ8eA25y4rdQ6VkdR1bQaa18QKLJv+0EWw
NsihgPN9Ygt9OCF/jiOxI97mHi+5lz8nBhJVpglDpS8IIh3aUNui5bWidCZ78PVk
v2a/uONeHHMd5/AgUre3oQfCpxfhPgIgxHmkWtRl7s9cAEZrTYJdfNP1l3HFsEqa
PTGnbVvV7V3a4bSjwreuOWYdY6vH3pLbnzBgqivCwSa78eSVBgYpcqG9qAWlJ86y
PQBaxgB8tCkSir9iVmcA8qA4ZvcxRnRZ1D+jPByxJ+Fto4HdgMIH2V2eHMckssMA
goSZpxkYEsG5j3KtS/T8qlY9gb5+EtyROX6TalEDxxIuXU+6UEruNJ/lPhZf+ci1
tn/3SWAOWFftoT0RgVC3A5O41QCgZFvjLbi0oy2J/K3plJ9DZWPLB0KUnd6L7rZM
xEoGwkMNZ7HNlZ7LTF+Q6TbKC1hSJWR653I/wfGlAUDrAqd/REElALzOfIjTFiVs
E/g7P9p6T6EBN2mzkZJgOIgMZohFaua+7JtWlq9c+m8nJWeJcgK7u36TzioQLM5t
hK8C9ZaAJB5ZKkVqiVcNTrFhJN/JKB2Vr1EsR9bHe8gk6HXLHPsurachceLpA+v/
6+SxutM4iy93IsACLvMpl4cTjGhMVF+ZoYMwhISvI2WsFBnUDr0cfSpXtetiahcb
zhCjFM4dKZYw+ETTHk7RxtLW9E5MqOhVbTwUGHUpew6bB1oVIWi6xcnyu6PkwV8F
79gutFZBe7Jfcg4v4zmoe+s86Qp+lhhJA75SgRsmGYJ5yhR53VhnbT1/TV2VRsRb
PocP5+CIzzq8lwbUsYtNmQMzxclgaDEfEfDnI7rdt3/iqQ5XisTMgiKyxZijrz8S
tOY53CGE9allJKtVC2yn/sPseQmUphotXhPbXwBNDWwyL5A3Mza3mYeakqvOY2jh
LdEWiGbQsP0Zxid8UFo4j0l2wnh1WDWNlnM7kwnlWa2q5pBRayt3SMVZ+4UK6ZHl
gYDIU2qClEwXuCKti9s7pDgsPghaWmlkcblmCY/wvZCagtXnRl3MmEQGjJNJBCFU
JdnG8/5F67rdTk6JjzvXTgz2nCJFw/leyy09z0aF7v/+WYTZlozMSYu579xD+rhg
2I0OBJz2l9qRtQqNcKiJCgOtT1JEsZo+fwyjyCJHhVD5QzeE8u7TebOpKTUhxx7+
W5YkYzsnW6Zc8P+n41AlYidPlVUJLUMiFC6NnPqPSr3rouR9Ieme8N6/TABOMiBg
rYz5TqmCu77KOIbmMmODrXsoRbF6r13bjf1AcfqA9kpzwu0Kz0XSNloTyH4pgdxJ
+0/O1gNCZXvx+tfPsafL7MhfxQxcZtbPs4sWKTNJqe60X6SQof41QA5kkxfOzQGY
Gp/dglJ4PLpHsGioto9e3h6/mjySgkwyaPlfE/DeTuNlqt4nZEgjmNZsmQ22Gk6+
ZY2uiiahdFOF7ZnPeKqAyXxrJHsni8Gmk8/nWskgJReSyBhDvLceSG1UZ73/7elV
/brvT1MX3PkCjBwLGW+Tx9m61TO0XKDsLCLzqIzjlX3zNsUeUcV2wM6hn8NhwCxs
4lQtj1/1JNWMLKIKnWx+NSdTS6iGZkrzdJ1q2qEwGr/0Xn/iLLynJIPLwVEKlfzV
N1j4co3uS0qX+JG2VW8QAStAFf3vCL/1FX8a5GXRjXiI/oO7JO914tEW0qTcS6yF
0KUKYu1htAIEyQO4ctTts8bFFJG3ZJroFhrZXgJ2cQca3hu9X8+ub/aJfm6BKIXF
ela9ksdwo+TGw8YKaQWbbOBCVe89H9e3wIOBrdbb1DUxEPB+W3v2PAR4HUCrGqCf
1ZI3SobATx2YBYRe8ArnTyLeM6wBdQeePLdNIsMX4Le4n0IqXoN7YaWu/75+EZYr
7gYBvESmCYmWG6K3zGeApjWJ5HZ6/H5lIxHjiXflWeH43Zhy4a+ra1E3lFjVfkRm
Emr4+GwILTFDLv0lGDNsfVxbvvRMJux6RqNg7KWyoH4CKvqIIXAmQRSilULUASv+
fWGMneQABNaNIvJt5CJrrNn1FBKpXlF1k38JXBRUEKew6MltFtrxYpEwkM+FyAyb
c3JEkDbO/y+PD4XKrNYkbqfjcn8ecBSXA2ztPp6a48Dka7hgnoPB2ll4Ump8e+rK
ln//1yy97MtQo1RX3J4SAKtsH3zLD0EFEMd1mFdPcrDed8oKZLuQiSM4YWfT1awC
8CUOuKczcK3PoW9D/y0QslITAX4pmc55kGSgcFBL2l8UzAO4UXFYSG76uAIdMs5I
hFWGMz4xRatXOGptSC56AyTpnU+C0zFT+Cs+zprzrvePIi8fxrNkOeSUW2/r6PV0
cmmOcnIYvxb3QSxKH662MoR3LBl4kDzZu4pqO5/w7F0cBwIhtuBgTG0V1znEN4sf
mBrOEFllGkXWHFjUyZJLzX7bUSylPt8E5UHDAf7YJp+XoxMDVNPcl4Fq2lXbQ9hS
BhZUSYXbtLwEVZfq85r0/K4VLGW9J47DWkOyclEDapmGAkr1UFoXV0+uogABMSUF
ve8oYDaQ7c73PgL74dN8j5fC4agM0Hwrc9NF/v6RC2ufku0Wu331A9I7qX44n1Np
FJXwiQ6BWeXgM9JVH7P3zoucnvDdvvDGPXrhE1+7JA+LT8RZURsKtKfoPWKAAyws
03UsL1bZL0vO83ixzFFo6McMz53mUdCZgMLj9jZdgQ5hk8ErNB76inJAnl/qsCM4
NqfsflM1DzTSp+/LLDKc3F8cEGu7bYUD3bBWR4LYZCFerOQ/V1JxfciUe6rXykXg
Jv9mfonazNnrUIUjGsCLtzUrGUOjRhZBJPj2zIwGPK6HyHt6f0xAemJ+0GHFY8wq
Md7VSSTGuyTzWqYm+c+HUo/tYUazrWlFBqyNIOptP630frPGtVtD10Np1F+ZLtEt
nYf941zicNirKGv5ub3/vIRx10iyaoil8ArvUcNUy2OsVbME5xkt5RP2ojpeJn5e
xvQ4nd0rjXXRirIFSYqtVSynXykZRbdwByCQAVPGO4ELlbQNZxKyTlTRAgX7Q1kZ
HR6z0Qyi03zHp/wRBL5Xu1PWGySCUogTFTG1itQBwKK0n77x0DdBtWSJDSzLCkJX
lY3/S4UXW5XoRt49CeB6t3eTQgzFB42nzSCuD1IR4oeWlvmLcMiHTNgImzPQ/ab/
irPVCigRdtF+YNNS5pO9PLVvyKbLvE6JTRI7ljARXdsMAXqWBT5c1cFRxytBUiLk
StL9K0Zcu76u5/VPLMpteBA5UPp6HE4gjczxv6F8goYcS/y2D8/sdDhGFcZoqg91
nYiWVz0Uk29iHvy8jhn2Ts8+VZYxTvXLTaNlArEj4h5i8B2k6mSPsYyIV9jvGmXE
1fqEJtu2B/+6FXiPUq5O6/jXsegIR0WlWnUi+YFdYxrr/N/9ub0GQQthgsBZP0Qu
RTS+E93x+/n34+EwK8kI8EM7GibfGXp4qaXwbgCebqnhHDOfUaWLqXq9zzimXRQ7
76ml+wH1cYQu2ddLy3OgvTP9b2kuk0AW4Nb+rB+eCKA+ZeBQbWRO9w9d75kPuIxQ
g+DKij4QqMZUBVJDk1lGQiVtrmijx9KlQten+5v5tXwC9vm8+UdKMDoMrjFpsqw4
yKYjxiXjoG2uHQaRK2ZVgp1p7uNo9X9ckwitn6oubmdd3Hw+SVUWrJisyyKno2He
lBZzqSoY84tJp+uRXIiXOS8aV+F91nBeLhQQFjzctVMtVUMacai8kK1qVynzMZk9
VrfLtLIirMkXGpw0iOwH++czvueRXH4ayfTs4MsJNzD+irRNHgyu2q1zHaBjG90R
fCkNLt4UifwQU4+rNKmcO9l40v2cof8PyIpE9dOLL/hc92/GoVTgZ2PQHgEnfyhE
sQzOIFB+PDWbdr2SQivS5SQTB6X2tqL8x3maELPVqrKJFknVeyVtOTKrObWyyrq5
biOilzENXXKohCkl8o07fjK4ikkierBELLIWz2RzlzE/CmZ9X/zSM0W6+Tgy4FVg
Yrt80tUBo6L7wTosCoEQec4jBDCxMl9u1QL1lrhQWwAPF1qns+58HqJ2kDwVzHV8
TDjgzA4mqLHIj+y2knqyBUXvAICemgCtya+9fofV3JSpCuwL/q4+6+OB2RdJc1yK
DNOA6Wa7tc4i/S/OFGAGHejd9YN/Q1ZLYPMbS+WSnHebrTZYh1/2TSeS2VNW84Dm
Z6A/7uawNOPXBeXVI2Gb6v9Q0/8CJhgKoDsTh4/P/bZRw/RQeaZbQ+O0E9+qYAys
Q1V440ftACTstlAgYK59EVcqjRZenWMizp5De+wD79R/W0MQQqp3Z1GhUQ74vGCQ
z3g25QJ9kefkl9eq2soAjbMjhFS7d0sg75zac/52bFXzFRTB/0/1IdfIE7eQ5aVU
Q7x0HwwVEGZ6ptc162sG6FQvrPm/kZgMUAT4sMFTLSjolxvfMOieVoedVTmukVrL
mUFFuxE32X+NEleYGgNsiOzqGUR+M0dG+U7QsbPzY1U3Hd+6NjIDeut4IWjYwpQF
B0U87yEZzgpUdAn/GHkxOeacEX84Fsgvy/KcBM5TPIf6PKlyg85BUn8b4bFzfGAu
RchTSZsVpTzWB/VJSt11z65JJs8GLm/zDggvMtgaf7sHgiN/2iPF9RmiZyPDsenU
CMyhEMFPlxSDqEoNFtCaBjnmcrS31r2q71Fpfy6Hu4PLja9bes/tIeskk6tWAHvo
caYFTvZ+eG0mMu8VMp8Ip2adAhmHqeYhX+hFS27yaTKhYjnMQQOJ3EYcqF4/xHd4
fgVqv/9IynNq8dLOaVSgRdU5UvM7RFC8a4RVIMqG/uJkB8v625Jk13K+donKdwbt
p6JaZ26D/meiwd9CHV8PtU04qJPj6hRCUVASHApnmXMt+jkePXe0VPV71H+qnINL
s2CMh+h8guRKle/RLTYy4vuhcmbYzj3nh/Ji8WYZWUl8IEG24LWkr0vn0uu1Kn7l
IQLh+uuf12xcM/jmQLIzBy6mgX8G1Bg04qPIFquJZ+4GA+oiyvoyi6fOEGMaTqxJ
fjLpYJF7/XVeb99ScQIC2eiA2gCFMv7lRHJMDgfBx1G6yqxrr/HP4S+az2A5U3wB
4lzJkTz5i3AuuGWhMx5cO14R5PNJCGfQoqVIRON7kVnzgINVh94vgW5mWlZFi38G
xT6/eLGDxjrted4BJZiEqUK6Zg70am69v5wi33b6Q//NPnehW2bxe4Aaj6QUAHtB
rdQmfvkgHHeztutlpt7fAMKcennR7pVOKgDMkPAQGSEgYxcllrXRFtmFp7Zacc2R
hSS0/CH2eckTqJ9A2cAVctECC+JNaK31EAF4fD22YJosl0GAlR+j7iJIOnaCYfWg
CZ3IP9TCE1rLFZxPFLSQ5sewCzXlc+vBiCJvmbO62OE2IejWmw3L7MOH4QmpQIqh
zr5Gp3Gr+ZxERw1H5B2UiRRJpGPI9PP+T1D7FADfv6PbnmfQgob5C220kP2r+1t3
qCUZyyiT/YZQvXKgwIena3y8Pa2V6tkEx91ekFAEjpbQurbYFfYPgnkmD0kMrxKl
73TY+b/kvTKIrb85ncJTYdXY8TSwqvX6biI3xst8piiyERzOqqrqPhyTqeFQrIR6
oAcQqERxazlqcuYU5RAlOpNiQ+CJ9o3EQEGK6u9rIccmvKzhqeCSMf1paf8pJawZ
PHYIYDfiQ+jtenCdeE5DS/J9INLu5n91LJ6IPkpXW4z01eMrGC87zbwq6hPD1m5M
91MtQ2lMWK4Dh9YYjXIIt+kMzpFcBDcnhC7kWjdyoE69jGtBYqXq0Vc/+vOaw26j
kEHkR3FIPwk5fbkip05OVhxyeh8YfsjaunglznWmmsHNR91luuNDz8siuqD1jC0l
wttjkj+vddsqvKK1uZgBvtq3B8fMnu32tArddnLo8gdPPXTWqi9mMoMLdY9/FDXb
xjJVuVxnR0ud6KKyCdamuNNEWi0vRCm8tMefjfInujKuliN/biO+l/qgmumm8CWG
qDvt7KhDxyDuDHHaqLzu/hXgXHeZTLXImt33El8LbLUwlox+Grv3cu6RMzC5rcNi
ForFgNnbyIr7gAZAwQYgs8tNQa5Tg2R9Yt5uJT3ck25nPOV4ApKCnmOXZLKQdGtz
ornNmPOLRriVpuyl3NalymwxZ8wuvsutIv0/ws4e+dDSZOFEpCZ0rAynD+ZqVvIA
YUaxOCbEiUdWn2qiL2zXmP5vztoe/9kiy70i/bbxYolpsIQHo1tl08Fssp+ggPJK
Z7YejmspRi10JcuxIUCGgWt+l8B1HVKhMUMxDnU/6Lm6DiUAytv9XDcyZ9Re+tHk
G7SiFD0sARMrBGxrlFlA4mu+XG5O58HmkzJGId7RBp04FbN9v+LHPlPr0AE9lWJK
Nkl+PQ6aXVIzmCdeOWez2sJei8dAXodHIHOLudj27fRtBrMPx2Prz1Q7wyxIjhZ/
H8sCUSU+yB70ZfPhm76I2QfPM+l5dbZCVLrLuOQIB59dXGnhWWhAmvTwln+mc22p
ts3LtOhzViJAmN9d6B+ziJJJtqfIEcMz/H5npCz+JhzwQWY6Wgo6saX1stwAjTZ0
edmOP/YQN9x7iA+pdSuhLoPPxSaPPVj2aaDol2kBM11dved73Z2yNqcUVWREyu40
3xQ7H5tys96FrMEn7xAm1TF7VoiUY48k7b+TCte7cEA62Mjx00KwQxu2IqYbzIm0
fL5/2G4O0w6SBfr53hcIJi1jTy5RfLPZBISQpC+pwx7zyj/G6MMhpns4akghSXCP
JhH+HuVjpZocKG/yl8riYJaC62nceyuzQSQ27O+pgPbL/028LZ3RdYlXNeB8W6vo
uLLeBSrrVDDxDUNgRrxtPhji7/azwMb5B/+WyN5FEdlz0PaRP145vSmXjWMwfa1M
L6v2NqzOeboGIr2AvZ+x3WzNZxlUYK2qVZaOVi+4tLCFNJI3gf0ej5zg89hQeIKL
VYTaxHWatIS7moDxIVkMcn6N/nO009EM8Kb0u3K9x+37SBsYkCPQfCcC32DbzvYS
8oR/vcwNqPLeBR5GQflimX6nMVu3W3KNVH0clBSlH4aM0YxJ+fJSu2ZADELIzAHT
s8dpMrMrylnqPSvoDWoDijwDjKhN2U8sbhF+D/DwbFRdCAr4xvjLnXSpFaGER1Z/
lTrpB/mZYRxUqMgCQyLaUabLNsCYC/4uAACmKsAhcm78+gEGDh6WGo+TjaVuzndv
CmcjBk103PiHLBNgO/iJOOJ7i8PpCeUJ85P3XjMCWSBUy1yZEcnq6vP0Q5TAlnoO
ep/UOjW96glkm1Luy1iJcPJTgC5odbWRRKlm5Olqi9lTqGnmUPN7dVJI9omlBLOV
fISyzYrGysZJW7rLmjPSc7GYJXLGXqZSzxpQgYrse0yYE5+IeZv7Q0apcYF2r1sa
7LyR7MA2wa2s/hCbv+/lRsEQKOPAY/RmUTZzuhWQg6LmP8tnJ/XkeuLRvjTgpVuf
shpPKC1y/sHCW5UNkwJcbke8sNqUydJMRyTzlP/mh4JnOXGYCRTG1CauqxjdauEJ
QGypC6cfyNxNAz3TpHUvaFy3crtSJOGYn9QSxnu2rxLVWdcy8qw+FM603VSAJncH
Zj974a5LkfZJ13l5YQoWvPUPjPCTbvjh0pIfd07CrRNWoahDJTtK/ZDcM9ZPGNRx
GCG70A5Ku/d31JeO8xfIW9L5QSe7KNsSAuV9TzBFZOMs6C0AMMT/pgQ2DHorPbUu
HARbeUuGtHAuzXYA1T4tIV2fE/WrXssgqyUgLtq8ZR4pFrkU4uiCbhhuAHSDZkiK
v0i/s2WSlYUTwcHOIu3UvA/G/cAr526AAQvDwKoG8XH0ja1VhQMcZ3qlj6Xec/xD
RAMW8y9CAHwuiCgoXHvhPxh8AWmiK368zYgAauURJoo0+ROgZzH4IOtYHc8faJiq
0wiYXiOyypzFNOHyP7oZs7EVJh4H7/YEJDqEoXxboyuWB/5Hc7AEmQTP1K6TL87Z
LPpb+a3IIuOuaxvtcPBN2ZrG/i17qeUuuLjlvCkiwosNSNgQT3pzWIZwrD3FayIe
BDwYrpUPOWPyKZOieySCMT8ZVi6AC6+7y7HKTASmU8Zv4WYrhN8Tf83dS1rhBqQb
OIrYmihy9Tjpvrs/Mng7ERNbLaHoB24IGOT4XEeyfvwkaAKIxhHyN3fjZZ82sxgc
`pragma protect end_protected
