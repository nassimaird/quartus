// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EZyM789rUU/E+IcfGmGYk7JKLTVIKwYS+8qRM7oCKHgSMmKyMK3K8RBSXJJLvXEsGnS86CYFTt9L
4G4JRgAK6dxV5jr1RQTHZVqD2Fw78H1jtx2okOofSTtKxBDxjZYRuPWITUz2EgQmoUffAFYzPtr9
e28OkZjCG/doOvigi2CPqn3qfTMKE/pxedpoQ/EO1emTW9Pyw4nObZ4L8xIotsei/ntR70qbwB73
7lXyyqOvgDF2At4kwNDzqjNnqfqWRBRW4C1i8b8Z5tb8u7BAw7nuNChF9i26zjS3HuSgFvAN5ZuG
VKAX6Pg/+0weROJdINxliiDZjJO6F2LgU/Qb7w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5552)
fHsGKb7u8vNV8932wDSwL7yUOFmQ+Hh6xQwo9gy2/u+2bCV7hYQR8RxsamRNplALRssWa003uSac
Y8uOcbipwtPGRNX/mK5FNzd/i6r5Hc4IH/jdeXXRYpFN2rzhBmxW7l4LkKw1TER9owZFUPtXXpo3
ouP7zTO4nYPoYhe+jT1rb0GejWmPYYx+n30PzakY1bquL81ui9bGovORQKUDF+a/3de4UL92d/RL
ZcEN/U0zqABd5p1Xv9DUcC+lW5m/7W09MI61eU7Xxsf5rRqkx05tiSABVwfJ6Kjaoymy3PcP5SkZ
N/YgSagCZZnwVU6vEkRMuf/z5riOAlKVAG0Y3Y+teGQxNBWtQZGrKWLHDpLK+mpRPH3v4r6sguwY
TflCNg655Uj8jT6RzVYts0j3IJQAhQY98pquuSi7QyLj9UzDs/DqnYdbIAJRz9y6UhLIuirzAgAq
Mq2XQyV0uSbZvLVr+bM5pFDCNVGHdBUDh7DM0Q50veE8Fe+sT0540p4RY9WShmLq43Wft6bljn0N
v8p2casxYBFQMeKGTkT7LtHguxyKhFtQh6tEjrUYK36tDyoxXAyMZakL8TU7+EYyUpu3NG1k3f9s
rH2R6TrB9yr1rxlBybN5K6j+AjaRBu4s7dXfSm0JbuNFcEsIb6qnseaSJQZqLO5cCGTE2MC2rxBK
q0F+ho9P42d5pXWUd5fZWpKYD81xQomYWQkhfMoh0OEFjxmt0GWlzaFLx9u+v+4jeM2Uj/ZVu1iq
1eeyPsTZ11BK9vMT89wL51iXbcG3zR5GV+X+C03t7uYZmSv9TOEQoszCUPd7YP4u/4K3AKph+RDk
gx8tap6Leew2CvTyofUENJq/4sn5FbfYL4ETtnJ4YhXbfffMRUHaFkdnCIOys+WHQh33USl+JQYO
mglEwAfyehs21tCh4RQ5It+WH28vNISuBxJd1qL5AY/ZK57n3BH8dzouP6bnNOo0bwlitWpJmv8u
BNYFpR5yEJfbr3QIEsL+VdUcYQKKFFszeS+IHLKJdAx0Bb8GCYxFhdunPbuN4MJyb/uAmCew958z
Rm06IUummGtVnxvK8vTbIl5lHqiA3m0BAfKW2ELM/pj919VWnr2Cq8cXYdAhoYeqI2ity9d4OaMG
WwHAEewITtgkzMYOd70jI483rtpaFQTQaLWDRk0UglRZZN0zLjp+926u2256aC2NNr9thVbYzHMj
q3QwqetZABW4yItgwocB542Fv7m8RgGFMTTcdsHOJZQO7FhSPiGrDnz0bkW2etiDeoxbzmR78EFQ
2jWTognK4GjgJfxXruac327Otpgd2/2qatefOrSCUMChVSCI1QEdVqGC6XOcsF/vJ0JSH+t7nkDR
m6RCDqyZzYk0tk32b8C96UnNg2cDbJJ5+Pi12ZkksRX4ulQC/d2Mwhkejl4R2eMAEGkYCvtQnoNo
fl2ajbNjMEzrHmwCyNR6t6qZBf3crrsUpjRmSG+O0765uJNBpHys86UDzHU0t+mcFK3+c5XROLqq
tpFbKsSECmh08Jh1y2HR2FBKvR6sjlvtuTbFTfiP7yNF/F/+zhwGiCoaYvY0tfxmwyhlitokynqv
wEj8rSzqiLlVWNi7OPThSp+n3MDF7E+fchLqz8hSH6RdbG6BEXFrBJtS6rX5cJi49ke+v9i4uV06
8/FYenFhvWAdpPeAOW8l5nEtlV5qWvlY1Fh08Zag+wtqPSykE1lDhz1Jf6PsDN4WGnjd17lSmR/w
z2Izv6eAhmttU8Cj8eB/b4cDkZ7h43Nl2Oj/gonjVkBEE3tP52SxguJ6CXK4UKoPJ/eQwbzbPA2y
FJsihsBHbaFrFCub41Q11TViKCugBaH1BNaPd10zZhFntgof3R/KBfvYRLCbqXPYtAYxZau1nP7n
vE5W5yDtByD0yked5/XjooKwMEDaOd+jx23yXef9GDXdm7QBLGIMoRMEkgZkObGifrGCavd/lRhX
NS1lB+a64KMTaPrhXHCFTojCS2FeRfGGiXRYbmtwmjmMq+zPNCIkREwMZ0OeQ82ubQ9V46OXlMdu
Xr4W/bBlw3JkFynEL2xYocTlsixblzZvqXeR3CyduFYva6R84lBsNg8S5SE9S2Str58V2R2dzWIQ
u3EK6g5IHwEYrAAfU+wklgZwrm04YEkNHgshZIOHz4I4BY4pX42DAbWzOlV3on18N9gzP5F3Y2h2
+UFzxNaDkMkCN/Uuz40X9KgS6OynDkTlDzXUNYXxc9c2CLHajucArr2LkhpluCllOX9falNPM3GF
JwRUvlu/HlMs8ygVr5ocMVxijrJ4X5qbb5KCV8Eq/s5In5HY/JaDBy31QSJtQ73b9sFH1jApev8H
C3yuK9PHsthwp/A4n8UFHjniyVlDytxv1lUV0+IW9fBhGgfXijRN2rWce0bfXuX5YNmColpd/Tff
VLzW5qrcUVmN5GmW6vzsXZL6SKHvmkjsX6R/dfpUUFJkfesVo3EoISeEhkx/bRlsTeLPqATNRfkF
P0+3EhEJrFKmYuCjgVtL8YzQK9sf6d976HHdpj7x+Ef5ophQN27iVujmQYCavVBHJs+caVO/gZPi
EzMJaDYqZAGO4YknbG1OB1jSWeW/AGX4bEEDzGhCINHWl0khqDW/snryzDAZ742YHlp9sIC2ch+S
aQzimQLh06pvBejhEfelrMVuxCBPsgGELcBVBh+6XlncfvfYY2EQxJiHCMb9yWvPMtyPRqjuhanR
VO7E6iUi/Isyv6p3mDPwvQwoUFbILhvce8e418AZXKWqstM9SqGOjeIMRSqT9594TP6HBcNNpfPW
PYylVvuMZBnfAdPNFiNYmqKgotXE8Xa7UYbne/xEkTdrrK2N6ISi6QYKeNpsIL7zyVKwLPs1ooFd
2CfvFE1WwPBI0yI4SkAvAu2EOj9YDynh7ruPW7kfvoo2VORz9eWULIKnGYHL1e/pLzoCX87TbSqA
IEFxany1NRPM2m4ery3g8Dcld/uhYcYQm9oMuj06TnTJWeiXZFJAbLWKVQlOpXcxQjW+mytDF+pw
3Im0qnL2UBP4oauHfHl1z+kwuIOPmfkXquPemYsFHcMyhxfVvmALzwjFQ/J1EgjPeEYTe2RiWbpw
qWfoj8H2G4tFFiPvCF1az7tdfb6W95TgitOLk92TBZmWFho/X0VXHp7g95ZOFR3eGN+z/12pnVKD
M2dxBQIg6+9WlAVDEkP53zCZ0NJ61Sp41c3quImqIDDYn5020FpC49YfbebsVGFV5eGZPH3gxMbf
2uQ9dr3qFxIHX6veZGkfUeBSUS4NIsOFnNOlwGmGyMXh/uzwGzENyMLoopfwGNm80SffIXfGaIK2
POr+TIOOKuM3xPQx9pEgIN3cPW4ZNbf76XHWJkRwunIyTscqg63ezDZJl5EizKsybVkScioef+m7
MoRdEZudVc6ZnV1vS25c2KWbD5X3K66K3brsHMjmZU1Xl/XkrrrY8lPqAK4/n7Q5SKlJASP6esBt
0SwQIolhBlCoIF6XvuywgtCqT6bjvnxv8cH0SAW1RDQKDf0veaQz8WPKoUJWhU+akLQNEwyXQzm6
8Aoc5sQh5qnSCfL/5Q7dQTUnsBgbfHXR4kapkJOILsyfZuGkxFwHK0/bSRqS+9TaekK0lNlfSIyR
04B1ef1VujpIAUEul5ZmdEI1yjNPhvpceCwCfPlWmUUi5afB5MC6UKUjXf4Us2glBXz9aVKvEQUe
hVTDoNdtLBP8/5qnC5wQiV95SJsZpCJDWFWPOQ3MYFQoGQbRiwJ0dL/MMglJFipJ/a6xxZvSCaKm
zXb3lzSQUqme26yKOcsfBotNM0oXYH0X2Z70zERxmp42vSt/HKqQWxcysJF416el00OTxWMkJDcc
OlqVUeBy6Vh035XIxOwGFLLVKXlwOOeAuvdDNetBpHnb0eGuOn25qhgrWh6t1o4UZY2Hv2d0VMt8
BW4BzhKdijRkDMFdgV+J5kkYlh1LdTGLKGxpCJe9bUEAvpxyl7k4sL8aX/T5ww78poOP/CcpmCb/
eHeAFzHsLtPqzqVlavrmjcMm/fSHHSZj5RNNpC11K7IAFBJUOgIoS8YJun3lEXL2UJ6JErtzC6Mh
95I3bRAD8KqP0RmagYkH1ujHHgVIvBKIwLeoFI4gQtnv7kWE2Q9cFtYY0KVwcAaKveTS9T0UC1gm
Oh4cG5tG34VQLZ0H2KkPhxERhcVGCMaE75pLWAFfLmTB4HzUMOGKl/JZJD1B+hpJFxyvfnXsDR2a
UgCzt9ph6l1iLcSYNIEDZ/+lEr/W3ZEZB98csq5eRZFx/R8YaV9jj/GSZCEbIox/6BJQ/gKNQCKU
wmtnitC/0kaafbHC8vFIrQaTM7jy1D84u8NvJAXmRXPNebs+P7Zp9TeGhGUBx/d25BmyfyQXYPY4
YrCWikEZuM/6a29EiI8BPvAwcaflGr6kX2hBGYphDI1BGbcbbexzddD1PfDF6t445VrQJyAuLELC
VtpFu1WEbr2EjixM0SnQIzmgRrzQEczBrV6wsP6Qyg1CQ9LmW7PSV81LKatcgNpOGpwXDvyQ+YDK
xmCe/5oK9GV9yBhHhP1DkELOaLTEDTjl6wHW3Zbmm/Dzh9SwIkSa+SKtScKePXXHHPYk+rPEsrnb
ChE1YCItHNv+ty/AOPnJfmqrBj08Ac2PNhrowxaBLbvkrajyjdqAi3oELfyQtW3EgprZybfNMsPZ
RO6pq4J9HL45MxTBmQ07CcRlEBA8f+uWQcGPoy6IhumGQc3FfuqzASCsZq236sHMzLe2j/AXFrNO
hMNXxGx5sTa6XeQbdtJP2mLKxE1HLw+nzwJeROb5Oiee8QFNpIRAyeL/V4zVP8/eV3aDh+xx5/kt
QVN14WU0yRzEqnEjyPMw4+Gw3iKvTjgpc1LDNlYUmrKd/8TCtTtyZy+nCqGG54j/qkdhXCd4tQC/
UPisjhF+z4+AsaN1/MGCI5IjZj6W2YW8OBs0y49cvZpArRPyg/gVVu1ZX7yG3Ef1zeOXX/sS7O0V
LBe8L6me5YkyKqdbX/P0tsoLWqwo6iMMpZZSqJiEyosiroZaa34WzTiwX+pummuELqppxlMSuraQ
qQ7OaO73MHaHqQ5RgkgRVcIhZ4IIh2hbqEo6RHsvHeeXQJUoOvXqOsT3T1BAdV+f7SVSIH3Q7e7w
+hCJamzNQJigxB7rLhXV1upgMFD/HmuZnAeKxzYYfjbyCl9aU36WOclmzOKixZCXfx82ON4I6vhd
r+SCOMQ8BdnjHzeLEFRlIo8pbY6fOfAJWgvaTGjjmVGUkUIoSm3BPSu2wF5Ol91/WFOUsxM4RW9S
hNRGH8Ptk9amrgH9nrmceudtgBDA2KSvTv4S9Av29xeGiENYOrbY0yiR/FF2mI+HHk/8f15OEAtO
Z87V30Hkkjlihmek4lXJu3IznRSwHGdIxInU2DNEwlFfFUQaXi9BsbiIJCaj45M14n/jpZKsufy0
33WmktpLnPK4DkgkfRKqoof4X6E01wxix27iq+sJ4I8WefgxTdWWG37oOZGaARVv51CFXl35iMvS
+1EapB7B2rdR3/tTtUXXAzRuSdyrrrZ0kNRjNCQz3RE+8l1HHqSTyCIue+cgFp0zDjaTcTpLtUyS
bTbU4JiPsauJ0kCRVJnwcnP7ODCo//t2hJMbVJ9L9/X9P91K0F9SdJrJBncJjpTLg4XnCEBh7mko
KdTIVvzOqI2vHdwhsjCVyAMi73tieRzcMJSOKJYmYnr4bP52LZ9TNxrK+qHM5eLVyEZRla2l+UWA
HxPp7UHrSZ3KrI3bOQQaYL57vFY1pENIo9nB0Pbf6mLb6TU7r0zH5r0aLBZUX9bkQsgmrqeYzCwB
+xafVvWGuQ+NMx7+LQppnFcHyJbvr8dMOVYUalsZDRSaETKroe4m4AGWKIdchU54WZQhzc0ZGeDG
ZvskYFnhSSBgApfZLTHOHugvSb65wacNfkRro73NoV+HKqP2bNTe3Mhxj9uR8efbHv4p2K+LvJbW
csW7tU52bzpCuPMh+/3edxvPNbEAsJBLaXRmkx/iqbnQufWr8jdl5qD1BgK0Zy1ICBIWOkUWxJ1V
xZNFo6LVbjDSrJh6bNh6mcI2LYcpZI0YiUTY/iWGJbyWAJdLVTbtWR9er3CZBVDHesG0BKObowKP
iv4Y1e4x6LCedLUnbNceC56/qcEZ4yKPKKO/TpkazJREMvlstkb6yjwYlp9w+6wS4NeZFz+anLqN
+9pjV29I6+oU5fL+B8B85rlRRvF/1iFqyiyEGqrcDnwBMQYPM78Fy1UrGt+u9mqTxNzp6bomxC4v
1K/O/NlfmpzO3QTwsT3pMtcgPwxhrTv/buIHiTeGUYO1P4BS0wkT/7cF/Vh4A3byFljIEEbHQsaW
biBOVUUBlNJnz1bYyG462ISmybs9ZSsLShu46T9Lia2rgIhYnOfFF+yTXKrppFs33hGt0ikk28vh
v5tNWBcojoGdx8XM2IyRrYNatj+85QehczcN9S+MYVLB50fyp5zSDS2neKZ8PnjCJjjca3jPl5YT
HzhwmPYiETyRrUSRd0LrIuVFShu/vBeq/I4o7IknsMvbHr9/OvjzmW40kgjeJ09kv4vdmuOMlUtq
ss1f2AbWRgkIc7S7qtzjcDgUF0L+/HQYYoFdeMZ2sZsEHKx1aVb4P8nTudSejSmfAMzyEzE2P1NK
XOCsWyezUuqt8e0FQQwVmhxJ86NrTJvf9rm/jSjNlo+I6ZYoK79BSx7HO2w19i67m06ucvuU9wbc
mqK4LfcG0ik9yBZuaGS8DTkweCUSTtIbVnVBBmRBeKWufQ/nEd36b4QYjrVR4AMZhIO77DA4LVYY
L97SrB2uPfqBvWX6lK564KGAXHSNVYKS6DYvbjmJ9WNbXNMkQNwnin0/2WteDbIGvhzEoVYeEy/8
c3pq+7OySvn8CsuEGymJIPa3GVci8LLBdIj5+Nto8T9q6ckexlWk6HZRhzACGmAW6/Ix8le1LclC
g3Hr1dl/YzAYZfIg2VbaELiv57A/sSB8cMRU4J09uicPMVITkA9kGf3Kh0DYF5GizVABvLRXazae
9J/XR1C2ZOB+uZnxbIj36jigoEwrNoDbuf8HJq2JbCYYSeiI5+/4SXDJ749YYsFmUQ/ZX34mQ6PE
DuGdJ7ug+HElwcQoXhfOqzecjNpiDn69uicskdo/E4SBsPYktSX6fydXW0nY8v9JTJqqYDWp+xII
fWeoC2p2z8L0WFoy7xPOTFK+RrXUfNPsOgvf8zVzZrHroI/49Iso9H228zPzjYa5e49WLlq6nefW
vX5RKf9Us15mOsynBIKUa/s/KcSGYZFNKxbmVs1+d5PkY7FOEzIGq9FGaG9kvM4HpW9mJFnZ18DP
Ar8FUyM3wOfmCpcPdFa1yqBT7+5a3m0=
`pragma protect end_protected
