// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ivA53R5/C4+l7U4eI3HF632xYBwAmINwNqxL1hF19B32gVQhlgNAsqKJ3qbCrHNzuAsZhGL/yVV9
T3qDzWC6QlqIyWhM2sCbraVaUiUDTAG5Zw8qeQ7LpDFx+IYFA9PEp0FFLGZfGiE3dihYkIspyQvg
Y6NIhNnmbdq0wSq5WmkcS/hc6lElopb/xOU846Ftk29muKVORcqS/2M/SC5J84WTGNk7AintAq80
3/Cx3hmux0AX4az60m1qoZ02kgagRHvN/9HflV030SwVW/swRGaeLfVbPiKlVnyrhQhra5wX7bc9
FNUBsBmScgnmliHk6fCFpE2zcLs9eJsLvGnIjg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 67584)
PBtfkqMIonOx3k1VdKd/NHtU0DSLO1/1V/BoE9KsyZJVFSaBZYvFCUIainFC/WJUKGT1FRaEov2M
p1/yHTDMMeT9iLg+MEm/5OVWbdnPlMAi7X7L8NlNlNONFJwFm5Db/hYaNDOtFNcniMKQ1AoPf7la
87u9rf9ONolMb+nQTnx79uT2M1ux5Ccpf3ucRwryyz/vWJLnWc++68SGXSogNIXrPv8ri5oKeysr
yy58nJc7I7l5e0NYgYQQjokSdJmGSSU+TT6qUOHKPau8pTC6WkoPeWX2Mvk34qeRvNJT5NGji7Jy
wGNz4us1ewnoRE3/v3PMQosbo/jEi5nme6KWNkVY78NRZHyGYPHMbLXyZIUYhRM5kWlTs3k3ZPVv
h8D8tOetYuaelcq5+Jfsyrc2DFmO++CcW4lI6AgKHJMFUmS5XMRUUb1XZHs0qhQwp4U6sZ6qD/Hg
3g8HQ+UfEQp7juNn53SQMJQL25/fh6JCinYYMJNml2M2TlOOi8AUACSnqtTnmPvHGCUZf7V+cvOr
CF6sjLAXoHLHMu0/0FhoXyqKMANpOhHBv+IXuf+la8ZNDBk0f0kYe8B0iDmp9w5H66XOhAq11XNJ
cA8V0mWCqIN7nFQZ7PJh1LuHPwQofd2GR1JswDPLdTrWrGCJjP97ayfGdit6971/nfJH6iOu/1Gm
6vSK/QdBipSolfTMKjiID6xhCRc783yfm10a9AFEdTvErjx/CigYsP3MC/fb1LpSUlksTxkcgjmT
bvvSMvD7N+ywR+U5FgH69q4THBwk70ROb+lrcpQecwwPSMjewAMxRXyEZd3+4jixvXej8s349mlM
cEhohIdDZxTDTds3NiavPHyw2bFyZCp7vjXDpEd0F0/0AoxPYPO737wdJ0dLftODWbKLzVpGRWqe
khIN1fbzou5JfgEGyNz4DK/kR3IYgtK9KnhREN4cafDf1TqmK8xNv82f4+zRkDn9rrHqQ7ZHXfJQ
qMznc336NNFbMUyk0a+lg6wPeIpcgjs/vSZrhog8tFG80jlZc3TmIeV/Ir3XlMo1eplJAuJ4PHvD
NrqfGyAuQUBr8xJoSCDJTzhBkZMWpt3N23Sr86ux2I4H0+FZkxbqq9HLdLy7hvmqsA30ZnQHgfZZ
P/hFYk/s0QfipFHECPjD9Q41Y24nojo9tD04A1Qy2qvfvO3HrZlyK0FmpLcGu2l7JvljfRC+x76y
2HScWnIjpzBFnLFW0dxn+yQEe9/T8d+O+vJ/o3YCXJRfNhVKFdqlqcz3xmHntRykJIVRMQ/NIhwE
EX7qRHkMZ7mJXLhnPgqYK08q1zUJ8bF7fUaluqmBMVamXxnMUbqPZtFxOnqjFYPWYBnjecPsFTwM
eOt7ySe/pe+BEaVodnMXRhfBY6YOD/3Fq+qf11sXx4QcVETBHYgvRH8O6YjnqE+piY50Dfvdvvhp
jVFmk5MJGSUHpSu9vx8jicnw8e4Yip7HCLXJX99HglMWpYkMMxrNo5LLTz68me7cfftT7daaRCi8
RQTpJkwLQUaKdeHrQOzkQnKythAW16KzEW+Ey697R+BSLRlIP4qA2acKliSeg+J3QVNvLWcaSA3S
LeX4cuHzcRMdRRd/54WniNc4iGlUzg0lPruvnNYWC8Y6IqUVZiTc1mCC5VjQ5GpnGcr3KfK+qFP9
S8wseJpM6cmOA1JbxTebyfj+wUuJORvCJQKCIyvNaThW47dqC5bVM6djkzvql5oM7q22kxUgG4A2
VeA5EZji0O+oWdTaM1xGTcUlsPQDdWQUcvps71ybehAsCsxL2F1lviWEw1ReQXfE8fChBwF46U9e
EYsgai+VOLr43VlG0DiWnXN9t41J8afkfDAvJk8oFdBgeBNx5k66peVEsK89ZC9slmbcQRmq3yAu
uA1gb/+zrfdhf1tyIYMrRd/zSVcnLvBUZJFkqlWOJO9G0brTlrh9LEIiF7epOph1ruzplwF89YV8
TK48w6JxljfXhhaCl7U+uTEj4qBxyEErn1GI9r6zW2RRf71bx9miP/8rfI/amDJqDiMYkFAfBfd2
VEAlFTgDscaoUNcmnv7/9lox9dF2ctEu/HNWEdmD09iFGyfS8YMV3bC1ljbBdn8vWNSwofYm5Hcp
xkfHUwFBgYW0AgmYexIfW17oKhJq1oA210rXdrH5+0VC0Jc8Z+fdsga42roHIM7pNK+RQ8PYz/9B
kM7XmyEIOLWePat7j5G79r0TwzCgj6YKa/dB6yQ7qqyoCnqAK0D6jWBdnWPQpwP8ubjlbTkA2pU+
y4d4wlLfrc2Vb7W+RTQGy3JlkuHcn4VDRG9IiFJci0qWvfTFNck7n2FkPCcfZNM/Wxzty2WuIrPP
NyGL6KcZiW6fLWeR5GLYlTpAZ4QJnxqvyiGNxuvm9EnSWWkhEROArjbfyq9YHyJ8Pm3TVV9LtBS2
VUPd5gl7S2d6+Z619g+OwiGyxJ8SlQOcA9CqwG3UxiwcMN4sVSg7AiysA2enkTVxo1yGTt+2vOSe
zQ66zfs2LvIXSarsaaSlWF8HW/C9acNoQtRM/ND//2OaAXNbcOsdWUkYv9+vbBjMMJiVWuOKhaLN
xpCc08j7NYBms497qaQPj0l8K6hniT7fpkXnkhCJRLwz/U9lmLPtJZgXsxiFSiY2943LhL3bAY1U
vzZ+hF4A5KpD3b46YN5V/h7LROjSEiMm6St1kqIff79SbGh3+G/P/iEgCvYJv5uWDP3LRmbzqB8M
PkXY84EESjnGx0UhyIePJP4wkaixzHvI8IdoQbJkaMn4/ZoKl08O5myYo3kQtICw0zF3tYyglcG5
rWp33YTk87DWLo36SX2PRtJV1VIOFVnxLsr8sXGF8w5jJ7YHFqkq8IKRLGUHtoxmwb2aReb6PAaw
sNyNgHBYr7eNwQ7sPZFyx5W+dK8FsVCaix6Phcy47zt0LIoerBPbscX0I1aXA++06RCvt4U2zdtq
mIfa7uXuahe/vIy8yqVqJidWEIk+o4Dnl2LMfb4ZJ7h6C37PR6Bp4mFlclQMmRrj+nnwEk6jV4tT
iV5AKk1p4ytoUhNcZAKRHQyKFzypwkUVUt0BDmurXLm6sZJd6RBPHXpr0DwT/lMJKAIsv2gEh7Lp
Wt7enOYI19q+knxk9zipkpc3KrBsfRB3j19nqRpzlm6Y1gQWc1JAafI9cHeaJ2aeAE1nO8FyBRgl
UxAjE21fkWkAlEQRNmG3AqmL/2VQ4Ayy1oMWplR2aYN+3SSacEDZSAY6PzaRhqgeyvhyhpA9JCRR
uB+pcKnGv6z/gEuCgE+Qjylpvwl0M/CbJSB9zSW74c1q8ZFdQVTaIRcKYNUOE+wayyoHgKoKANEq
l9BSsjQDvnlfigzKUHVq107rHvAA8I1MBm3FMTYKN5P+No4s6zORxykwP1BAxmvBUejcGFFksb/q
mIDwPuwDLORLlEREnR477iSjnzQcUsg2X1AWQuuLY9Q8x8qYJup+M2701yq2kIOB6HpoJL7CEvSY
lWkQ/in+TfsM8VWPm86JJctZjL2D1CX1vugtITfSFMHYiKYMUn2fSGt/ztIorNSlFzFnIkXWZQpd
DxtT1GckBrqO8ojZHxSjfGcwOyHxzOlsFH7kaha+DWo9o8lF6O7nNEyqmq4cJinTI2Ay5XEYUFrw
LvlLRikHrZ5C9+cQJVbCOlsmIrerNnV+nZ7nzM8sWpMKRj4ojKHcTSuguFgG5eBZmlJGkkxVCaHU
b8jo1Nlm5GHjk2tgbgzu3mpiB+NQqrf4nJ51Qb8A1BCpPiQutkabeuAI4ykrIK1rbOTmeQTfntMf
2gAIezfoGyYsZAvoXcW4rLxlFTogPHZE8KeNKowk8I3AncODVPjYgrg7O+++urjoRXoqXU9OTTPC
Ba0M6bd7g2Cd8TLe2fBiSEV+UzZ0ysOEjCcVImzCIgi6dcV6vIPbZoGBbjbbXZr0FaSFDZ3RPRiw
OFAo2vAbGsUgxpRXDjOFy8d0Brrk00U8rWfVw/myi731KeEZTb0TtuWQFObIo0Xbk3Fu4DrESGWm
rq/IL8XMNuiGgjeAOhZpq1HPtoxzq6JSjPHNrKlQq+dPenbozWESwK0Mdb6qFnSOPBTlnEjqAs3s
4eT/HBm8dijI7atHchtvsGWkkUzjWC88w5o+xGYPy45SmTX+a/c/ie6AigIarj6PNwA3namql222
uPZv+6CjfVVzjF+9AMqMdgXAdl4ajzFH6CNWl9lMP+kzHo/HQn5ePeUkCLE9bXB9J2fkd03SQQIL
TOESHBW5F3GvddqsUIuKLaRPIsv6Qa3NpiF2CcBpUo670cb8xY8EB00YkDiCnZ4JUNlVzpa7sP13
4CU8XybjzPVqrI8vx+vQjylqocoN/MC00X0yO52Y4JNS7q+eDAhkgB3OQj+sxNyJXekz1fyX6YEO
vybU26Yk2UJjUwPk6wizE6KaU9GNp8Pa/ucq9CD9mHgvDj0idU1k3zFumof+Gi0wEnaLoff5XO1j
0+KVxgQutK6xI8W3v66yKBWsRzGFneJBx72dno1WjuFGYgt9Acw7X+TsG5hUuChjYDEuDSocbz4b
Un2pM9Ja5xvy+2OfbeadviDtmj5kYTlHG9z87zfw5f40e21zgbjaUcuDMLPQCEGl++Ht6Q+2FRiB
yX5BOGvtZF3tCZjw0oxY8smoFEHh4vXcxI2BKVygw/ZjwgHZ399wrEJGTc5wkJuIhEMIh2zkjvqF
On3r43zMqBOCuK/9q6iTtx3SlpKYnBc/huDayEeaQN54kZ55Tqn7YEvcc/wZjrjpy2k7blk1/+tb
8UO/vt45aW52+sLezI3FfnjRsHzYOQD63g6S7XQRcRxYNc1gvUsvNaVSK5qx2Shll7D06aCcsaUj
I3imeN5SaS2v6gxhc/dp60n11XOHZ5LWQiG8AhQFcUCVRsQAP4dDPHrkzD0ZymzedrNxv3Lvzx0e
co3ICILWFEdMzWbLvWl/rEZSk0CnalD6CBxpX3PitFEbPTnyRCndWn/kFjqFU1avTfSF/4N9ASWM
tljETB70lZJVtGZ97XsUas2kK8mVfHgDZLE93veFf+Mg3zspR/ySgRPxHfm3gNOo1ms/36YAGkGp
5rfn2uXXt72Egeci6+biVTdHBaGocKkPVDOamOvNp+nkOl8wjsy9q0vs2W+BfNO7IM0uKfPGIm7h
V3/pLFcfuZwua5CjgTqbedqcab0cbEZpX7gbltfbkMWW5UOELB9QkVKZy4lV03Q9ry/DKvWfJPUB
Kz83l2j72ya/77JP/SWS0CGkz7GD2RKLWSsWaZD8Of7Rg3St0nMQQ5C/7NglsulKVKtx61hj2rUb
Fa1+MQ1YXHzapZ9iVfq5QzCi2xXGUdrdj/gMU+huoJf4B1Aiy0s2q/h1r1bo6X3YvXuuNbRc5RUY
2idQy6bpyAnebLr8f7hOmjdn2DLF9ZgeG4X43Z72u+nDbd8zcBRvHe/tkDj9nFQZjCGij+nsfxje
UIVFZBICq5qdtPf6y8Fam9bONUd7dOoWpsRiicQCvSiJIDrvC5yjtF4X5Mb60hDPRQKoAUkxeluo
nIbirDZgv1X9ueivNJVOCwabfIr0OciuFnmXFsJe4LW8yyks5BJw+pnVqyyacBejpqihEq04vtIS
aq7Sv3JsLWDKqKZk63TdPUbIShWNQ0ca6+8VeNEThuN9Ly5ECuC1wN6nLFxsn7sQ+xLxJTE3me7l
PS0PH+zIc4UAmjtuA8gNGOy5YFL5v7c9Z219sRVfSnHl/nuaihf1uhbDmcf6jOp09fa1mX4qgeKk
T2djpTCx8gX0iZBv6tBXmFTsGjTcp0dXBChtk94xVEfcZIhdDbmu4d5Buo62PH8AwbppxmmsbaPl
BaviVY6YNpVPSQKgkj5eggkFYIRO8TEG9M9Q4im9tb8igHjPOGH8Be6q2sr2jkAH6/gnNL+w9nVh
e7q96BshJzGAYDJeStbJUiPQhv9GYY5FT4JzzQAp10nu0BK9Uq/uslXJN6kys30htrw2UgpXjZj9
cFMcOh8XwRkAMn+xHlgrhUn0uqhxUQ2+nXxJBPKXiagYVr9ofk/MPSDdaNgWValX+cskJJDfGIs/
hGc0fEow1L/qqgMwkOJ4cyt9zbFVmrFHLZzmbbv0uYrztCDnLH24vbKtk2WI4prOaTttUP2k2nhG
MfOqyMCCrb7uZ9AZt+Vq8Kx3J6/vTIB+m8eTQI+2OOTn4Cl6XzOrwyY7W7GG89nm9g+khuCA2SG/
1KtMdIec06/J9a9xX4o2gsbRjAnmflXVPcG8wI4r536EgyLxZY1rzph4g0fmBcNfJ7dSuC+0eXvZ
oZPC6FF1waXMXSRo11UdEwe9hKV9pb7HYfRSHeHIxpewkNEbZIygn/edsX4NxsVexQAfy60Ct+4K
GTjvfHqxOE50YFJfmCTYxQ5ADs393x4XUMkRPLIOEt8aZClVJ6ffwvJThkLHVAsytMYxQFrW99AE
3qx7A0HivYykMX32GpPi9wGkYskj1qNd4rQeUbD825XgwdsQyDZpHqrdNjfyQO1NrLzdYbdLH9lQ
Ghj9yTX3fi5kKvjwverG8g2sdR4+XpVf42T76Rdbcb9GZW2CsGyKWSqxF6iS3J+5HgqcNXtMYwJD
T+3Mo/UN59B5o3ez2EWDqBRzVH5Qawlzrq0aGfrFT9PF6+5lZ4p6CYIjX3DUvJCWTrOZ/DnwS7YK
nZsRQztfoHy2jtp7tNVcYxAKHNc0RKHIPIgF/lrLUshiQguIx6EIYAeSSZnF/ZxbybBq8tvpCIxY
jV86OLjECjlJ4/vTppty/MTBhRpxsy5AV0GLlfeJfrIrczQCSp0e2wIN+745uEAmDHa3RLI8n8ED
SYK1dH66OyNT+dDYIJP699HVY3qkIAJFV307jf3Ks+lFmX4qYDL+/7lV/yQpJ8mo4PqhCaSwBbnT
qiGrhEEB9Oi0Xn9smvHb9tZ30kyo20BYzJfTJ7VEJXTXbxqC1TBSqHZz6gt80E/MeZNrxkFY3T2O
iw6VypvvClod/3FuSk11NANf2umy4BmgIx9vOk0XkBQwlFrO0ZctDHQ5anfJ4BGh1KEGvCSLyGJ+
IN7+0Atg6IaO+eDL5h6HLsX79Xo972oQC1Ges06fwrh+ohmebnrFUBU0tM2FqtO2hBWXV+TwjLRj
GWrgaPQErJq4HowBkXwlWNA9lys6x3Yt9kmLkZi+R+ApqLxm126d8otrEECXGhnbTuKOoTqTzfCH
4oKFdAiDUcpGFq5ea5XU9m69x+b/syxFzvtB4WpjT38yZbXoShZJI/L71Jbv3jtX0J+jlrqvqIbB
dDJ24byMuBrfs9p+iOOnGHpdmyll5nqI399m1qaU0FDhvNvxhadlp4S/U6XqEBm4y8nHYlEo9VGO
4yxpRIdo8vDdPnuBdY6tsdpuguTa0erz9chXhLXXxcdHRsYam90j47q4BfTZ5CZyG6x3xSdwKRJ4
5dGbAgW/fNhqQ5ZYAI9DMf0pxeCAeJhLDtUitNETG7YifQxyYtBq0f76m6+iF15XQMX/DF5kLRkK
EgCzFeT6v8d5YUED8eH2oDDdNSu9lWkWukrMDy/rcf8KlofxQ2ici5BLWWKW5uKfW0d4q08xtw/7
AaJ/5qy33DCu9JwNhFGWAeb2D+kz3AzQnR4QvEWKgTTo0XmJ8g5sVQg9ZatmTE5UcLOF+AlcpRgM
/49q+tki/WC0kJCkeipdXPHlQ8s/RX7UYkK1PNELVq8ficBiQ9II4+SLsgA3rPd5CRrxYLFMxXr1
NLZ2LJtoOlJXS5mTx/FXsHmeT0PUXds3FPcLKMw1zbT6UeaS47OxoPtx89fTqeljHc/wqObDOV7O
+BNDD+Dfkw0tHUlOAVPk+2E2wSFSnVDxDID4fJRaG5HSJYk++IQXYqjlOcF/0Z98LIdqi6i8ce46
rZEw+mxQCB91FuCdKzTnLprmo7y+nbCR+ix1TnmiWdxiU+4a9b2P8QBLvnJfBJ4k54V6Pgt1UymH
cGhvqLvBttlcmpIzgsam+DmTK58g3BW+XrX9W3dV5tY3QJxmLnazClorLmKBWESPW7hOwarojPRL
QaQx3bbl5KUyFmfFvVXMUmLdVy3JZAcD2uskxilxPKl2DJdoGKeQALyQ98yv+OBSxDE6Oxd3hW1x
QmAYVkkqmHOx2UpU3rk1Bts/UZ9EnQSO7eNIvkY7uuXvO/XChuqfRM0z/MEf4bWA/Ix518peeabI
/A0lHh+2rCo+yxAVEdNQKlY9yJNBlASbnjBj2mhYZL+jl0FqgqAzbLPoUx24hsPioKuRJXTXlKTM
n1ne0WxPpVsDwUz5sJiaoC6aTATdZs1rcPbLFCCm8Z78/rKCsrRAWhaI2Q2o+0Uaxu7O2wBVyRgk
2+oX7hWVfuXoMEepi4/AhBzVY4ydlKC3LPxvzw8GuFjdkbuZgd4ZlE5NyYLOP8QD0lgugPVhenIm
h/NRppB2PM4WojQ1XbT/FI6c0YboiXR5cgMBdNX9bv5vtMBXkX0KVY/BelmBkNinQ0AKKNiKfwzV
NQFvun9r8PIrr/gnAKc8QbKbAIt+PoX7DfSGKu1+ml1DmrwwkSPZLwRMoZvUbJjnasmWUmNCNURq
s8bym8vfepPQpLanX7RtFAHtHn0yf71iCgb7kFtl4WUfNgWhqljrW4aetTWUsAdCaKAnujfdubeB
F1+WoHTYwRnypd58DayrHOiz6+XzG4GjozEXAmHr7sT9JO2E3cM1umL7vFyGgPF46lKo2ms9VFU7
5QuwGQqKRrzz+fUl0FBYp04oz7j8FLUR9uQTfMcYdnA9+x3sFBDcVOOkp7TT83VL6bFoKN5AiaWU
47W+G+6mwkf4Z87XxV6xfeiO/CwlBHFeIPqXGtAEg4aEo4Svgs2q1KbU6Zkte8ZVbGb6tWnEzCCj
qSjmTBMcYTc3sdyPQ1ZaeMBJucEFX0MT2B+/RpjDwaTK3qixGsL0QKpVRyIBt+j86y35zeTOAzYB
0Sb0FTzjrYMQyg2JPa6ShhQLrA5TQmH7cPQC1x+DYwZ8r0CWo4ZH604rwxFKeEX9V6XcwEbNeJ22
XLhcPs7SmLfEEhEtTZe7ZG90Zr4z0umd9qWP7gOS7db2A6xU6ejcg9bo9hIjZgdpuvL0xhrUxjo0
2wgVte62EJWY1mntaGHKJHZyDBktxP04O14Q8xxia06LXU1IYx9gMYZZjWl6veMwVF3mFQAi+aGu
iP/vBxRNhQ1IHrJIwhIZhS8HrUdHpuJhGjgphrDYeWSP8ZfhuiQi11kTQxnpzTLsBGDjZPIGBXOr
uFDiacuEVe9QI4soW+uEGUxCHUAIeIocFMULasNeTZT+/BU9IQp6yI0eZwg/IPW4Up+Aj0/pcjQ3
MtKA/Q3Zv2+/HOIPEoAoX0aCYQtcH79tsoT16EmsO0rMpTbGGxkxwlICp9bx2lnUZGQ0lhT+Xne9
lE3UuvMl3/TbToUYAEo9bK8B6N5UYks1jfjFzsoBzn0elmuxgvSq4RCRJVoXsRKOUMrbIVVgKZ/Y
HLdVbfIse1QCpKbswq/W4rEcDoD4vxeJukrVeeZzrFcV9C0AbWaOju1s31046k46nPeX4RzcSe0O
4uYle4/NSgof0nqg4cCE4rg7pYwvB2NpUJDLrA0kI9030L8WUWhAbsT48aVeygrnW8ApLqB0mfNb
EVy1IVKafeMhUEcWlpjBMqp22VKz7UI5UprGt8wnLhRCHKxexrjh76x8GZoBHVrZclTu9bmxMsTt
C8/QN+SOozsTNGwFZsBRAhXxgl6DXZ7cINjtyBwqOHwdEFGO8cpqrbY32LCe8vVGzvOAJ8Ue86kg
UT+n7j8XH7CRdW9zGnELM9KQNSHZA4vRVLlEUl9GQ+Y2Co1oa399eNW8X6Z67Y5xaTQdHsuCoL+r
cnKWOFe6Ag18pCXvdx5GKZe2l/nSDNx5R91rQCZ7+awVH4TRKCjbyBVGgJKYpSz3BV9+19sbQsAl
1oyrfpebUB3IoDrJipUlYwfjR0CJ4h0nCQLjhL5SmKzhiE1QmdxqpV+iFtMiKdv2yen+mPDOCRjJ
vxrMbkKq3xRWpPxwGujU8ZBHFWeYu3TqXMKVjcpP7G1WNH+LagOtmrkQGMdFNia7t56iULd9QcZI
xRDuRfwln4mvDoxVdJiQfxUAmV61hWLxX+4EyYaY7xHFtwHd/MPQWigmedlmb72FCPtuHZleDb/R
kOUMure1YSeMuVKm86cnk5N+RODhxF4h8exOTWSdX6RsG2M47WaJlZrbS/13aLW6D8hN2T3WPYrf
gIhshJv/w4bIFmTIzI0ZDzYvMnBIR4YQqfLuzOp8VtezL1hhLm0xUXTGZ5FxlmjFftVI+tn8yOzK
jZy1fGx+YEvIolMCkL3K760144ffnOY8nnNWGRg1qaPuC591vPcReBN9IVwmx8eaTbu5m8E913zP
4nYoTQFfY4Z+CuIDiUjff/VXauIh0b/o59t9rN2cmckLWIxmZLT2Lcpxnkd9vlH3I//v7pOJuYpw
Ro8QRp8fhvFrC+AdJLfNif8XcbAJ9ZPwWCPau5/tfA9+lV6DfyNM/JogvfQUGlhTxKEcYVtPFSFq
WiUwbjfBrAGG+HEbKV8mX9qHqD340xYg/eL8wQCtDv5JSoFe3WtA9oCql6H/AW3dcDjYx59tSN8H
8lMum8ioYJk0OSGm5+uogAJhqQEuENkWL1BU6qHweNJjuRVKFyB2kx7VJg3+CCIaVrD/aAgpfjey
8ekwrIHfm29g1OzigYYg7Woab29gO+L20+z0wXv/QASFZZJRTV/y59aqyDmHSSfdSuetIMtLL8Ah
fFWindhSVstRSybH9OeM+AfyHZbOEu97dwsZ+pAtvgHTNjMzc5kMK7HV2jd538mCIk2jzM4tOyTO
LYKyhSTxKrIvaCTLxIx9pEmQHKnbsSppMT9U/02NIZnxOx0GunZ/gSRDpkb2qlxSsED5SABkP7L2
2FqaS6qMWkMT+ckfsH36s/3oOSKwZGuDjKTp2ZoVTntqI4DxiNFmZQWnTG18visOPll6Es0z/ffu
5+JysH5NLIjftmuz4525ao4aAA6OvZeqEEGMhN9QKIlEf4M7ro3KaAD7QnSvWS+kPvEOGHbpOpsP
45ros3Rq8Hwr88lcXJVKxokK2xivqxzmIeZ2DiBL8crkhNUp2hoCmk1zVpEpRxonrvfTqlh9pvbQ
lwb1tvhetSC6dhch7/BhDTNqaC61UAcX06kqTbPAiEXUp67X2HmQrfouMPpsv1JW6PnPB0gb9Wfa
4ZyeI84cY7Y+8YdaF43h8w1fXQvVqnQS5Kurg+PbV/zylxKDq1v2kLjXPyCr92eTS8nvr11j3Nho
yiEPkrX0udjnJdYV1DtQnksaa+07xwUGMsPhr7KjXWwG6BkdeWCJjgrIIeNGTx4BksW/QjuHtpE0
3XqOAFILYGkXIY48xx8peedeRw9oXBQzHo5gewtWQKyg0UBoO/FSJ6UYTZIjJk9qc8T5P8lbzev5
1KHrx2r/s0luqeGiaYjFgvZBcNONfArG1OEoKUa69f3rHLuiRyPKOd//g1oDdjQktW12PPXT4W/L
S+KwEk1qSFY/AxokHGbIUVyuDzrtmuFClxPip4WdKA58ZAwRnBlWIHKSyQWyDOWFcIs841f5nxTA
DOy3X1FW6Xu69c2C/E7Yz8NzQIeo325b97K/ZBBBLicL0yGQh05BllIQTcrN+eIZ44yc/eEWW0dX
V2K2MOfozp3R8O4y0Fc+gVXQdEJg5aKoHIo648eiOPEHWVAXmDNUO+m0ASmG8fBK4WST9P9bnyxa
M+GaNoF2n7xOmAR0hhwUT4+NEvmTwhtvr1eETIlyEAAJ+Ktc2F2V8SE7iKeKLuaFUYyDyeKLKjUp
JBfv5xjtM3JKE5xqR5UjaDvQDXXvGTtKP3ESBY2pDr30VdzenH5vxfDfCLRB85l5ZQ0eo3N4Eupr
ETG7dadeWBblIAj1EBhx2HPMceaCSegNS15ImPO8rnJRvwZkiVTtgaKovEtlwBzzu9s2s0l0AL/b
aggg7WCGnXRclML+os/vdg7eKuU0M6QTxAPqBTwP9bbEI93xNi32HGITZBK7S8syTRjQ1P9z+hAj
EscGcycHtg28kHgdIdzGOfLH7qhLlaO/czkfQTYnDzitsDyCQIGC/HGbmZvSpbHk9CnzwvhrOzvj
gOMPX7C0CN85MSc6S68tOVnpLdDOxAsI7QWPvPEkph8a5XZBtcxDAi7/OYt6WdIcyp00fD1Dsq6k
Xzic9EUJ7mofXltptSOHPGE0ruL+geMz2UjoU/nIZKNomnaF5vSwlBB9v8qYgSJuoXWWvwo58Nbb
6fwxHdFzSBhbhub1hHRj1wbOiYFVHJGd9voZH6P+692IKuGYBf7Li1aaOSP59fBYLBq+hSK6Iou7
1X17ML8FgbrYbr95QVvG3UAWprEMVB6uCPygTLi0yk+THgbgMglO+sGzpSNaGVUxGRAPaG4sNsF2
9TmZNt+/Vp6JeNQd3qtxQVNYdrDDrAf8IjhNwIgmLcm/pv6jFv5bJKJqSElb1pe6vcJqHHZj2AbK
8IWMZs77ESqiliOaPJ+ni28sr4a3RCaQ6WyDWLy2PbnInLggH+E+k5uqN2ik+xXKiErzzlUFgPg2
YLl7r6UEARLaUt5RCXv3yUF0Anl7kwk7QL95tgZljlGkOUEKsoEekDyHItp+IpX9HC3CObZyjWcS
qZq/00zt2yDk57FS7BSE8Y7tmjSMc/ZGY0YsYfGs4CmeFDDIMHXD4ZXIGygbZ9JNBmmWUhvRKzzh
S8HMAdzNYRCrPYyjg9JqIRSwDabPLeW4EWBzwIj0ogHBMrhsN5ZMBsQpJNmklBYiqKjYyo3O3tGM
yQZ869HPIuSFJBWacBlsAp1DNlxC6yqTRnexwZaJtJIhHg+cXDMCNL62ANTt/4smzCM61cmiKhOu
EOh0suxJ6Pq8s5q7C//I5RhR5QBbW/tI5xpvfN7nWzelYQXUFNWJL8/KGwBVrJi6yAkwoyJa3+41
EZGLpOOFl/O2iuWokJKFlaYeSpJ2ybntgVQchySEnndx5hMywQj2zBrFcPVr1vAdRgkza1/YTFLw
WbnurV4JTYaWjm3VgqsEVc5JbEX3JHbOfnU6Sg00XEWZ3Y4fYOdMp/kq7HkX6VUNHhcOM1UlHLAZ
vvEyC9CDn4fHJxtMs8/DIN48/uSyjrqXeyCJ7/ei4tEEu/jOqEkwi5XIefZhi1zV+BWYMDGUobO6
M8S5l6tCV1+fBDVXk58oQ31+hnEik3oU8/qC8U7kkVkXyBphHl/4zoWTH5/mPb7XooR+HhO1m1ss
0AsAa9A/WYix/upuOD2xxpBypUuRlsp3n4M8ClnJE1Ya53clD8SP+EXX1FLPm1Mz6RWvN0bf00/l
/blVQuBt/Ow3Fdh3FZYx3AhnHwlIwgLZv/IOZqw5wnPo4DihVJ1pHlPWCATlNr8xyUi/2N/mzOrc
bvC7QuQ9aX+tp7NtXm4J7wOj92I7nCpcKXUnQenyR8stJ3KzTZSyqY0IMPKFras29xNxeAE8avK0
8rwy533bNXIGMsksCGkR5j+X/sRVB70B9Dsr5PLOJNjJk0fJG8WxwOp+D5EgA1jYOLO3XcTfUK+V
67jVEKbtlGbvJq5xMZVScvCiF3+QsmjPBgBFl6drVgN4rc0ZtQX2rFyBDmPUiClR+T2+yHgngqD/
P7Q4F7H83tkdunDtssQJNIRDEWQG4ymNT+dXnDJQItRNOT90OnjDxvsBsSflMKu5aHmtxPbKnCWh
bXl57YEmuwkdj9BPtUyZ43tys/swST2dHVnlaWsuwOvrRgfUHkgiCMg4t048sR8v1SJIXJk6bwo/
kKutQGoTFN90APb4wayjTFKkMS47jpFJk2264jxcBMDITZLdluorfJlXoOYD8dkc3D/xGkFi/4CK
Qqs8pLs2xott97gm2DdzcqpGIz85Rj1PvZnMzJvS6hzva7lvPMWqLf+lJZ2XFuWKJtsIQwn1Mt8W
5coClgiRPThAh3d5xIk0ex3AMEHRxlmbvn0MLXH0U04ORKsQI+zq4M1saBMB+Y1Eg9ba1ERvJqf/
WGd9gtzVSjHu3OhpUS2HBVSYMhwbfbTu/kTQ3lyrwDZ87UL8OpMfv2nayiVHmyleNsGi1CD4jaWD
00C/c9rLuTKZdglNNACyGhn2Skwhe56HJNwiAkm2L7umHNyNdaPReqHK4yonysLbOmS7F8WJcElM
Sh1liT4oTYP4cPwlKNcemAJKtbSTIXuFtAAT4SDl/mlbkGyRTP1rFnlE0JztLfHKiXy1T0RgzEQQ
NyeVRc+tGQi9z/KmKOiwFjjU32omrCG0rorQQcRq3IFdMnpe4l5NgXKy+2UZ1Oa1O/N709uJs1rr
M517zLj9XW/0R8tllNbx1NRBbId7/eRvz+vVCjJ21p1mn+q6N1Mk8JQRgoncD6nHLp4CKcRxjUFw
kHxAZb3CvsHXn1SCmgp4R2tKbtIaK0/XMWxZvcJGWZHHoz++jU1jpjW4Q1dSsfOCYx6BllclFZAy
RAJn/HtZvC8dtU2dOh3sQGXF1A118MYuCZvkZNFAGdBFdJfPhub/QKHQFKFU9SZoP4vhKdvQx7As
CiIX9grO+rXtWIsOrSE82JjPxB/j1VeZSJhOjRPh5zqlhp6wBhvqgwApCzKCUehX8W8yD9EmBSha
ZASfLToOLSEVUVj4wvVBmaIBjs0by159Iw6DbTC1v5r3E8Ag88/z8oIuPCPfM06OqTZ/BCHgDKh8
szHjq3Ysk2mIrU2zSscgmRzAZ5K8TUVt/PsYJzj2BiMEBJd7nGzSE3jwOWdh1NIpoPhRGkuR4obC
rxsJa+EPJmrZVzy9JRGi+6YMlMsNqZyW3Ein1f1jfugOVIY3F9yUEkOnEERl1tTtsv0JIHXiMA/H
05qC9oIMWKYU5LFZE+VEKXYM/8t6lhaR3jJb42MY9ciNeLIV0n3n42mmDbAz9+Q6W63cwYEdhEf4
Omnh3wt3niMK7YhdpAT8UlmNID/ZpEY5FazH5osL96aMl/nJCDsuD3yue2v2xav6DSK69hL/wj0Y
706HLc8lkG5IcRxyggyOmTSotOxsSWgw9bkKIMMERq9gyXQyuSK1uv9fEutNjNac2lCGVBArK6z/
g+J1DRQaV3T5plZzOLOpjAPsNIP4e+GX5nNbLnz3fcGwkZT7rV7eiEgWxGU8cqHD5JsM1jt5ZoFv
iOE/lUD5A5ILIzN98UzgPq4LvgbmOitZE5C4UIc+R9Z7Ej7zzLazOLmG0CPg8PLDxC3qr+Odl6nt
Yw07yhWKuB5H0D5LG588wBDs2WDi1w9XTBi3rws1Y4fPNJZNLR/1L8jHTIkIQXctcjFTRAG9LTBr
dSLc/6w1KA7X+qBlRMqcTE34lpqhJYllWzLBDqY5hGUcmjB8uZk5GGMs7rIfeH1U/yfcfCq9Dj5g
8ztgs28Y+3mAVKuLhxhTvw6oTj5BBNWp4Ga3VEnnFhxFeRjGhSp7wMBSSPv+0JHN6tu5CmQdg1e5
0FJn3syRdnHH6vco6nw3/fP0DS9mVXIvyfPj+ximRNjlp0V6AKYKZvHR8H+5CdDwfLaDO/34k0tU
2BKINFkR8s6nJEILBuLAabByAGcTSlJMMwX316dwXroyMPTGOfXDiYxILTO93/gcvmRm+9T+DJFI
1hzEN6Gg/R0lQPMaQQsiKfxl07lgTZ0WE1G8gIYiCldZjJKv+AlEfgQj1vNW6/PLKhcE/Cs1O9RZ
NvEHdkMW9eppTJZjoFxotnZK/OwitSmmVjGvwiJyGlvSu3nTrEHpbhGDMNlqsJ4EacqFwHEKkGsi
7nwzP3ZxtTcBnSrAZFxq8X2UHaijF9kJ/L/96vT8uvhhgl1JIvln6H6GWGj8fB+JI9rkoA/1suGY
Z0x2NsLlI2pBpMyVA2J7AaKLvbJzNE77hjrvuQLaMX1TflmMbzcmabSp7IMcBx6LlsViZQdaoZSt
OvHltrdIXlgWbwlKM/xrESqwMcahyclzdNxMWLV/NSrkHESJ1oOCXyH5qn83In6jjNC7oY8OynET
ldYZce7nfVtIScZ8cpM3kjzW5EVSjWJ2jQDdaipLcNZhP2JbfxDs7uxJKukgbOEtPD2zOqVZj0ig
CaQdbmXr9QpL//bkBXOxVycHfNdtFsSfbZNqgYssZiCQzkFCYauR+ECCyN0gM97VhtYq2g5wrKtV
ZFK5I4nqdS5gSJvtIXosYZAdNJDtpUAoPvLhJxQAPrMCLcnScXz5/kCLwoCSN3C6o+/Q0zbOF57u
ab1ot/RtB4Ln7S56PA4fz/uUnrhN+pH1M/OzqNyO3H95qcg6wu7BoYIOI8EYFoymG2TeNg2lxVSU
nnk/GG6H9LJDZ5YUJ08gWFlRa1vfDFvL0innjMOyeDCGJC8q4coptYf0qciP3hX+EyE0aVirIZ/i
jRDo8MUWR/X/5cg/MdJ2ecmfRS6ZPOHjhrprWhE4cPJx7cCfW3pYZ0E5ozzl9fECpMO7AA/4p1OS
u2Lq8Jj0h+cC+lxcuEmXvpQs52X4UKcrtwhaabbSHbSFSe4TdN3w775v58+JmivlE2bfRRZDoIbc
LENwzywk0FIL9Z8K2Sp4kUCn6Qi1UEvfOEJx/qji+dSAbkosE26Ived++a8RWoXBO1/6i5cE6TBa
xGo4RtyzIh7pvS8dIyrbXFIP/ugo/Exf6wb8CkVsEtp//3fpnq7Qxwq+X4jJpB3gGiMYLR5Z5T5y
baekLUiDPztL7BSwDJ539hwxAvvITNvaUQ9VTsujsG03SoriAQ9y3A0whUf67BPTUEXdr4vH23iN
zNx8obbcfPK77ob8mA8chT2jn+uhufb3A0Lv1gUb2vZVdzuiQS9zAC2iOhBDGji4IeuM8cLUItBM
WZF7FyH+R0Vw/oQF7UTPIRCx2h09heVrbuqurO1J/znZoUYfVhMrnIekrIt8M54JeHPY0lM26XjU
kgMpmIFf7JeN3zKHJ4RxZFOjf+ukhypWWLjv/K4tBUv2BtbcdbqZhhaUmkddXnyoZWaaVcrKGbbd
W0j/yGG7HEt5xlipKR+cV6M0SZPaKSw7+Zx/WnFkzeXQjCAWMq6edvKeSD9T+mVePdlGrTDF2Cwq
IHY+ELMl0bYY+FubGF+2sZYimHlLkflP/GtZecwEXNx9SEGpV8npFx9RwP5Vxrkomyg8EMOR+ZDf
1znx0JJdpNwrOjiWnIYONrgfEONL2t6IO0xwgkKVaP2uBjloVo9qoGMp7KZxcUS+DdyFZvH7P7HP
Gb5c+IKLLywskpUMRTc7tYV6aI4s7Gplw6ynnK8Pu6CcZTUtJK6vS/gBvAERYjEvdxL+umtoTpxH
Udi7QGJ36UiRBTJqIfoqqg59z6HVJn/7G7CcTHgiM/4i94L8TO/AHppWgcpNAQX5oliATz/7pfEo
U9tnIaF6760x06pBWfHz1rb+nbzQQ8YrETXOqST3lfcs9SUneAlci18/3/HloasmB1ugw0r9Ih9c
N73dEejdwbIkb+4W8avwUY8AuV+Spp9qjkpxbv33fOuFoC7FBa/X1WZ9wdzri/1CX512uDdw6aiJ
7Gw4MB5Ots7kSZtO5ybq08QJXV6H+bAiptlcGYPXp5xAYal0TK6i7iLfy71ULeiK4F7hz9qB/sJU
48JI1wr+ZLv5tX9GZ8eFde27NvlTLEIhOkDXXE0oGbTeyYbsx7dOGH2LxJ7RN5hZyXi+gGSxlh0w
qsrb5zRj/tPiJist8/uXmloPwyc/0g9k+VWXDlJs+UgLwpu1YKt56xpXHtWRiJXzqVA5yrO1kKFw
O/8Xfx5WJYRku1frP0WaA1kD49Zn3izEz+cK93o6mEeZ/ZEXsLGjBvid5N32FH0QU3Qgg3JZRjlT
3nHlmKwSbsHSe9PoGP7ROsgKr/jGYUh1/OfX8TVGoXjY10EzsuSVQww2BEOxvwgPC4hx0juAigJ3
QXlMfu0UdHBx9OfAsmkUbOVEYoyjPgwiQQQt7EwVtQSXOolE6w39LhRnwiEfCRzfxvFkqI+h03Xp
M9G+vwJlGD2P/Rx1+SHmqX8Cq6oILArYqDSYcqPCOMaTleGD4PHtfvLXRIkPTvseHlw6pKeXpF/U
Sc95xmZizzQiBAup026nwd11JeZ3CmS/VK7zFRbFbLlTpNoWP7hbQi/KkYUU7/DIKpuwuByJzXZ+
wY/g/xNdearahiIqjIMRIasY0lD4pr+TSTXjyGEdjn/ZObf/KsxqxwtvSOXTktkVNHVtuhUJ4MzL
4DFSpUMHI9UwrPMHC86sRzAzLkLRmmvhZaEG10FF7oViAy4p/p1XwAgAn+ZlY3Lm4ygFxo+rUK2y
GY1sRDiwyZ0+vBugOjFE18HzEJeX7IJl54CPK04TWvgUuFIe8V3lgoNZDsk3smCAUsomZiQs659q
sGiJsR0eqq3u+7haxl+gASEMvfusUuSmR29YdXHhbYeCcvI/errudi3GvSYT5RkfrsQzpSMaQ1YH
SLN+5H13OQ0Res2ijBbq989DCJzOlIYE4A/Mlegp7rtUR2JLOTI8oEqqSXVEuj4ozEh3uqLKas3N
Vk7qRO2WOJ51+wXovSM6Vua7dOSFNWjGx6YgySA2EwU4iXlSLjxPu7UIrW06AgUb0EgpcbzG5wLo
WisMeJi/P36vtJcv4a1HHD/K7DLMcq7PR9VhinheEJnEuE8MPW8S/E/q5f6uWhN3icu14z8BDqO4
ef4O7sV1cPvQPCs2vMtiDF9Msy/xcn/q0j+lBICSaYcMpQ4k0zIDUAE+8YKAB4LGgOUls6BYKrSr
oGfXQHZU+lJdGutyhMJHAbww1lrn1/lMq1BAORthxsQ4tYcdA4BhtW48DH3ig9Bg/fSVkcVqSpmz
OSS4LBrkMYcCf9bgEHZ7C54RGClJM2W28aDpQGEy3HJ5zCtbkN6OOV+6e0SmYsrKzkZ01OBXLjle
kiRM8daLo80nonvDM9Wj+eHm93/HPJi1HEE7EFUWhhSQA0FwAcOEbKV40UhhgQAgYfkuEgpmHmQY
NRM6c7X2tSTL01AOzT/lr7eb3mbYDnm91TokdQ+/vuC0LvDZAPVaDX9vbTsmPsdRs8kuS/3aU7+/
MxrRzDTKLfvxsAAHGdoFhuJekeV8/up/vEcrRT7t/iRuFDXEI9lzcjPdHKGkGrN9puWFXfmBnXFL
V8e/N8Smr5rnKxs2CtX4YpVyLY/fS3VNJEG5t6WekfeHxLw8Xr+t2fDVnFGIVqmfDTiDBvmKryMW
4oxX5UalmMSJIZLUduAZPfTxPsarsRkas1SRW9OmNjU9Dea91e1fITIRV6qHif1IyXD+eph+y+Wc
6Fggsl9H1NLGQS2sA8DMMi5bYe90CcrmNqXmM5lFxqoWa8CNvMojOtG6bu5d8LEhD1SxQZv33kjY
7ieDZTYoXdV10VtFgIbiFVeLU/D7l1rqa+2dyZd+NThJ+bdDUxtbBUlcyKBDWrF918MCg7Y7ChbI
29rbbPO3yTFFRX2sRW7mx61iAuQp6s26GU9cYslZ2K1oooGPr+bPHrBAf7Eg/9YQbBqy7s2iU0JI
HG61EuRSvKMlhbCGyEhcAQeuZQgiITfP+19UOVWF8FRccLTiFM4JH9Cq49NmU8uRMYP7aOAspIzC
mPcRTVZMXosnA/lOUro/bRc2rSEQ0LBQCElrbuavBCKtQPH+ZsMsYNoxfvngpnAg63tzDBuAw7fP
Amra+RELF1SRqnYTXFQwcNUWEwivU5JEtViEig3LmMxIHzE6ID9OObFrcHrfp9Z0r12UD9eFGoNK
PEoJDopTC+JWspjpqAsesIWxUOMBHVK2GW7Qu+j01qS6E1HpNOGw3sKE8lULrTW2eIJUDau6MMn0
hCgUVlS5AyTOSQWRlAy+huvnnzaTGgQaMPKBMNui6W87t/+mJIMLnJ6IsDIqAPx8bBIdAvQYq9Pt
YqMCLcxx3jl1+s9QXZkhdi5hy5PLIQWhaXGmWeHb7I4WKqOyAi4rfBE0LylzMEh4249TUHXRJwVi
yccvE7BaVkZ54bkg3zcnxREoA54AN8Ft6eSQsxojGhTQcTzqPWnRjRJahKZhcuZrt2XA32PTucaq
dP5eiuTD6IpUmmXHET4RpGlxmFi7hJ3o/5yjCf+LBjhbHqBmF4dlESuiAycHvZV4+XCOOp3Yfi2D
BDqYludcCVF8y2bPDYvy5nFBHv0KC28ByXcfvLLzfIVCMfMDA3Lxk+YsJcCIvHq4bpkccUMyEI/I
bGBnvBNJnAN7FHUmSQtIew44cUy+8nro/e58qO26KqBHRlJbm6nvqLL/bBCK/D8zeOQggwCN39ij
f/8kLrzEoznkuuMHyM98jJPgeeMhEKeZIM5oKcIVNHD4eLo3DV1wwNaPF3ecMgbW2vtQ8w62GKXN
zj6v+J1JjsbA0FTSkLLqH/khwvp46wRj8Y59jf8hGIrNMpFw7o+P58WkZnBxHKU/hinD97XsMRBI
korqvYh4PeE1GJGIItK8AE4fEsFJOeKTHX1dnwtocTz2vUyJ2PlQ1tF10I5wBnvf0bQr6J6s4di9
IWiCRUTVaywzyDOX0qzgHis/EJPyVFtjf066nyXtlXtvVAEWf6cd2Big3vUBc8ld1dZfl2NzW5+e
JNbzDqEOvJ0RwsXDKwijEFqbSORQDyrLNS+WFWEpCrLGW7bWm87ACUVdzN1ZJUJFrf0D9qGqJrQC
us56w6Ex+eQVfZu1N4AokT3BuZDeN1PiEL7Ee6BKWNfmgbWZGBFtlO12W/Rcsm9D6K3xDEDExG7+
70wGNXfqysfMaLpMYFbho2hMmKa+WJv4L84/rdQy9W7Omcyffuf5c6zI3a0Hnr0FTlVKMAvWOndJ
YZBT8yqDdqY6kJO8Y5deh+GHhAT1TWGAj12BDedXMATZMPv72tdGP+JanEl9dlp6G508LhPOrgZx
oOEUYo2mjbqAxHUMVmHCTd0ZgvMwe+x2o1ctReI2Zyfc1fxleMP892ikHh5IO3/tOlHGN3WQFPJM
MnJ7gBw3rwIL8tyqXuFpaiE6FiQKicIEYLoutOLXKIT96ahkPp98HZ0HQL4PnNmxaoukf1lVyNS1
2AGD9br8f27bJG/8dwhxyMPA5RaX1PHU9mCdIHAv5NZwzMxFxjQZLjKbnvM9w4QE8D71THgjqv8G
l8iNjKWlWSPMyUgJ/NcNO19PV/fsrt7sdW4oLwVktmu+SNy2jbrspcyYEdfeDNnefawJrVk7t/m/
HsOGKo2lgJoT5qRUeShaeQSFoMS5EXYFJMDMMRA+IP/1yzMPlOfCEo42qVeS4YBCN29OIG6Fwq3s
rdts6FzS+3p/XsmYIvUPmsRu8rGwnWnd2xnS6+q4NG6UM5ijqhOjDR+o56XSJuYuySvEhv1HU2Vp
P19wqkqqzm+1Nlfya/780uAcklSHYxLtnjp+s58JfbSLVHmSZK6j2e0ybHF7UzDmStTBVYEai9wr
VXXZhWi7QZf2KAXupD5cVkJ+Tk4gy1Xuah6HslHjX5P8QpqFaGsH22nwgZw26Z3kznlLmeBx58Uz
VeD1TeeN+zuyponmbFxyX2i4DpLB/15oGqLXBD41YN4bsvIxgCsxplwIBTwA5R9l1cHv1HKzZRqr
PDb7kRAbYAK6h6mjvpC1k38s4U4CjLTBX+vafgA4EPCJgB2ZedSsh2pCs/KLwZn0H/w6sUmYxo2H
RYN3UnYEfKYxFcG5k8HS8+1/poZmZ5XzuVAk4p9gew0P93Z9faZcsnt4sWw0xR4Wvhv4C/B+ZToI
9Hrl+5VosXlaV0K64vff8DcDWBf8z/xDW7cT2cFfoXpvUuMNHGlff7tmM6L0sgX1ykGnf+HeOdJp
7SDxGj4KB9+sGHMSTcUgChvlZuXl3m1SAvWZp+6myVxz3dHD50EBYjy0HmS2Cv7NzvrqcQeuPMeb
Ne3ZuUjORde11Bkl4J1cRjePXZbJOLn7XT0Ctd+cC8yS5qr/uEg95yF4AFuP+LEVarxTb9e/U+BO
P84YmGFhzEVIqkbj1rNmSTcXoNVvt5ksnSCNAGwGSGDrHC/ylBgw3wYExyXg56S+tQcoL9EFHQQw
p5/LVUVQ40jAKfOc1woB1AECNQAVzJpUAYh7zT8rgtaMUhredJQch70hMu+jv9wbd8TbAhhApCUP
OsBfOTNQ2O3XyqU2xy5AMSfswVcdx4ej+amE7rXeA8nt5O9qREHgPcghPVAlnaOyoZk6yYe1v6S1
hu9rstitS3m+bHhjsZAVGXpzsuBTzqI6kw+HB+HSuCU99pZLsPariygxwZLL06PJ40RlOsmGx+uM
p20HXGvLvDharfk1ylLkXumDca67xXRVxXw7AxUHc6jcAl6uXbRcHd9cUKJ+y5EkG3XmIkv1Rryi
VhtXcJxBVr1oqLOXXuSjDr6DidZWxg/NzRMIGZv4MQ2XrJ8v8m6R/GujZ8WP9col9WLz3awybZA1
3NaNWtJghgW0QJEs9QtJ9zeBjQSFwbgkuv3HZSQ26qSA3EuXtPgb3NMj/PHgZZ8IL0RuRzxanhSS
5upfBEqyjaSNeewJQgniZm0LUtHVIAkqm2Z7mnl5iu7C7sTzXPWjXg5w6OdZ9t8Ck+B1inostzkm
qj9nXGcAxv3120z/nYR2tV+gZAq1Kzw+IDXIWJnR/6baH8jirLIsnUF4/aPIjuV+CqfXz6/kupBJ
IZWMAcxOfW9JfY5QfAYS9x0aKjMGGVNAToP3nIGuXUqlVXGP7ai9H75YQB4iBWHWH5W41rJ9zpsa
lLSpZMI4mMvRIPnOBjJvJYRbajUnOmMiaZtlIM0UXOm01yEZbNPQLj60sFWtiqlxLlp2ZMsv5nWY
yj052L1cr7oI1hUWMbGhtrLVuAYLZdYPT8T67q0AojFKa9/k0jxNqyPvQPRjKQmGvr/lvdLXq2rX
40M05AhzimwrIQz15L+Vvgl4WsBYFlBUvdRB0prMlwaQqc752dfPECjAWjzPNC+zd2+8zSaJdGjI
5o6g8YWF3x5KAg/qvRpa/KrKNHVyOrQPXhpMvS+5cdJCc6yYIUpVvraqipX2sI+WRCzpN2tmYbEK
FJgUzMzvdgqCpt0nQoAeDO8Vr/U3Lmv2E80CV44XevHFL/Tk6nu7sJz3bnCz09lY8eRv+BO/0m5q
cfCj5P/Yn9ZemTlh/mtSTA7ngcQ/DARqHiJ87YVt876qBB0aYh+3fc11ra5vMAM3r6m8XXVxbpOm
9uW6i+JeX9Nk6BZs6y/QE/h1FVPohN1PbysUUWmfyCvRDGE1hSSOnhfzrLpjNwbJeQHcla9NIQ/9
xmg/EYgxZ8OZE33tZd4seX7Vane1pq4ZSB3zOOHSwGE/jVss7CCOnen5Bx53K6MR8Z1BVIjHaZO0
sU0n9Wmikaf4uY7jE1nVI1Tu9JOz/Zrui69QN56YBtaxfY0voUog74Ri32x8cp9kX6QQtmupfzwj
th5+fEW43DGvOc71NTmVblup4FxusWPbQaC1pbQNOOOKEaBgb6m239HkOqiUv8ereuaywwcB1ZBM
+JxKpxQ0kOwg267TLXDk4EisrAYpoNQAIZyp8Iile41QrgPmWZndKxhtdCDU4N029Nk6YsIvPvgz
EvowH5lnOFM0ku4U9fDQbMYyi63jMjLz4xOgG1NeXHHSNalA2eCmvZG1c4D+RfitdZEHzYUQigkZ
zjRx6IeaXTWHbOjG2KHKUHls+zUNeVYBTSQmxtqFBcXQNRxXvf41FxDG+3iU0k6oV0Wa30z41FhR
G7fxmzT4SzfpaWVXvo7z0h/9mqbiqYFsiMgSBi0WFllkPCx0RnlgWyGYmcy6WNt5ZNlGeDXDJnhv
D2sJO0Pe1CMFoTAwqHyYiUvRbIsrsXqdB/7YiAVDE+XRP4RnJ0B9R61rDLw4a0wg+yTNoYLagxI4
nLimvJYlLsFehR1dYdLVr4G8/BauiivMJ7SZ9A5V0PGSvV6bUG+k/l/FT+CeR+aukR7c2k7KMSke
I1IqTQHzxT18//oZ/lz8nr4QZNA6AoFIfnhS3d0DBDd8IAW8b3QWp7zmpA4QUfKyyDmIBQ6uP7pE
tNmX2M+nzKwQdvxMy5FOEsoVAdWQ0LhZRj87BzB6hUaruf2klXazcqOLvWQ4CRiQcT0Sj6C41yr0
IcMG+dSIt/UZ3hirhXmeYsG3Flc3SyNBhVpWhnwemQzyfQMV1eLPC1a4kxKKUH9jupSDWq0G1U9n
K9XK8m5lB4oSBKTLCsKj9sv6l50hCz8UCWuhf6h0DSDPedPjY1y6ur3fA44Ux+jFZ5lUXhkDqIXX
daa21uMQGWPdMD2r8LzWJkR4O/nf8UaU0xqLa58Y3zSJ5sHCrw4H/j8qC3FdXRDQ4+UV25zqVF/9
43BYv3J4iKNdjuTCzIIYi5+UKny1wf8juXvtk6ZrJwDhO9W6lnyRiQhi1I4EIylwSKXd3LGq8M2+
wfRnFShoW5wG14LC6KVKg5HJNJrueXKci/Dde/JKGgEqrGLiGzw1VBbUucIIlnNdBEXVimASpCJT
CeLXvSxPZAgdHYMGCrpJP5UCQ1iX2Vh096wMBTRhNcQfnGHeZHTkuipQBrJJClrYE1GzBkjl4KwU
De6fHyvFFw06QiA/2TmohnvqzHFvk5ElnRxBPNSODoEwReh2ICeRM+j6ueeQpAU/tSke3qPU2xw0
8sJHVH2X26OHkZvmdgi3qqMNYWo2kkzJeQrAOCB5DJElhVK0zN7U2vP4S+Iddiwuzw1tzNnSrTsQ
6hKkMIHnJzUGzFG+ZRxEGWf+HXv7LjiT5ThntYkvISFE8+3F1RI2OETAGKyQXgUzAfKgN9aAKZAI
ci1FmiBjlElwH4gCaXELRKTiqxTCovxNeVafblbijz3z6DBZwGF5EG4xsRgrG6Gw2U5n6EikM9re
3fdoIcQwlrQQ43vM+4T5O7pL5WDGFByUqJvhqYCuOXE20pafw9cmya1kBUHR+2LYvkCeZrVVmoa/
AsmAFXTYvJAhlR41XmkLi1H3I1xNJO/LiOWW+FjjwyXQeU9Q7O5br6JZWsFlvrDX9sXhDzW4NrvN
jSyfLWGr3JZapZTx2HOwi8vqTIX/me6zrPoJicfgq4a9SSY8xxUQ8u/oftgJ85Xo6NdRvlGP0Z05
GY6F/iaiTo83isV6VcendCMf/L+aVG/91+1i89BuAKuvZQlNCBHPA5d8N1wszCygXXQ7x9yu3LGi
2hsWnrE+RGlOqNwENZ0eQ5pibq6HekkE7X3xbKCY4CUeQM6V8f5FAk3QkZMtPur0Jrt2c7DkC7zS
oRcBaeuKGjRV81f2Boa41Cx70loEMRNkQsBUk6NtEXE435+7RmyD8zS1eTiH0VoOHVsuNdecdj/z
5tV7sPY5Orvblv3wrcOC/cOK/NDSRYfYRE8ImuVlkyUl0RmjSVjGgdRJoDik++wBjn7Y8MkyWVUz
3y0t31qg5cTcExhjy7vyOR3A9PYAcSGka2Gg/NlAVWOcqSmZW5LgWv+VRzvZ7o+AaFXF4L5j+PGE
ri5tm1X/Z6xOYYosBgOxHLDZZP42r+qpA6hy6ps5UEWGy8KkR1ZgFSFzsgWYjOuJZY6qhRm1eekn
ktFgtXCPbV+JTTu25TfTGXR84oBdUuNWOO0XGYDogxSfO2X4AX8gpumQblR9mqDkD0Z7qXjbWbft
Qn9L89R3mbr2ehKV2KW4ZXcvRb9UC4ZOdA1msR22GMr+K55XYgEz3qUiWLZKKN6H0HC5zwXlaDNi
j8A+nPNkSDPaH8EK/Hbd5tHV0YO3ysKN9GDyILXViymKavfQrKOVSvoJgzvFj5VsBWNTerKKvnul
3LToYWSm4tcg0Aykl2iljMQLN4iImF6leKUopdo5Aivpqtf4JtYc5sROyDqiLlCyqAt731dACM6D
LrsMNIriLjxw81QWcxOAm3uEGnLlzNMT3QBh02uVloZL+qb9eAJC1BTztvBk17uHHHXv4dIfC9AH
pVGfMhZq5d/AoqbCq39xRlhnx0oU7DYwxeMtMRqb2VZrV6n0RmRQkkkRlvz7dGoPRY1tZcpTd6pr
dhLHrN0e8XaxAtIeARl79vMRx5QzFFxKV1HqpbLdIeY/6MGetVZprcZZ8q8ZBzSh+2mnbBqD2D2y
qHY6d+7w+0EgeHvQM4M7q0USfmE/8hulNsVhsG7CdizNIdTvz+Vm5s/Kd0Pyeeb+z+Ecc7gXyftu
6mL0TepfYeoqLkjqOGIafuELgrrkoGSoEDAFl7xjB8eIIc/fVwXOW4sWlPdcxUGOP8Ece/b+GDNM
x2oFWtNGAXHMNdFnZ7spiAeODBhqvwDCZNp5iDHNCfJBGJN6QZwgNEvWWLSjZLOeq/y0YPQeAp02
7LwzWJSHqY/l2p8YnEvccOdFlbmmjbR4EZ74iIFDVwqmrw8zI93litRzCtGx0Je3p04HNSlXNK9c
cVScplBHgKc6CDNQle+YrcIuQ65HlXeZd3YD6hT6yA/5FS8JES2XlxpU8bbNe9CRHhJY9624O8T6
EUfriFefds/Z2+70L4Lq6esj+J7Swh1LhEoNFhGu/h61Pfc9Iv4us9rNW6kGivo3TE1vsP0uBjfh
WOpZ0xnOYFnX0OoJFgdas/QaMJHlyZph2/RuPfeP4KBXLFV8kzsG1UJz+Os4oVhDUoNyDjqlrEpW
KkQRaC9CA1gOz3b7HlquFGZty835zOqp3tyPcsjUzgWnOa+sBCgrvKR0wc3iLHOKFDU2UwE4y+K+
6ML42p6m8O4DloqI55x/ciesAAFU5wi/k+VB6+12BQZK6XDy9tqsD53AXgPObMSFyhGOFOVBGDWl
DwBrQxnLkZ5L6ncgSaELJ6pCxjxxbFCBGaDtGBT7jgFiAAYe7LEVxDBCbc2oEXIbRjjc4lXpOm2g
jDNI8jT51lv0nF9V2wb4CD2cUcr8XXXytRv+9BgtK/vV9TjGWMztDlSTr7ujESSWd90Wmac0TA+l
ZVKshFYed936qD5W4IRc6Cvl7WN8ZPqLyKzM303XDeiYsC3mjwO6XQN0TG08OX4hOs5pUOqU/5jU
dczAH80S4od52H+pPJnY4ivYcQvID82dUYmzp8H02Iv/sl8d5fCk3HwZ0rWnrbhAb78ocXidL0rx
YTRz2CGcrdAcPmMVPdxdS2jACJInLbp8cMwOwG6ZM4jcKL/H/VTUOO9x9251N607288kd9VCOanx
wCGzpZMRUSN5PIatpTKh+97W5XzHdToNyiGiPYlRPaCd8JfBQPL4bKOWnqTF7bjvP9lJ1WGvAeZ0
tliXr5CPs2YHDKlG2AmVBrxvQgOHjQnrhKMb8LKR8/5lgpDBZe2MvfuXKilqB3i9hFOh2KmI0KtF
ZC21DvGvFisVDyDN8JksuCveCs1GeBuILooRupJpHHBgqp6GEgo0kVrsKYGMDrWcwUVkpF5ApJIo
BMBwnQ4wYm1rjzGwvViV7Vma3nTCCO+hL/TEHwsV3uOB0Nz4YAOKlNYExgZsjXZ5E2ya5limkzUu
f6OgIlUnrRU+WYmoYxjtOrBREhO3RUX6YsFQv+6YMX0m5Mz9Ffb4YChX49qwZBQWvKOcLfzFGMyR
LWpxyTfKQtKyUMXoaGBwfqE6YE0zjDj9pUqkPEbgv8YFrBF+rIgseBbsgzUduPFXqXv4nhynzeka
D9wKcv8f9I1PgtJy2/tDYBrkkGeJ3BUFw0+SYfXgEN0Ibk9Ysy+1bNJtQgRNQjfPSAlRHR3T+A8C
/1+kpc3A3OyWR7z+jnxcabPWXFJsacjGzIto+NRir82eFMz2w5jGKtiRDB+HpNU995iIemmY/7PX
YsMTsplO9WcLlF98CpqyNKNoHq/snSv36FjU8bmPeA45kP7XWOi7mWY9M/i9yig+Y7fRXLVyUGRv
W3EyVEKwQrLX8SWlyXJF1oFuoTMWicWVw9LrwcIpEUu6OjxkaisomO3fj144uZ3ac1HQBkSLa/gl
zo5exg65HSNG/thWK72VqbQiKx/Bj81+Fhx/cgmCZSGdRWQkdW/12v8yetSgHpMfp5IrEczy/Zku
tjSw3kqVzKUCMfTGSPHoc0sqaJGkhUJl3Xsllnh8cX6VOkPeKtMtLRnfuPOa8vm3tJupP6KfBllS
4Li/cmpwDYwvSQXFqT6x4C1r3KulBij4X3BZh9FPTFbzIAInUjCpDcwLHNVF/t/7BV4Am4V2w4cO
xly9lmz+jtI0QYhO29t/29/b0m4CwtcKU+kn+nWOEPN3BpXWpLkx/qKVcq1Hxv2keUjsDHrtIaUG
OTVh4xyYQtP6qR0yOvA7N7/YSdlgvPxNUB1wXP6BUoS/D/4Ue+pXp/pFkVSiktRci7iCq2GGOnLo
kzc7WAiGM8RxOek4ggvRrJD2XbTpsxpZ6w68O2+4tPuhv/dh31aOceA5EcUfwuTZpijnvvj4xcwj
4VxJPMNQ986TaNtHRlwOLqJ9ypV3/SEhpwz6q5vqAIcPsOAh+yKLPBfxCybI+6iE2V36x2TbhjVZ
u8Nzn4LvQlSn9iTs3+p2oag0CYffYzFlsF/32OF7yepDehczN5PTNwawd7FkD8oWZPsOQw6Eqj47
2STNJ5Ym6/e7SY7IAJafDazmJX2CMBAm6UKaPsEVm3FEjd+TNu68s7FGXuwfWfXMm7aUaczd2ax0
uSFJNwrhBL9iqUGvaVuYMi2rrmaZM1iiyG/QR5BYrfwBgB/hIzo8o6H5CJf1nM68BLdFYya9x460
/Stqnpgd8Tpi323dJzp/apvG4/rpScCwx0RQoHKQK9MTeDiI4UFnVItHIMr+67/WBQB6lbU20gCk
rCitysWPjtvJ7fC6o+BNARWXkyJQCknio8J0AgdAxD5/b+OHXi30PK9GiIdiSJ+yfjktGP0PuFVc
Po0e2HkjuVqHYRSq9oYVJ3NA+rxIrtiV0DPRxQnTZbylcbfxSngHTANCqTDPBBpL5uiVnJnJFYMf
nz6c/Twq25zOp1gUZw1CGYGsk+wIusltcshMG44Bxdd4KL3onV6ped1r4a092RMfTa23YnKelvXY
E2QjhJcmAJrG7crMTFj656wmryiLZTwz0VM1YwrzezH29++WPY12BzZjKjHiTXIZAgjxke4ePSHF
gvwpmYWN0rGJL6PXNqDAvxvdHcnU+OXaX5C23xz4GoCyeAEPuySXHn7YN8ivYj1pIhJjHfIsecQT
0+bSkfSm7aMzwFQ30qTJOaDK2YhOQtn4FDY0rlBkUl4XsEto1Y+cVwFmpF29S0dKEnAitGUfyYTo
Oh4WY8FSsFPBwYaihPiNi1xYEbcAFK69sTfuyvp+TxxjyYI08pFNVS3tg0UWmAMTfCo66WQoOvkP
bmyAPFTEfhI+Rjc3cYcV92oUC9jORsPzewm2criP7jySOBbvI5HYwUlvuKItp2TBCz3pc4NOrWyV
uakdfE6UnScLehu54DQq/ZdLgUadQRff704+eQLjSgtvGstrauUAS9K423VRQJzC3Id14GyFrfUO
ORhzfFYJU/dz+TWUJSS4iZMk2p3+gQ2kb+uUjhRYbyiTzOk0SE3CmndSeBsjXh2ls+5YpbYqj6Cj
jSR1IBvOqCQv9fjCI10QVeIn3m6yeRMEqrMJGXghPMx9eso7FLT4OjAUaGz4kRBT5WLnkZIII8Ll
VGeCDN7XbqkcyO8t2Q9oWOH17W227CDMtnh1d/x6CRMHFDN7xNi0WY6aptblYsgDYyHt1Ip1CiKS
p0jdxnmYkKCAqnxcd46B5EX9wClxV4CnPMLYQtTNg2F5IWCby3hn/dd+OBhdnVMWs2xcx+wgXlsA
y2J2mV/DrLUxI0wLfzhAxupWYQGGWx+ifqwqItZ2NJKFsbfAqA2jWPjXhFvK17scUai63hb6Tms/
Gddh0AcBQJBBrDrIPODwfJo3NAwC/YeQdW5oGEDFKXHpHz4MN4QRumhppGA/eKIpA6BqfkJYsKYc
NcOYyF46nogphFlDzNqDKQDZekzqHADn23RvVKaN1wvzViwqKAT7AtgHkO7XI2OcT2O7gKS5UBO3
mZOQHTm37D+I44QXjXuDg/dlpO2pRAgBufKAsXn3U08nZoD+AFI1SYELWa32QEKqIlieP/XW/dx1
T5kPXxda7f6bxSHSSRqDjvzQqekbjWb0ItrisLvhe478lOFESNgs//dso+IMHk5rUIiOLQ0zMWUy
SRVjZyOfM9zdqKHcT20Pn/3hVivYFH+4CMJ9k/Y5eQTt7jwp3PJDfTsU2usb20y7VJwmLwIoZwpG
4dNtiyy0038JpwXvloQoF4GlIzmHVNo7hEty+LrY4Fdpco/41+tKEYgNsVl1oIfgn/uiqILAuKaj
SV4fffcVXF7nKg9gpXY8H6GBzLWTscRaIkCKwlaS5EP3DNfTG1qOdX7aMfX5hSX1g0gdWyBqo+Ly
IaiGdea0yDiDdUM+Hsalo0Y90OnWoIaM9nuFA0I0reZ0n/sN8PyR7bM7dymWmBbn5UGauWfIesJ0
lMr6X8xL0qoySeLkeceustJbZZGSLBJdVLb9qyuuXeaEODj9PXFv9jAU5lRrbMcvIt/VlCceQLge
MaxoT5qM0/qm1o9fhefuXI9rcmN29p8d8DgCDHBJGNBHKAYC4vHv0qq1Y3cUcUDtuubLAtBKIWup
qjGmMHeUtYzGMOlHvdynMTaj+Ht1cCqImF/+xTqVh9b4gCS1EavOFzop90oI14qTwHtq2JDH9n9u
nu7I/8loIoiIL1tncezDVwztg22A5aaPVG7JdhRE4FStDn92eWZPdMQgVAlqcGBYJbSNR9/fGSc7
wUqTGp6uxfFuDBWnreVYCfRqskj5SobwdtDHhlWdvfNoLAKOs4IGjXIMoDDLjrWoDkuAC7502R/v
XZt2ORHdh8Ff5focdNJZ+4mZQST4FSIVu1zJdtRd5FL2sUPfksfQdkQFfD0aKc8wQ8Xg69ciNVpz
iN57SN4an7WPCh06JkLNzQiWjinq+OtT0Ibh1WaplxLccH37X8t+u2oSTpP06WZ3/CU9GDsTmKYX
//kYkOTVKbKQCQV1v+ErMgoDoNK8bBJAN4au+pvng2RrNsKINqkxwQiYfgUQXWqkeWyOn7FbTpOQ
fSIDgdg5w6HU+nWXgBlzaqc3eB+GLj0Ld99MSt7eaECmwPmiqIVQjr/hYORSb99o70MUhvo5EeSc
cUrVi14W/WWMfpxsxMxLOPoKHntQSkNw8GjotG4R+q3SB70BCbTQiccuZU5IxayQ3lSjtdZ963Zt
lT7ckzLUeesEc749Ybg9pRr8hi9VMmbUX/U0bFxOLABIeY6LEjzNyRxS6NtmjTuTGzVhLN+Et/VT
wub1l4b6JlTv1xWhyx2Qle6HHfH2aNaDTLyoqZfF2b3yF2uxxLs0FkQAXc/RmLMNRqkBpRdszqAE
WIaahaXIgMpvUSpejlPb5YE3xdyoLKMmveELmWSHdEFjzPdgWNBQxHDAaIVVrLrI6dNVAg+KKsLQ
vcrNJa/z/ZH2z/LANGI+wmysNmIChPP+0yljctFwm4/iMFrzPhVe7i4+vA2OW7SJBdzNhA4m6pfw
5CFLVRZ/m5r2bpzVr22VfB37sNDgaC7IzQxUBtwoZsABB1UYNjRfYCnwmeOjiHC8dSifDrZIRH2H
6gCIpvqPpHBinjrXloMtJ9qXGUomtWhlQRqVVZjEq5xxV/Z9JH66/J46GZ6ueRWd468vXqMOp0uZ
nlAIL8+YXcUoYXal1LJd1lJJD+phbKJgwvfNv0i3hJ7Er2GkBK3Isi/CNFgvVS3lEqXLZOYoalY9
KvAXZ9OXFsoQt/prOuP+QAK7KDqp7XAFNZX3pun64hE7GKyyZgV346QbiV9+aJnxkzd4y3tbGy4B
uQIZv5PletwTjDEMZhne/wCk+Vex2OQaXIwkyanVKQusnlJ8/DHs+AzHCbXndSyjNRcQU9/4nhZ4
losuaXNUTnrIkWbILnXU1sav3WrXhjd+ZxzPfVicY1odn6p818TridVfMagONa0Jx2IVQfhjuJ9G
2BDyJJMtF1WHTKWcmEOuY8XpUMAr0jcmFxbqByrgeCGjisgVWdRwnBstc/RDZMlpzjIO1il1FJGG
nFTYpnZrbnDE5i0V41DfLOuTg7FrljdP0biKNfTcpIGCY5K12oPwY2I9XbBt5zM6t0DT9/gbQMGH
TRx+NVT1Lzph7xEcO1k9eKKZ8hxL2On1HM95ajg3odpB381cdhoisTxVJDTASBI0Tjb+tsBynE1W
T4+nmbmMxviw5ivBHuj0Eluo2Qx5Rb6ILD0TNI/cNdnCKGY12KhYCi+SvMLit4PCsQYRcBMe6we2
J4g9KJCt6MIf89dFkmiHWSN/ggEeW38ownTnAWAGuH39Z7GtsJB2XRVa81Ar9eeWF5Ftyur8p/13
T2fi0Tsa6+4DzjzfDXogEL43NPURXnBmwXMqWd+pUwjRArgZdcrAJ3j8AmoDtzl7ztlKN0In9lmH
8XvFPQ3tEeIyU8IDblo1T3czwtEm8Vw1JzVL0U1gRrk/uFJi2ZP+MYpwcc25DSlIGzjoWtk6HZo+
DwglVVZ5jp/Z9Ib4Vo7o3TXT220cOpIvBVkhr5pcpnx8qELaaLB5+g9n5oLlCFqITttgEgxGS6dx
IcfAozmWhA6kisqofMXtYawnuEfDdrEj6cAv/m6II/b1USGk1dc48LCfoAnA5WkW/r33G3Pbc14N
L2Jo5vbMwIIUNABfhOQlSOkBZboiOlyeNm5pKof03YP2jMccqPGKb/Y4CWkPkwZps1c31cqpkCvR
CmJfoiEQ1J5cQN6EWneIx4m3Bt3T3Pe4wUlU9X3H9Il3JvpghLZQEvJxCanoTNis2PNSxzD6XNih
LYAo90oJ/t6qhRhe0Ll6yXuIchzgoO8WaCx1+LpqRdNa1uasUuHZpOIDG9QEfN/J0k24PxZWBNu9
zhIp9AAQXVQnup+Ygd0VaGzCOLlug7hT2VylK6UBoohJZfFz0AJlpdgvsoQNaAXpv48qgaeZ5DlJ
a11G55sFcXz0b+KervzqRZnCDmAHkqLB54E1K/jmtGqS4I8xJSYH8ZeSqSK8oQAJ+fc/cieOyRcx
fudXbJbr7r19J/boUCKyAKuRt/48Npzsn4EZvfB1Q4fMf9MJlpJHukjDPKSzV9xOkcCF8uuTOQe2
SCNofNwXeDEmWzhSIgjQEqgfWIvTBR9GIToSEEDyqJxWcmt83XUKtDBBOkYNfmVlWL4mSxN4TjLV
XtdwwFGi6tThavfTwf0IdjHYaEkV0g08UHbTdmvi9CbOmVMHGH75tgBKvx3T1l0aNm+SEzjR6gcO
rfCc31g1mz0EN8Enl5SKha9jeOPOmNe57fSQczeEwVS8jCRQfM1EuhZxfAPAVqYnckiqYZ+TAHJh
dwzhXgkM6Fde0lDPbmwI2cg9BsWmVqW1FoRItFVvVKm70J8uo92dahYUlrWeCotul37Up7EkAhgd
yuWAvtL1k8EtnT/UoQTHvNnIju9LzuADUF4on8+jfYw57quzCPx6XMu8BtRckk5YPoWyCdPUNFPg
NtmsKc7DmVSqY8zlJsZJzX09AwUVacjonDBc0N3n2pPIjLoOyWo4lS2fmHsrajOBUUCHjux6qBHP
6834h+bewkgSxHECT2lho+T8Lvz+S1MU5BsuasRQBb82/PJUjmNr91p4Hch6LqbZSkhCepc19IgH
Qk8guqwXzWCh6gJrhiS+14z0iuG+sRdGi25OkKz++C6qmZ+qS5N6tXXFDjVAC47FW1T3p55rzSf1
Frf+j9sgBMpQauJlmMsgzWCGZXjK2SotS/3VudseMV1eN0wpzgPATW4bxfuz5YcvvkCnAiRpWhwO
IQjdlflByhL//w1asLzAoMCZbcoX5CKzx8TUWI4z6wCbtyu5i6jZBgOf1+fWim02qQ5z1K9jplLq
ZCwll0UOCjMkhY+r2MFpSsfeku5vjPJxdQ75SneKG5Gh+PxftcGinwyM11QXnbsdDTwdxztvECVs
w86z/yxdQ2Q7yiXUUYDa/HY9s2b4i7agK4DKfZ5UHJpP4XM7S1X3q9lr//IkmAVfyo+fsbZGenSt
/7qTYwOhFjCT1YqxkxmKVVenFabAzpaOaE49z+LG3Kz6fQPnOPHGNONLFxJmkrpcg3jRf/YPFjQb
8LF5kDmn0cSX17pCRCyg8fUHFpQN3eCXvt0RJN9Ww2DQPYu/RRDsw9QzHbLE1emKuhHvl0BxQnUX
uKeJDoeVL/Ra/ASNnb48+mX4K4XKpxsE4weAZ8n7gW0wzlBdbZaLv/s0VzBTF4wXbeqxEeOj09tj
BYxKByCbIvAGzF67JZD/ZVy2klgD6ueYzprxg6t8UEuMzmfNOuRKfAWWT/1sXjR7UlV4NM4fQPgo
ZOpxbLFyPJ9JtEXwQc3vvaVNmiiikW9SwBS/7gQ+rVUwYQlDUpSCtMl2I8tNq3QVqzdoaBiBdJuK
j/OtosCvP1MOU+rarwE6aUv9S7tZ8ckboeXaZbRCvZ/pk7fKp1G1ZJTYRBiC5zcimdNBBloYT3W/
EIbEdCzaq2VxlvWvC18/2Tqvp0VNdACHIvdFp5owqvVvCViQlzP0wsNv4tBK/cAEQAzI/JiruXIm
xMos+OGIVNxGtugLH6hqwAaDpO7liRpgzls/ldMm4ioziSi8WkkGIjggDt1tCVjBc5fX/kTcegA8
/LWHG5swdWBI5gix+L08CumpxrpxcuCAo133SYdLxf/QcnAB5APnfye0+w3gWp3pY6xia4b57vbG
ecURrUC+T1/pQyISJ7X+dyz46VtjkMD3F8lmJId0uLS9Gf/PlNOdWIIXCAl6fpguLFfeBIbICs3S
33hNl9xjemtIeY9eOvgDGWoQq8UCdFzUO5+MEhVclTK8T1ln1O7UBI3aMcD9FqU3NUWoG+Ir8m00
HYV/KmZeuesuy3J285Tg+oBrew3iJqYY5ViSytkB/4N3e7tamUNsLROCuFla0TJK6M0KmPlKaFWd
UrapH5hFTmcwyk6eWmXdvXXR4XQgE5b0CiYaDy2G3oP4zivfiBG8NsLqjyI+cmm3ctfLchMCFCQ7
EcEnBahTGvVJLw64tsmKtktgSyET3SyPUZ5EL+sZglOiIRj+JUon9Z4XvfJVnjZQu1gfgCY11d3n
RsWj3vQ7xowzoW6brjZZxNUdsgfXzEj2G6+dPbzD4c7DDKYp0FNh5JkkL8NN3mAapRwuWLse6vET
3jKgl1veejjn9ajAY2wNOHKZOCZGiZ+mTK/TWKTQl76FG/tqxf8DnzZ+NFK77Rfb/H+TaN3fbrfo
9VL6y6uxZsoBvb2E0iX/ihCmTDYDXlqu2OavBfcjGbkkn1uAipcHDANc8NOSm6xkZDHbVwwfYGj+
AdAO4j3sSUKYlNIIs2vZDSji0bvZj3keWNqucK3Fly4PyYCnhqWrhVpZmMnL8xsT1Fii342zbLpc
PUDz1lyDGFvA5sdJYIUiyygStoXXWW0V0iEOe379/LAi7KCyqN3F1ZLHg7ziNweUlU+giSy41EKm
PwowQn51fHiV0Ung9cOQ7kXQvHklrW5xbLwfeCiGn1JJ3sOEcO5CTJs4gpV2DL5HhU2mG6PMJC/6
zzyiv5eSgPKRz8vc9/qrgZej+mslyWzLQaOxxT/V6C/yUM/MCIL7PHt8zD25+6gmRLS4MrSEAK8a
DqsuRZ+rKm1P1qVEmMJ9pqMJpwpMKMEX2gsBBda2PZVaH2MzgQ75hxMROUtY0U7t/QdebbLClhpQ
UX9zwXA6tAx/k/pa4et6wz/NHOhRx4URV9s/Qap/yiIwGY4jyJESO+4fxia+BpzA2Sbn3iN9irDt
5wxWUetksPrMyCEepOuSiFjaBWALG403zTm+fSQ5qEMVSpe7DRYlnQ6HBU8lxPWCh0qAcVbq/qJI
DBpotTw7/2EKNsbqp1wNSb3oK1rtXoETLP6WHJoojZEJQsg1dDSmadAwbiu/39YTAqvIVzThOGXz
hi29XiLbEwW6EgQcxnnvNPu5gG+zOsZnAH8aVDbEyuzZtFJHN/CgVdyBwvEkB80jmiWxrEowqzoR
1YjfyALFB0h422XcHPKMwRieX2KTEXGtCOYbyUI6OnF8ZfYMtNw18LxzafyZRwa0L1H5mT2acZTZ
6YgdENlVh3UWjxYvdWnMy3zcLd5pp/uYx33/+NOyRpxM+EOY4RH+fpMBMGcvPRYPUeNW90sQ7beg
zyyeQdHKUbiYz2QQQuCLqev73H9QuMp46zJNAXlMZnZ3MBl175uOm8j67QSx6ArsDCugK/S5rxWv
Gvtra9LKrEiZI2GeyBijldBRwoFP5zmZTMzcHunZEOQ6mcuVv5xemRskxzeg/Lw49AM20zF76zaI
/Za/lTacPz/hqT+WN4nmFN7ZU+b7pF6FljQdr8nVhUgeomdB98K3gufROvK7W9Hag6QzrL0MxBtp
/3Mq28gzq8DOuQ9x3Ov9LqbAdR2IZ7YMTtXlVbxB6L8E1nOh9ya7+NQzyxgXoeB6mpi72vgyR6M0
4YzZCDlfEXqKw6N3oxjikvE8rQgtNdwjmbK75s85PxalCbwR83EExyJfACtK+zyX3Z+FEo9adpmN
U9eE2mDVREsIQOZqSJrtx6eW/EDQDmxn+NXQo2mzEVDJWnV2/d+T9PA9TizYGo6ciWQ+DTM9r9O+
Pu7lyfeew05h3kTSHjapl600UOR4NhlPrhrBzsOM6Mr8JLKCOvd/j1MXv+Eai2so4d/gMFaFH6/R
5VaAt5jerZ07O48avYk6YGIwklQkBq1C68u4FB81INgeLEmYrRxG6qD0MANJq+xCywhbWSC2KBzx
ZV+cHeE1iDeIi66xxrfkDAbr/ZaK4GdoTAVUWV4LNsEEK7KJKDpB5BJdGkmDrwHN+E1WbQJFB/ci
Q7NG91oAlgk2FMslflXcAST0GPCV5I5rNKJ0eZJ0W097xpve3/vSTZxp7Q61Or4QI+v0bRhGG61z
NErlKnYQt/BLLk4zne2zr2+RWGMSEK++9v7jk4xzqXRPJ0CrsYoNo9M2hr1J+4aEGQ3d4sLprZ8q
4Eyl3kSW46fVkqcguZuuCubVsAEhvzU+WZxDZBVoRradgjOVyhoAn3WfU1O7zKXBkR/t5A+uMoVw
d9JaYYl+luS1ngFFxLJfpaYlQL34NCFtRFiWWpviI1lYQzdXw9CzKkl4AgOEtGE1XaCeIxqTnu8S
85RO4ZJhOZ6WckhGNHPQJc1FoxvAOv3QyObqAxc9wo9aQWCVPSA+OVpwWZjVw/Xk2QKzI08fc+aP
Jsol8fPtLzBghAjI+cAVp+QU5cG+uCaQVa+TcknWNAy8hI+IXgRw3jLKYrFtjLsB9ShqRoo8mcaZ
WTZCJo5NyYQ6H6PRdRBVlK9gQG2IbjZIi4LVkN0UE1I33rcqqC5MC+P8crJbcmK/3x6WLVLb+fNS
KljkY6/NryPC6RAWOta7sPSHnbK3yo1n5l1nqi3LDm7fNbvgSOtMKWTNg8U1EUvpOyrQDeCDe3jY
GrgAVVNk9261G655pDrtdJ20t11ZyjjpamLMwjnIGr/d3dfjiNiXML3PVN17K7ohznIg11MM5YbY
K09Veps/TUKd2gB/iXrsAPXOYtbFYdelZvnSapyeQi/wV0VMATVJudyIMYcBkuBBgYxZ3w+9Zza/
0A0Dx8lwn2rZCUlwC+Z9yeFGdacxAS4T+SVesz7jFGazsjBJYASzTiGWzkdNSJVpkvgwl9qvZm1z
GwAo4ZQhDr0RlSbiYWX9pVpIG5ce4p2GQae3HgySepr1Y0GR4gvk9IBwM2RgfqMrI3YtHp4MfaFw
ctYB3FKd5B+wR/ZA91reUM0lmPCB2hz3+mgKTdoz++YTmBA71VKb5319sGo5pwL5zqEYXliKNYzW
TmOVL7qO3PuX+yWl7AG0vbT26WRLGfEkOUWBTFk8ftMeKTHOgoH7FPxTswVq0hvYDckvIoLqOOrS
B6P5GgSwghHgEQEYtEN70tHrasZwY0Iy+ZTMVc+/SAGe/h/6SE8ll3AwtJ8Xr8QXe78SJRzHcLNE
CwFh7dfeGPFMSFgdYGVqYAvqw9+nWKx+XJTJJHGwEUpvpuI8LZJW0l0vMU1O7VDZOfzIm1j+dSG9
OQ4SIPfd71iIYw/lnNtsHJFsZvkuIX8eukz4yxLvXxhvKfzt1gCfYQTZ8t5yZiSld3DkimcaBgy7
o/T5VB2CvSwf6++icwaMuwRJgoTt9bOXrF2ZqbYXTjiNLfWyDWKszA3OP01Cd5ZJSCZ+r8vUlEw0
WvHa7SaTz0gZYwyjPrNoDUlhJyMqPp1MW5cGWG9CqCWylOFcwxV2vxPFHx+LXjOjQCSdmqt5gCU0
J3w/7dwGelq/cLNFC+OjzitqvG0VUkzHCnQUypEZdpWOJMkks98BikmG7/aZl714Ao48HWNK9tw9
cYDY7Bivd/2WHjfH/7R9ZSoWmWt22Yi+t1UXwSur9huQg4t//tpwVYSZwkceR8Hqt5HL04g0WxiU
j3kS+abLjDE7xGY5XsI94jnaR+fZ60Q98e8d2U6b4Y2NlVZG+r7J5jeDrJv1Py7wswlPfgS/56J5
8gSX9XgGIAuRHFeo/FiIJf/dChhc7w54RsszfEnZiiPhYIqH+1PzVGgwBEkV5Qt6jz3TKY4WSqaX
LEy4d0j3na3sE+2hJgwuOG9+PM4CzlIiY5ziA/WF8laNOcGhhzTCkRY+pg5mQlBYOFVDnBKmColW
Kgol5M8Qsr8/brxjKxQ4LtqTX9ZSXsnv22Hz7q93Wuwz/U1XeOKhwzqtvkqsY5zxAdQf7rL2U1v4
SK5C7MHEFWzK5CPZVacsXf+78SJNAFTssrYAhpDpWM/FiOui8hmExr6Jt/0/NV11dfKn5KjjI/ga
Z9LF/uO3rIEcUiBDlNWBl+8avCPpAD2rx/mw41jjNx/qDh/SXwVOpf3h5xhmwZfbWPOMerOgzFcn
Bqg8nnbPgDz4Zvoqi6137v2H/djW8hdW+SLNL8U3raM873AJpjTfy1TgqAFExHDX1VGZlitz5D1o
moqd2yjPaYKOfJ6n3OmfxBk0Oli93fxC8fBZv5xxV+VRq3bulXaPg9nWUd1ghJcST/5VLeentI+y
SWGkdP0IprPRfVdVsUkk9OeZUBLhcDmBrvCOQiBMsAxF8oqF0jpeJHVZn//1MnESq90749BSLbLL
RXA5/mZnIuXwHOzUtDAY++Dyjz2umZWr7O7JfG7uYwCaihCnZhddvMYwKPwMMEtbpsK8ofsGWVd8
9nPz8YVq5duTGCyH4yZDe4nXGEwvQrFs81qKbBTiwvnBHt2TkdmIO/Cpo9JuDoZQzf6yY5QaCXWJ
YOcoqls+lEWqyE6z1LXsHR2VaI3d4z3SFvDtC0kr/zct7lL8dYm3F9lBjPAQqbv49q4dkmCRHc51
ythOj+z27OHZIRFWpkcwuRFnglbTtWH0vkan68MyKwMiV516TQHsxrtAF4Fhc8/Q8sLD+yirHqop
dCs8VPvC0nOw91QUtH6mANe+YIXWZBvBPCYnT5FvaxbeZZnS5dAHpj58re06KcwheEw4BA9FMfN6
VRg/BjU7uJHXPsPmHwzs14TJDne3AirvumHJlI/P4Ns58wmf6qp8F/j4QchlWVvKxvv0TYmVW4Xo
WwL/jmo+0l7ay2Z+Fhnid576SZqvYUJwbCCkBqeeBuQ9hsy6CnAyDZv26ElyeCiSLcm8ft/BL5z7
qQAWS82uLIJ5Vv4KF/uILMutT+44KQAysn06pdhEjNikDnqegXjUA4eRegfGonr39hHgFqRiO/Oy
tWPVZ17jwrg+FvYJ6jyGoSd7VG5a/P0WP/ajr8vzD94452Suyx0khbdCbFhAR3XjW64zKnDxE9Ri
2UzzJNV+eFntxcJypyBKdTKH0zIqnIWWi9bIfs72DhTCYO5nZXEPx2DV/FM7RXENBTvpITelBwzQ
4zmK3tbjnWtggo2fdiSvKsGrGotxjMJgyjOfosL3L8k0rVI9WhGtm3T86G4rzT2e43Dt82W469zy
8KaPAL7HJI8zVE3SwAdYlfDOiQpPxTHeqvzn9lDrsj9UYTkX3L+dpkwXRWqEq9UZKY5Za40t84X3
ctzIIbpp8Cqk3ue98edvYFtFXiZS7Zy9L23bJHTP1Cb4m+sIP1+AzT4gskjUq5AtRwXgXF399Eni
6Ey8jsxT+I0ZLernKik+9PP+PojU3aJlvfADfy044RIV7SDPSLqi4CLzQD6h0X6NWMdOGO8UqKra
YNDiFUaEukyZgVehCNA0ddYhQqOFYhB3CUJMda2JgB4OWhGFIwugk6UD2H6AqgO0QU+1cxV+OeyQ
UZUPkAg7H1eiG2tAbfPPJic7zgEZQT7ylxha3AEt+XGxwfX3GhPffWB1fO/Enaos5qJydO6Ptd03
i8ImOd+GRpVcYCKRMPODusUCRWBgYb9PPvyLpi8d+glOzsXgCAXfN8kOFxoEFRXj2Fr+4GImXBbr
x344I7WrCb9Fck9LHSTsc804MBwnrUe8I0uIll/KiU2lJoUiA3Xe/Jjprb9qYmXEUbe+e3Q5VgJL
hdxW2LIaD5ftX8gVapvB2rqMVRouUuOvZ4L4+O6zccGiCmBlGTFIlJ53wTNh+nK7s+yf3FkIjmZN
7d4KjYdCid/vNofq+hVnSK7c9kpaRsI3G8ganQn+ZJRnTkMIRf1oNK/jxzXtw52C1ak5A9mQn+JU
8nzw3pJCumORKSJR1NrhJ3F6Yl28IHAzO1IVccBHPRDTG5iPgKQw8dw5p4spINrsHvqzufCr5nRW
vziF6fcAlB+Uopu8z7eEvP9PpbRcvh5AMsDmH4CcJfO7rlyRsIrICRWFWmnZG1OOvye/slxSLUQo
LLa5bli32bWq5h4zp/lf6E+BVVKKcPrQMAKBGK0RNiFF0mUUXECKBln5z6RgiYfhq4ibX1yKT7rt
ZkR674b+D/ojjPomFw1cXjXVeD5a9JT0nzxstCxNZ3ivGe7mMkA2QK6JHyx1FllafTfdNTMQ6ti1
gIZzYEET7MnbPsGmPWOjy++UQFM+YPkPsUp3c7rluE8qB+yhxo0nmBT2eEPaY7LffZZvgO1dbH5K
Y2aY+qu3xu02XsHxvYsmSqzSKM9+W/KJyY5dJY2YqZF0dJRLrF12YrhsJeRHNwd7P5B4u4woUo/s
SS9aWwDWFzzfZTY1mEiXvdZJEJGt+bzWjDtXfl7EmFIQ9VpU0UpaQqFXNR2bFKmX/O3tReqF0lbU
3dr4lyP2UcJhRnxscF6NDDrBi3hWUc2fuCNWAgjBx01Blw8yPxBBtnMZRmaUR60siXQuVMeVrhE0
lFx1u/GReO0XmZ6M45p73WC0I2xMBi0prztoAP3J7KTHdphFNdKyYAmQ2uynDoX0X9GLO7IRRAlk
rboYuK+KTMLqYcodSU8f6uWnEK71jWNN6p0eqokVoLS78mKQVF1nusbX2IJ6iAECzBJLS/QPdS4m
xp83ZEKsc/hMH5RIWPnmdNWiop/j/IiYVYbXOnELZ5OvoRctF9igRx3rBSNsxwalRcKU3nWzogvP
nMer5qOiE5poJo67U4UpamRUQMcMvvgECyShjnhUGNl+5KQxbtrbcgM+SEfQwnXkz4CNb1cu1KGI
52B5iM0wV85k77NpwsBMqJpi1NtQmRMCo3UYHvHakxgglLxV6xoSJdbu8j/7q4SbvIUvpxUXyqZW
YNx52AoZha2Omva8wxk+v7044jqhGkh3wkp/3HU5nT7+qz7Bw2vey4vZSLc4WCu6cVr0n7Tca3Mo
V60N8ihyQltqEd34z8TaZcspbaBhODca2kPQyHhQzE+R4Lon4WWBudpysE/9vxtC3OONwlM4+Aq2
ODGs97x4BxCTO/8y5pKI7H34lZlmsM4lqSIpMPShpB/JRKUTrPcTDrng9UF6npv1yoSN8uWKBoN8
p/g9rpWY4coooMiklgLMSLEmL3fdNsIgY5Wk4kKQmes8UTS8JXuLjnP5bs9QCYbRe8UpQZRWgBtt
NjzpXHtOR5a/90ITMwaJIB6yHPSZ63vi7tbkwqWkYAasVVAXiGh6/oqaQeDyR0hwS9Fe+iUr1C+J
2+LanMOuA5JvcwAjbRKiKj77rPHpzVxUJ6t8EIx15hWs0JnONQHOSBqj7bkKRMc7kpJs1jpXIdRl
xfElmK4nuXaltOhp3H9wKrSUDlPHnoMQRu/wv63xlzqnzjt4Y5oRhGTcpX1ZsyIEdHm4TZ/k+imp
+WZSZw9Q/qnCXmwbJpKRKqbZiCH933FparzFRzTzy0cdS0Xk9Wike5eQ/FC0vgFp2HYhqdVrSeIw
G6a6nY1CGq8hfTHXL7JsIkj7wZzNDyLUFhd6z0HsPqkfC6KybqTQF1a6n1oEGuAlfGDrqRinDoA4
nKK9sDpDb6uAaAgXGs/kvPMc2PponRtGOdydQ6fHvKFiologupeLlF7R15bAHASWrDntE0lniFBa
Oaxl7Nnq1R2CmFusoMUXOa0VpvTC7Ax9Z+ubTSKhs2K66DW64Bl5Y6hYsum5flAHdeVKDbYYxPC0
0mYJ7fuyKNxgwqYnhUX2I+JojbvCviSHwPuIqq0am0FsBLOAZWVZuoMk/CXjfxf+LV/1iv9kvHJX
PRiwwvC9f4ruEMNE66Ss8SmtjPRYTxVTueKdQAyEs14Y/OTUAi0tZyEa+Bt6hwqcr1XDJ6l/yNNp
pBxBI5mO4Hfc5VJBzxY0Dadffd5AI/G7As8TdwVcNGxQrqPrx4VHU8ez/DTzpSVampOYy+2KJnz/
bxQxcoaPFAzNI5IlNj4VoBcgLId9YIyJ0zDRPeQ3TZl+5ER4Az0x1uAWatr2X/YsFm+ekYjhQ0BL
aQAotKb3ojpO6QFRsL5R85DqIDste3ptnC5tha5FiX33CmunLCzP4F23qxoIF6RD4ACzj9466Nf5
XRxI3w51Wvo0slS2Hf5FfVyVHv+03WanD27m5b0RGcSe+XHp+MX6tRKjvvB3nADMKz9tK0ZqfrQ1
3vX1KxRjQMAwjaGY7RtFcfVaA0HZPpOvHwrg8f5p6dQ6EbbXRXcA5Xh8zahKDO+dR42UyA7rw3lr
wRnEPrIw7/UkuXMSK3r0YV50jemdmsShSgSteHnpm8ktniVHIsiOUQFhm53PqAh215JCz7HA81CN
l7dcpAJ12UiSA/nff2mPgmiOW7ftp9Kw86q5qhOd7Km4Q6BMahZfm4hzuCLD9szHw/lMcj+F5rbl
lbnlPh/I0asEds81m2UZEhmwhV4XHmRoNEgjqkLiYrXa3p5/e8OL5ODxh66ECCTN2gHHqEaFfj+W
UUXdcIVCRb5UmFnmzX/3VT/Vcp/WOoBf4V/9lVomWdnBtP46/bdSRwG5/VmBHPqf/0wh+Y1TWaLl
4l13xUGKhls9FLvF+DAAqC0L57E9fPfOgqXQA9BGHBAgd8tgIvjtR2OjWjEsuQGXpR0s1ssXGZ36
q/fFrdDRD7vskPOANblGTP7TwMfnHo9rNgoOBRMcifnlzPQuxx6L8LmLVdFZWjVhqeMhtALmw9tf
IQNkxRa+2teOb7s69z4xdmgeQESKAkdMPkfbw3E4SkdOe82AzlZRhz0b1rAv5FuYwDOKjhH4jkMi
6ZKipH8aqB4Dz3lbY8FAj6kUDlVODDijonO4JIcVpacQXMJ3m4LwGqOiP4KENRO1zMcbclpvgeNx
K/VntIOjEyLE0roPJ4DnrYy9T1uhKjL7OgTObRXa+zgAY9lM0wuHE8AkVTarX/K4c6xW0q/VQKz+
btyZtH7Ps6w9kQAv3rp8HQUDfHbWuvrIkqiFY55mv9L96zu1ZmN4MOmVxLRgd6uHxTQNX6mn/0BQ
7Y/jqQ9dn2mtu82moYMVxsgvWgvUztZnCUi0I4YlvN9Apipb7+4Rne5k9BQmvyjpIU2Dd1Om7XS/
VPONNFpqI9V8wYmYv/OLwwRROc1Ex4lCayicqN9z65aEeeg3yDxPsbxz63ClsHSEeOAIPLlaI9ur
pzG3MxLehC+ZxsuGmz865KGzSk6He/9wXla+qEub3mDJ0CWYAnS70CDFDoSDL1la8rlBQF+l4lx4
ylmaig7imgOccnvLUkovPGz9srbEwOIh5Cn9faMdzJXVCcRbU2zHkD7M8QB2RkJ+zgeZMfhuvpHU
+pmZnu7SeYdA6bEr5Nus5syMnqLP2TlOY8Qht83vAE2Ha160NB9aY3DrdZBUGWsTY1787ZWr5L+x
59ZdKv9SIoTcFFcLgpHbC7ffGE3by0aVQekDWtthTWo9jZSmS5Y+pwri22lrmE+zXQWMN8bT+YGm
sUtqlulmVzwrmqBCQmyFTTwTg69M1jwuOYkmvmlo353FsX0KqXOKVYquu3KvLqbLdLKdzsHqei2v
jb8dpdSA0Pcxs5QWww/xuPNRjC/iNBfpBulKSIY7ie40Ly5pnHXVdbf26Hg3Yjf159lbhLHEnAvQ
KXnAxVE80E+gSbaX61LacyaO4EuNDXG+WBjqNg29SWD5Dsay5ykIRjwVStC0wb/NKj1kW8Rt+iZA
6O+MzO1UUeUrshnD2RODFfMF7flEnHmYMdEczPURMZ4qzpTOQEITopU5/7DiGTEqvpHkKAMdka+X
xsXiruXuaITHbbRjegwbZ1WEUED2u3bqbDlQDcoEO54mY7jOGpXU4V6yP0YuOWPJJRJSrb0ixmzy
BcEbLJLgBOge7FlwYA9KMc7r2HqMeRo0u5FL3a6CPB1XFlXYRE+6JGYnAUbA0GIQOIuGdNgRCcj5
bul4hXSdhlG+5LN4Lz+pyFum6kFAuHJ04taaiZDzgWi/AEsS+6TRg3KVkjxd1H1lJUN7O8bLcv8E
Uq6xHLqBE1X0o9rvv36qB3d28Fj5UjZIYjbzHxdQOOi8kCznDYVNSJOrb2n4gbj1iKLLupMfXoAb
TEWvQ1Kcz03yDEx3FfZ432J1uQp4Tke4NbNydm5Sf+9O5ETtRIjnquTpvdzN+cNZdBwEh4SDgw2E
HO+AnoUB3+0UJylCzBAK1NYAaMuv9aErHhUOHAhn1qGQ2kgEycVRuj/inp3QyeLokqdFxSnM25zD
HcudOsgt9EzD6t5CdiMpAvpnn274uy4DETVELGz1wYf7e3HF1ZZH1gnSbSWN9lofefhfqftfTyIb
cV7s7eGpUi6drkuFFO6hLHFd/B47lNBhRfx0n5g9m88Y5uOHM3tf5h3dxxBkWr5A/pcii7AUOi2T
SAl0rHMkO9QPMa8BnUP+4vWc/PEh+cxJ0Fuvdw9nY+8bt46scLt2IGGlNkiXCkXsCL538tUt42Oj
EtbaTVUj8yiUa2fAhqhRaOvRpMST0Lvf6q4dL1y/dV2gXM31MGmWS8H9WFT3PUcJkmmTSSyrZeaH
kU8C0bceGgOQ+KJWqIAIfQzVybTZ3Qydg8c4mKptx3lISZcKZt/T/AgyNd0KqvT2kItX9yebArvP
JC4IkgLtn1ZEtx7A5aI7buhK0wvezMcvu8FcQ7X8F3dLHuXUCZaW6qppsd7T4FRBVpme8ZTQC20O
XZGu6T0k1CP43y0TACtUT9abVlbzVnL2mtNYTA/IZOjcbhgU8rcx2puIWPXmIWjW4cvcWbtihT2w
dqp1Sm/s9l3gSxUGHq1q5ZzIpZF5mBi+G61WOYTfomnvNyypPr/G1UCeQDTWRhV3c4F2LVjXx7D0
FtViwJeih46VTb8BrZ/FXTjvGDMpE0URZK+fjrZ/rReD1gYTJ7rWzh+7tOV29eansmlBWdtaKbQx
jfaWTW7GAjqmdwrDPhUozP4CzElW1Gks3gvkbMIhtldutMvRwxYwOMZwBlGFgWPXyxsGrGKQ1ZxE
pmPRm1PTGiKv3RkxpB1jlLsjE9RlxI5E1kOsCnxx49mqBpfAuNYo4/ThvUdN7vE7To2wuYX9vj+M
RrBPoiQ1oD+sORiroRIUvestkTvSgKWihB/qDp4K5WNGtbZUZAHNNH7DlfQ5PTGQ9PmWz8o3rfwd
Kl0oLs6Nf1fsnhgrK7rr5ALpPrY76Rz7D/rNg4ygYbahhJNiwOg2wAM7CJ8SXH1P+69I3XxDV598
tuYli3e8SnQyH1Ze27gkYJlcxV0Pv5w5HVqjwkDMRP6eGh+w/3CitUYHQfByKxo6OIaZzI+MgvDt
OXt/8kS5C18rH+VqL7gtwLHvaY7LIhYyw9a/5cW4kLkvygE7MG7imKRjiMMSUQjez93sl0JZTK8S
6vWFUluuwLUuy2v5r2/1z428sCGt62bA38AwlamOOR8a/gHif6elm+WPAPH14/UloGqtDHDV8F6u
HuXcJ9FgWDLqcStjpoUJwOuali72y+GEj2uHO4nOtlxINREx86Q/B0oeIOAQhhLTt5gxGEoPUqlF
bktjrYhJS8LtZ+3NiEAOCjA3ljF0514osm8ZKswD0Enfo7wxgGV8+/P++0GiLAsnEVulV6jmSVXV
RlPa4JJzirOrQVIfRndMaE66b9O2AtT+uYeuZwT0rlxfUqRcyE30/QDngh9ActH1z2GE3ACX0CwM
rkN0EUHMWaNF9LkCqI1e28HZT7JArPo8tVAzSH9wCkGnHoWpw8aYD6+pEDbXd8I+Pi2mmu/sABUC
7McKG3yuD0E66X3Lpxy0l4/9LwTOP57l+0Y4ujXEkHTG7Zz8NRXiMMG48Wq7WKngDb2j2mtz7Pe5
0P2uGX8McLZ818FTiv3zdEw/NaAJlszCI0VRfTcnecmMOjKkPEef4b27wy2imAVSabWh0bkgMTIO
X0MsJt1odFUZhfHCJZMibpB2SN9AoZ1CK9AEXpYuagNVRas01JNxNftVDHTrg5KlGx6plTMFQ5SQ
KAY1u2i78JKWeXMgtRdvUgZPEiKOA5HFQCq7uaYg4feN/DSfKWxi3FzWbp1v0RiUrX8k7KSnEEac
SS77/Ops6rNIkZaqYuSNJDrkAibkGVGmhxdMuIIILbmm9o98dBSjmQ76ZjMrxSJ0CIJIQFZbdPcM
lHC7LdvQLOfb6ukWQY9Pi1qZtd0jQoqP73Vim52q9ib6tNp+k7EvCOXJtuud454+ljS7A0j3lTJD
vZGRL06kZUemN6pP+eofkLEm7rxuynFOTGkflk0JDPCqCh14OMJU3tISPG/fynObHWRBvl8prfgT
io+q06zWOg8rb6tD/ySngybM68C6YREmsEdLxxE5lJcfdxhs148P+mox399UShhosM2+ghfRnnmI
jkbjpaa16JSjy5kEBzwWMQacAwMTuMJYj2+XQMd2y4jz8ezy8BQJiMpENp6/a2gQmbbRHIvFu/UR
Gfl18XK2gtVtoOGkH48P/6+Fmgc27zw2jDZwy7X7UKn8CZ+IrwEL9e0sKvEseYRRJmJ9U5ACME70
gdvQUdsZ9mfZwFTPogl5lzkwHzJ5xnitWJTm9HkFMvP3KD+sVXvVdxsE1NfRMx6p0oN+xS7qAhDt
d67+ATnAFP6sJu36uq2ngYkaIEdkm1Rb0y11IZL5JplsP9hs+P2ReZ706EqbjaH6FRc+xI52mnJ6
aL/LEUl7jC/+mzYoptsbOYLdM1RxybV/Ll0pNpO2t5VCWetAR8X5E72hK8rtoEsMGwn4gNzXlffX
dpkF6k3uDv7mbb8CJMjd+vLKgOUmdHwW0oiSFBVSmapLAHceM+AQUKP5tVrfjNp2juqEZBzn/E6H
h6PpcgXxg69zyUsgU5AL2f9+hb4MQSN3KSSEVGoGT0R5civadzC5k5l+ArWGEHPPmABWN3753ZYC
UQSjRZ+piMbxChl67LgqYSsrSwhuXUz9Ym5Lb5fZwNubAf3IP5I3p6UePaeaXjP45djBH3MmIgnK
BiT6lC+mi1x8nxGnU22+hKhNHBjlEzsd4JT3xvNfKHznukPXxHS5ZcVDL1DBUW2tkjTydTYj106d
W7hXvCdI5zT8pujfwCxpaxkw0sFaU0F8G0l3S7SLiQVC/n8Df7hPmbN2Nt52WYnEsg+y0Mfx7xp+
93W12W7/lpMjU0CObi0tK7VrFdFL724DTzuM3wJUrMY+vCrOZaHTsjzMc2SnuNpTrFzbCFalFeU6
UsSZ/3SdodYQ/wTzPYe5hOF1eFM2ED0QWttB0MhOyuTd6zJ6mj6NcVwyu/FLmKQSCh8fuYdAyqhV
m/h/HDaakAF0/yl5urzpidn87dR6Kc3Z4uM4fXBsW2WjNYqEAyvnrSwqDwQqYYkb7uaGn3Zw1b1x
fA1mbbD9l+xI6r+cYWu/QAfu1JPzb+rxJ7wl6MxlYJ/LaHb2LJbSLlYfcMDbT5gCMz8ntSXBPZqH
3/O/cixsxe6KCju62DhxZL4gh7i8B92f1QlnjteYJXChrkpXYnGKQtv9X/WlFTTRto0UajD+2YPR
YrG3/72i5upG/RSdFmSRl5fcfaWD+DnOcnc6ItxuVUVTNa635XcdscXx7thkbtgs1iUdBGTLZf6f
8lSNA6+bbzRJuMb3gdsXK5y+eJSpcBKL0OfXnZzw56dctOJ7+L/8aY/4IrD/6rqU016JKItypKIz
GwIfhWxliT1sAOwIAgfB8U0l2XoHuYVvFUNVcAhDwPJcF+ft/04Ktcssn0UNKH2lJ540P1dfH+E2
tvsNNftmlT6CifkzTAz7xZ7mUbNKEO2c93mvMoyf8cWDhXMxVEwaRNE1vXoTExMrRpNwT8wJ24xE
8Em86YQeJYeg1Ys0pvEp+8q3eQC+ndWUKparbfD/Edrr5VTGUCCmU+UthakdvQaDLKqNRkWVsmz6
nCfOS0lway3EP/gQMNysmmNvdDHGb//F2oYx/aLWFdhu6nudUV5bPCm1eb9XB4MMXHvr9pU3be2E
IS0/jVxf6SBFIn0qzcF5OjEto4gDqG5aPXyfqdeRIx7BEUtyfwqdTNaQkxJsBNi/+/nN90UsDJsY
0ObaVhtqhRqcY28ZylNazLwsQ9ZoF/tVrQfI++SWrpVNdlOEJAGgcLW7oDLCeJcp4OimWCZluD/J
A0uLKHU2vcQ1BsaNngVi/9BykmDy1ehfYY8qqb7gB5+dng7yDpcfjbp1kS1Jes8olxSOPE66z3KZ
wCKsmPccdEoxVtAkPk8Er8eInzpRxJUz9x07Br3+9ROLnJVxfynxf0TrwR7k4NFghpZHJ940tNND
rngUtMx/o8LKGWPEtntmQIw7UtssYZ5shoTVv4XLymlKAwgOmCuM6zioID2kVWCv70Xcr605Kqjg
V5XBc0IC7MGEj+ae8lq2aNiN3lJUC4qXRdj7Lwt4S7tkU8Ws73MZU+4s5HaJjCr5B/DwN3TG8F5B
9dNciw9sLvSKtKTimnyT3F4DN0LO6qa8yN3vSTHm7AGpBF/0A9X9WpzPdcFQ6GtSH9BQE9Jhq5Ez
G7DStix9uR2b8Qdc5xk54QPEdWfzLAe2+z2E4bJI67R45Dpus+TXbXWHs8uyIzuAfkirkAyfmlUX
to+UGmQfaj3id8EK5g4xMfwNTCfgRdqH6g6tQF6aPtX/YGj9hPTWNyEXgsxox0zlkFrOEVcEhJ15
F7ryPK9dcWuzdh+7inp1TEZIJYaToEN8XzyEwF7758p7w+BhByktG8e8QNqh14zBE3jlCkXAnts9
RYDKXgYqm8sU4f8ZNI3hS3T4vDOFxqCdIcchz65qDYPDk2xsl3pmawCWZGiew3woibk2m7JQ9vcr
evGDaW1OPXYh6ihsHrWlqTczjHbSHuBbSyLfuB8YuPl8f5vS89Fk3X7yvWwRY3+pRSUhrdNk4rcz
yoknY40/q830dMBg0/3T7fTba1MkyLPlXo0nBhvs5NPZtbkHkzwFfTx2RZpH5AB/TLH/wmxuQm+S
Hm+mrX/68dXhkb27/c/fVY3b4I0CbGQIi9wHt/zvpxvdDsLlztzUurGouyg952amQfcx9IV61yZ2
SvxAMPzB68vhOefArrj02Hd9k8u0i6tuLRYsVodJqkECX4IsMnRNFugcLOhOEaqi/LqMRl1CbZuA
T90ZHSZKC+FurRw+Igp9Lt46jBZooCs+iHDIalTwbio3SvQ7871YP356IwaEtfDZQc0IYhptGNX4
WbSwtbhvak8YLnsP5yCdYNwqnrnpSD9CL3/DtA0x0AXJ7vc1H7W3MYEKE1trPdRN04ELzMPvlEFL
TDgelboVdHE3lRS9TL6cwbeNUYD0VzTlkBGALVI+TUN8eJCENwor38K/aMyIiwrvQKe1RtLml/Uz
TnPlCjgGbjuzQKuVZR3TYk2MO4XHgqkh/CUpeYlGpTFo6n+iHDguXACKIMcxZiGQ+2BnuXrSzwKj
nRfaWYZVHbm7E/5n70USWpqyyy7pQ4Nev/mJ25LsPc97tqbUHe7wiylJnQ3quY4qU9jnqCsx2nLw
n/9UaCiRubQt5d2phD/9HOmOPvOBxFsJN0Fq/whYN+bUNXxDvYWGXfMe50xuu6ZbtbBwRdFrCQjS
yhTK/JfpP1ja4WVonCE/mKsJ8XXzCzO3z55+/w4fDD7bPwKUkNZftg+a1JHCP/gOz3viKMGKKPf9
JqsIHyDarmY6KS9B1ZaL9M+MnhPfu/zqmEY64tjZCwwBf2A+CY4OTLz1cZgZ/vkO2UT1iiRHi1qt
Pq4M6yXj2f+qDXNjphxXZs+4Pfg0QrE8l79nj/tAJ8BC6nbzYyFkxVExlTN7y82XIERubJ/wnR4T
aV90q4C8K1Fc6VxK3EsXhIFxVaiERMUPtDv69GdYltxy2fwq3hNGCwvazPuOdRLqTX1Dy1Nf/xzn
JRWRp4o0gFg9kIERQKO/xab8LNeKujF+UGs/l05Oc5Z8abnF5NVeH7aBDEbFkj9f/t3Cv6o3FIMZ
vyAbvPmpOgoqRh8QoO+o5rvkCaR37aU8dbOE4p9TCHxMFt+HSmrhsBZKWexAmtBGZhXW2nXc6If7
KJmcyDTPHloioIwgatE5CI3eZXkytujU27pm9PA6U1qxml71L1+Y6aBD7EU3n0RzltIcvrMRQVFr
DftAeELwdBPKklrH9Yn0msgoCOqFg5kTz/J2DiiLzGkqetQECJz0YMgZBlC8OvkUzoZphgmS2cZ5
AkXJJxWmnMGezqMfCVnN//rO+/S2jn/XnJArWnUtdyQbdegD00RpMjmczLvqC38lAuPpF1K4t3Nl
0gP323bhj8aXN0lMJaKT0Ddhh2Nnyq2xkNYBG3Zq0q74pVmRDZglLG5iSakBwlmnta+4FU3TKFDJ
gh45aywDKRf3XVpfMAQaqMow4HQB5Rm6NTbpj/Rr72DhL0W1DzxLv0AP1qe+xCL016I3B38gCo8T
Ct37rtJ5D16K+BAtl8WDJua3xAn9H7MoKW+K3oQE1WPySY3tvXWvXb02C+Hdo+WDX+IPGVDdOiex
ZhTw9GOODYaeqndxW1m+JBSprJIAFX5OPILUA6pgTUTn5s3ZM3v/sPv2bm6hAFsACdfT0ZYybmaC
E8cIM01CimrLKwGsahg9AnSOTC8y1FHOxiXCaXDPjNsmob7j5g/lKydIB7SND+eFVTOGMcqf3LqF
fc8C4QfOklrW5F3feFeibuv6RJIYY4TrkjylmV7nH8RbDWQiMc1i7I1Va53lpYvmVQr8ztiItxYF
X5J4bDCBpuy0ArEYFadPw6VbemvNV9O9/DWqT9SVIXfuoJH3uieyMeJLKvsebwpee1EHOBmtTna9
fWpLHTku/Lw0RZKtTid+PYkTjTsnqO54PwO3x3dEZSdoK8SisigG/OxUZQVyyeDeyY5DJgck52Nx
lfVV+VEMlGPygdIpWVbyXgLmLhn7VS2Y2iq0SjcY3Q97k3XWmt8vPZya4JGoVkZJx4w9sYHtAa90
G/uF8ozne9G04b0HlsMX/DzOMYm3cjBErvGOubNhQUv6Z/eL+P9XG5x8JJCuvtbQyCe/HXouq5py
JgD0G1CtPja6C13nxzZyslrux9IGPkh5mzYqfSG1s1G3xqfyoe7Uqxqhr3zoIVtX60zpF7Z5W6ML
0aGMtliYIXc4W70rCkWUOoelGwU0GhCIGUQbV1ForS3OTG4CkRqBVX9yNYfPVlZEmvi3d2s6OPVH
zNgnC21pbJNKS8opNz4P762he+SbzIKMpqpRQH9GKNxsVmln+gEHZuUNy62HciGGmO2Kh9UyGRFt
E1ObIr90kyIvnkakb/U7vg6LhJe5VGWF631sfLHi3dqqIweIbbyzHjLCsdUDBWXt9c8pyrMn6+3x
B9jpJT4PrJzY/C8Kb+KoxbpZGH/5bzXmIJNK+oeXewo7Po/N+sBWk/T7FJoDHSEcVVCvn3vICeOI
dbGnGFu64Zu+mvbKmWGg5V3Bne+7O9QQpORaJXZ8ao7iI1wxyVdI32I725C6TUj5GGxqBdOjasC/
lP/VngdOV9BWHYISNmDork4JpJHmD8tfhROtsk2wRHX/LqzMDA8P8SsV0ttPIjy64feBGJjfPVD8
s7zpnksjOah3L5jEKkyHO8+k8IhSdi92/WhItY6F3jMd0wDYo4Nnln8SqFF0OaXYgqNGltJuCapo
f13tUvar0D3ndjYVrlMDxmMjsB1pvXUksRO4ljVaR2wmq2tOei36IYNBAoIfCn6hPtSCmj4a/E7O
1E7pTIbE5Em+/t3lqAUVWu786L4bOcofeY4jHrLEKG7TxdEZFpip2fteFApmtLZYzqdqgiOuZ/I7
zzkoX1O0zBQNGqX5tck8gvE8B6OszzKSX2ncGzLeQ3UyPh0gICk60L6tcG+jRiiasx8602Q89+i3
aJZD4TlpiFD0HtKyipd5pKnAWWI9nE3kBzJ0NtuCkUV26cp8J1VRoW1ePj6GygvI4Ay1h3HGniUk
1xixFmJnL6XKRSr2lI8dr+6hRtjSANQh5QSMci7ugayUqH1caAplB2NGo8nHR5z1PdgWYycSQNm0
Bpf0+Vr7CeLIYr/fDB2ckS6EV16CWHs62/2aAUqyGCEKjqcmKyEi5E9N9MlFF+/wEK1wSnxrirf6
dm344z0oW3lhI/tUTnX201G11sp1c0La5/dupqQXf6nDkITBYIeS7TC7oxyoM+4IUFRQntYuulov
oBMzrqNHJewaWyBbecyG6u9BqfyIIJFGPZZUZe4oQnk/eBqBLWL8f5/KY+3hMjYhTyS7e10QvHH/
SBrJ4pOcYcVUGMUMmC/nF0Iy7CAfkHLpqXox3A7f+CkDabb1MZ8E4nZ+geT5C/29nNmP9EUKpaeS
EbZSoT3+3SsXB5yWGjT+S6frFjnnndlwwnhFvWQquWwf6AmzX7hZWt4jmHGvIw63Fv1i6QoxJEqR
rHQ7tmvmQKQ/QG8DMHwxIvfH+aJjlgXO/WJ5uorM9y9OnznSay3BBKrPMa6xxabpTtCpy6zik9gD
+S99wcE0qM+JGjuQp1ndcwKVIiWW6/Sm/wdZt0vbQoW6zi6kseUCqFTgRvaLo7r+IH+5vnw3pJNf
hX36LLKM2Bk6P7aFzZJlF7MSPcs8kKWQz8KZBSeB14QMaYnFkuzZC0goUjCyxQluewrAC4RCVisK
vn1UDLuUobSofMnyBrQGYvNVLkMP1HzN3c/O17gYuxbs2U9pB5ZFi+c8aEinja/DKdwKZrXTchkl
KRi4cklSaLDZKLz9DUyUrUmcKVD7apXn+Sq3XlmvEx6MnZXrMi4mJjqjseJgC6nQVf/xewKAmWXe
2GErrvzJPrRvwQZBcV8ib9nZvMqh12mnRhP77f5MXAjRWVNEksNSZJUvcmY1QjVH/Vw8Y2TIWQqb
j+1LOtiixffQ0K6HYAG+97jjFVqx9wAQpuy3bzajL7l8B68QLjAp9GOziGtT3qTTrTvM6jg+KGA7
RQhUU8lWSKfEqt95vy66EbGmi8G95I2HkU0b+B+Mdmoc/94HY9aJ88X1oS8apnMzx0ucOzjkegvl
WdQNAMDIcsOVV9GCeqeHScm8UINkxkGMp98e8WAiRaiszITlZ2yeHXa5DyNWdqUMrRVlpxnbzmw4
ib7j5vznu5jhW3SmtxK768mMR2ejxKTIGcLs6T5zE4NX+4zX+U5IvFy/WwZOO3Qj2ybPj0Q3tU2j
cA+E5LK82DI/ELz886eKV4tkN6Y5BYuTxb3eQ4CFM8R+/vkz5WXt2KGzrZaTe9uWfOFAkG7xc549
2mFxdKeQfQCxODIewujBPa0Iq1KejRyGbVykHPfUBARz7Xy6opzq1KJNSUCemj/c5ADVmkaWAkdN
sxnKHz4+iREwO/f3XwnCnZ46buxAUii7HOymI1fhpXQjsyLovz7c2CFA802BQqxrrhz+IijX9u/G
gsGA95zgAYyTwH07156Y+UCoE8qMuFgMxAlQqw8v7AZRtscKj+BnZId/hSmVrZdHZ7c205KDjkdF
FcqjB1+0STiucuvHFUpSJF5kwfklp4+OGaUV3M8AhM3ZOy76RYA/xRqWOGaiFgzS1SAS309MXsWC
T1qMCIp8vJ64NOEINkRElq4XkzzcGxwekU9oPutA/QL6rF59Jwt3kQ0Scz1josf4c2MAR4n8ooG6
jBsVsaeBe1BUiG2o3EZaL4TgF+hb7C6wnB8WF64brEzHqxssO/zcAi+XZuYPfCKKp4bKWXw5903W
zCeDzfizSp0QZYlcBFc46kNiGuUpm/j4J+1zeTpSNfyqLVHAq/z6ilj+/Tih3/2zWqhTLBl0iRJr
xP9Xe6ZkQpjRXnbLVBmhTmCFehfep8r3ZrTpHHWzVKqM3aiH4xzvGE4MOT7S8BOFMrBY2Bs2J5zA
UL7AT6KHDrDN/I6scLdYkPKK4j8SDaeaCaiA26BtSDCBiv7NxO9c8jpLpTatliHmxCvay4n8qz4I
EaOa0UozGwF3F6gUseDROWRWFoYMEbuQjhcEgbPN9yIjSndB6a2HWMebpe9Ua0S2oMR5hepit38n
Twnh/0TtgWhAajIlJkf5X+7GYMWV/pcrKt5zm5RNJxO0FwfQcDugZjfZ9GejtYmZh3xj4FUwm+b8
V2DU+o5Dd1vKY+bs4eCZh3HCUa3HnwyqMN9E4KtaEA12dwACSq/ZJ3o+MhglvYUBbBFoY1jGHod8
sIvstK0u+Sf6LJkFv2WHlyzgRuajlqJfxdwBzNFx+OuBgdasbb9zVDryqic2semSYmscZTuBJl2B
yjT7k8a5l7QcucE/v0rDb/36Rrmk3JgUW3IFcWqhxksxcmA6MTKWTGrrpIG9rft11aD6ouZEJS47
g/nNKzq1LplhvKAjrXJlbbmKkS3ns9Z9XqLBAoWMq0Sz5FX173OxdZyMTSNHusT3+3+Wwh9gVenE
ulLIBpYSk2T3iAJ56zer7+NVedvMaMGmBoN8K6+BZUADieUbIbCeYQlYzcReeOPfx9rVVxcHxUny
QEEzH4BMwZhU+f+lu19TqKqsqzAdav0Ir7pTZWl+fIZsXR/qYHXIIYCMVQMhg6GsM+yW9GqXIWkQ
SSGm2I9+uhYkR/G50zeq7AOg+D2pmKNRK8adWcO0EI5Rgzto+1D4qH+j9ljuh3Pxa9hjzYtxf6Q4
yg6hlCW34ZszjHm9cPbKCJf7l72cT4HiRhtNAf1yEP4yBUJzv2sZLJc6WT2H/EeEE7J3FAI8lI4X
5kJRNlDT4aSp4h952D5XnTZvgQ7fMB3ErzRzzOzSNVna4VD3BeJKjQSukPmGT0ENkWpInHbGTudk
+0Jw1CK22ycoWq3qlbptVozrxxK30uHT8TlP2cpcSX4cfUSqg6OXbRRns+jibGLhd7I7/+iaRHMS
WIIeOCCb4K2sWIaGO+f2g+JHuOLPE5kMRQgJNeWDi9cXcwQHtovhXv/nda1rII4lvKI3EVSxqIXX
BWo5Gmi4Wd/xrC99t44Txme99Xlqi0BtP9uVhgQYRkEIeTl9SAv4RMCJRqOW3qWUWlClFMECeQEg
gLqndzgMuOj1mJZeRXJtA+NrBqS3K5bJGf201pEPIOjXMj1uNCvWy/gfoccX2agAi+WFp2g6z0Tc
K0vdsUj9qrM6v8nzCFH+nUP2X71Hzqq9dlFCOB/cW7qLqLi3SsIqcR8GrF9hPP8CLlXs3INZdHGV
EvLd69k1m3rG8JiouCjCk2hvL1R1noWzESlXBKeQg/5NgQ5cwy8xMYL0LqWZ1O53ZVWUspKaiI1k
bzCbyTZdmqe2dlNelVIEkENMxRKe70CKKQNcrGq1Ls1+qJ1t0ujrtJ41UUMbvWHozFBzJ/VjdYAC
hnmvoBAR7gDL2OW3djibLrHj3K1oQKlsYCyqoe9buHr6gTVRv5JDf7yWRouZOsAiEknOE2dXOcqq
rvFP/AgtOYyXrgcpcyanYSs1kljt+88FCCfrYP5UJNYRLzVILffYNTq8pr9Pku8s2zp0MofMs1W3
1s/8g49n7ruiWvI+G5pE31tZ3NuQ/WHQ2O6hn3sjxJ5Zu9wcboVB8MGdQgngVGWgVD9tCaDQMejm
fV/KvaqhQOsQK4K39+XI/++UINGSNHLiFnaXuMsoBy/48ytqTtRrRz5Bxnh0OupSwMUFi3dYJzD4
5a05lUZz8UTdv47FBXRQv+hJZ5GU/ukchX+NRmvxsH1H0fyMObExxEHr4uwvtj2FimkmeJGgWnma
hlDv2Q98NMWMjxGN7uItk2ScPq7OIHqGS/8ECx/DeVHtRY09TgTtEG3vq3Ij1exJElyNF31nwaYI
8oF3tMcaiHqUVfOdZgZtbCeJB9+JT21t0oZkDA5A7EPUH3O9PH7oCN4fXU8nPrl5rCM/kuzoNuxj
+p8vzV4XERt8VTu5ZPpd1TjepOhsuWPwxjQoEN8R/hwUNVxzSjmakxREcpYhznI1qfx7v5m28Sal
Z302wmeT259BhlWQC5urb9LaFQDQpRHD9hireVUBS6rnB99FjxAT38/itJEwgAVUTnJZuLvDiBc4
QmtXg3q+TiGmRIWUybsttQaGtq/5CsGplzEcRav0Jz8zuv9tDbWUGvyw5sQX6kNudnF8qH5UY3Ep
CoeRfEuq7sUZFjyV1INUZ0YEy+zQkTuv2WkZLgN76xBaaWFsK6M1J3f60kwev0MoHsGayf4yj2WY
dwegr68XMz/KifYBpyYHdDRP0rKBLD0letDCV76T6inV91Icgr34pFI7DoC19lsDjzMYd24uDkeD
1li+/oyqpjn+cLaLrKCj3XfbkPBSWjWyyv3+Baci3fnhaUOo3w4fy3qR08hZRugcbxtIPoqnb3yA
bJUYjqdcMlXgXfzdANIlYSQ7AabhqzEJxRX6mA/bhgB4MKMd+O0Hc758t6GVK0px9aTEqfknUvxT
8CcARXSBq+lXjuLU1c65+2jdfBHm8+HcCpaUjara9FGJIa1lUH1JQ0dDjiPb5K5tn792ucvuSuSX
G1t16RCLS9L5as7SwWdYH/MUYH+kOIEGsG+G2i3NHpqCUweWq0ESIdFBsdNGC4L7TImDWfk3AiEc
6TwGeqfsCFMqk6OoeW5mCpWer/5j5fj7KjgCMVqFaF2GTSqzKx79BZsJJRcAWUwRoU6oiDJUv5Hw
WwbZcvfpje35Kt5HjtPXC9KdXb/jlu5hrd6OylhifztJa1A+Gth/i6hvQr/5zhHTQSdoB3bbeGRa
haFtHn3twW90V1eRzVxn+XvDvc6MrizM/d54tUWl7so39IE9EaO/B5GbwgfyoTkHxfU7aDbC8VH1
2FHAgUlOLBxYZ3xuFt1NI4w+RnrDRRqBkbvhFLorwH20j4OldgVfhp9FOp+JUnLZFCxLSAMbqadA
4mdEYrVe0gRiyXS4MSo3qTaALWbPeiy97h0SIvBjp3bMy3u84QT4sAHJa9f2VMX9kaG//8oKuIcs
4wlsfgpLordj5TmKPCk2vE79ZLTuML5MGYANRgOBpLyLfPNNGs035/6HMoeH86jJnX3/lbEDhQhY
8CqHovAIFwdAOro7jR964Y6kHKBgmaef6i8w+D25t6Zy+4/xt5xWvhmzzGcj32mZRZg4yvVZswD5
aMPpdI2JQkzBBQPeX01Ws1UHsLbiG9+lj1SZLnoY5jCxzOSE97r4uZeH9nOI5H4tD3XLA0JIAv4c
6GWSlWJl9KM5oZEod77NvLkiMcXZ3SNRnxWgN8O+/inYIxFTQhqkO3IJawLe9KjJ+yAfS7Ab9JzW
i5phUlCkAYFZXdvsdT2usxysFqHCn4Sl7oveawz9AMSnIFYynYpSmFP8LxAla7lt9849TIQsvCOp
rIIV1z0IeSJVA/ddTM03MYn/DivuJ+qfT0Xw4wGNhq+Idf7AEYKkwk4sU4/TywTgLBGkJwk0ryZa
XCpBdxMXn0lytugh8CpiHagwAwbfy15belNUPSapvnNo21dQPBjlhAE+AMoLfrQB/Afysuf7cTbn
Mk2Q3YyE+K7JQZgy6ehMNvw8pqNAXp12dfEvxdnanjd09szdUrt0WBcreaJV4VMsJ4/fswBiMPqT
tw/9VVx1MlZvRrbugb5evcqvy6O6znM6f4UlrHcFvmiPJ1olVFENXBQWVVrN8aRRDstOmRIvSYs8
l9iDN8FzVnbr7EZqfnIH17Gqe4m9fi6gokQD/AUZlgJ4cqM7wIWFF006LaPWnERJRRihxH/4uygG
ItpdTu/NMYxWWQjrr8zsoey1Zk85H/gAmwnlRtj0Lg1BJrllM4bExya3XZvCS/qTc2LOYi+fCE3D
/JoDCqHwBTmtvc9Svm9aUy7kPr+6xLSnX09M8nGFCNzGVwVYAvS0ymwJOaaBY3K5nCzhVOUasP9C
Q6XpUIPgyuuI9E6M5meDOJACsc0kkbu+yNGzCe0ixkRXimnvDLsfyH+t9AVsPLol3i/2uCPW1Bkw
bLDPT8oOQoLDSAsEoPA2NYa1269HqP5L4QOIzNn88lUwhxXuXCsDjjfEoU7vJdIGrhgEFsPkYuLJ
OjmG+DkTme2/YPS8O21dvJdvncofdCU9cPUzHftxXaoI6Bwr8vNCkwG9/ekVpJ0KQKhtAKXNZ7/v
4x7NANIgoBZs+YOIPgfUvSPEjss2lVQ7+UvutMUU0DJpGvYjJmub7hLeRQVXxZ56wk0Av8Uojn12
H7ItaQ7uHCMrnpuwfo+yW5N9ncZFwFndhjkta1IT4cZFJcvATuPNnOtyuc8dDJIMQGJotVj2uuqU
G/JZBWOSZGkGpncKLcSoDz58n1qdpmUl2T8dH/OeeKZef9G4gFowcne/InUSayHrsiYkspHrVEAZ
xHyqJQDutNw2mspeSpLUaPoC37uO7zOZ2KCKtsZhzoOfOlMwuqJkcRfhiBbKzVUkD19aWO+BuzYf
Wlmd34mxuwSkLjlSo6bbH67m4RCW/XTfOGnGJJneXfhWkhsa1YQZtdV+lNEoKIhIkSgabnNjT3gd
ok4cYn0yPF7bYYQbdRaeaMDhTp81eFcprbqa6gIJebDCDb0lyrDA6J2S5FJWgSbf4UjQfqardodl
Gh9FPwChiiC/9Hzk02iYL5dxxfGdlFGW9HjoB750urYETKTAHW0MewGXsin+eYFw5Sjzc6Kn8zoS
otjgEbpeE1iwndcQXctTEb80/pK6iP0fGdaGbCE2SdDzLY1jvxVE2nJy7nw6+agUehGptNHLTv9O
XEIOY/2SWDxgQZeAvd5nfXbwSz3VHHG0+0OhSm0Tc348BUitfsWk/ZE5eDHYeY12j8xRob5lwoFZ
dojh3G2As0ai98B6KkbS9tmd4jVXUS89Zq/9PjvFVibXY1/DJemH495TVuo3Cf0PXkksKf+79LKm
+IjLwa1azfTQmBynrcxXB40mjHBSdaO2Z1efKQ9hE6K7cddCkaSfQZ1K2QiV2sWo6Ou6Om7yFFqu
kn1FdAp7hqO0xcar7TPd7ctXr8nCEvah6ZdLJRb38tpXQr+jzfA4lC8Fs8VQvqyyUeVy6poPI0ys
voQ8X+Rnp4lC5oHQprHMPUBFmfyFxP3DPpO0Z2beZqVwO7hjCkw4wX2mZG212Y56Q2/o4oJRPy5c
NZOuTW4405kx88yVrty4FOc6WtufbDIoaUrdW2lBJXJbp4wxNzgplad+5qm0HnixpxKkkKyl2FXV
weeKrclycWYrAK0dPIQlNh2+4QhNH7oRo7rvaP39T1inQESkybOixcUNnjax5TE2nvbQT+MPta8f
ECwlKmKfGLqA7dgYnPqxZ4XvPEzij7wxnDq49241BAvaDSB1n7yhhUCKepxu/tSZr6iHGzbJHJ6J
oE7SmqP88iEALjchBLUMp7K2qOoxOvr4vmha9nl9fOQqrBX4Zxj9LMsDvGC/CNSKKlT8VTppWYsl
BWxZKgVDQQAF2I8dSEkxtahIYEi49IiLsePK/NWHz/q8GRV+wS0sLnVXahk/OJxkZSENPTVEMe5C
gsFDugKik5sKjOZhtzgPY0lCY5ozyYeSmAbbPVddjEdpZA2RrC2aIXqg+cCFnw3BiozzjnDGq4Lp
8/EtLTA6sye4aZERMCLDcRvIGzoc9hfBmKenST/Eefn2kFWsSvwznLdPGHe/me9ZfhkGwcuEtyhn
qx1vZiJ3NqVB7cQIV0XQ2h4nlaoJ0I7DkmL4yz8RYibr61xrk9V7DHcc71Br+NQIqe59nE1Uf73u
Q2vbeq6cBz1vQjcJjLJ1RV/tTuGpF8uh/MbW9eOxgY5/01jmM2sntyk3wX6wB4pgTJH60kuQFOmy
rUVsjCuNtAoeLfAMimFwkt3evqtcJG297Aw87zsWahUVH1W7rfdnIAm42gpBGJD2z9bIOmaFEoLD
CeI1IhKw3QLbpeZVz8p6P5WXWOvHDYgTWJ4hk4sK0taw8ZsFd7FL8Xxxjb2gZtrKDmbosXnupGbT
iaHovqmtg5P1GQwuHjue0mHnmD9nAIis3/4K0SJfyfQvSr0cIpsZE9wEbdLlbRY8Fv6D3PceHNia
leM8AxB3Wjk6riMWDUv7vbQSzVc+4C8CMbZvRi0MV2bfFs2qxpAaqjR9vktaNQMCuoQTbzbiRbwe
mR+XCRMAE3CWr+0ruAhN7OfsVTflqv0GPcBPxngjKyywtS6F3YbVM2MQJ5QwkXOVC4Q3sVWKR6nY
N71TZAotEOYl5HFlMd7oI1isJTDbUFZTnKQG7kSdUJvESRhSsar4tk2d3icOKEwQwwqgk3zNAVy0
AjioN/CuBfgd9Eo08I6D1m/rwJ3WqgvnrJV953+RfE68pwUaTBLIezp/reckON+bDTIbrQSPvbWc
T9mwKfD6t7ZzNw8/hufx7dfrNim0WPioAUvQPNfkqRNmymOob2vMXKqRiBwzF40NsQB4XijtByaF
s61ROq1F7vFCRxu++DjhJrs7MlRKqDA4huPkdBZYe+GQTAxwgivzUClCVN+g1SsOt6nA5BVykWFn
tyzvp6KbAFguOaFxLWSUltYTBWyTifzdd95VqfAnkuMhCYgosLlD2ed7/D/BmaWiPUd/8gYB9MxW
s2LVCKV80fJ4lsy5771yMoZ7x2gwUqiJ+DjDKUZkCRB6O62QdDJ8NEJRRh7Q1NTYyNORKmrU0NGp
RFfYXzISBqstNNz2Oiqu9nhc1cFdvC/0x2psPLKKlaSZxIju8H/3W2Idhnq630l0AhhX01Uay7Lc
CO1sdIaSYRCU90n1XTowjfGk4ZAxm7+kAFFbgqkXw11kn0EjnNzIlcytgny8eW5/+ton9yNfU7mR
LbBwoAIQ92obUIUWiwq25OBiflyG6+3aQrXO/PrVwknpyVOisytx8n5cR0D1U6y36HTSyUFM1zOH
oLhQx034TmeMZXfLz7LHDXyftZ3wfiRjJVV81tRV4diPSuOOtpFvTJ0AxOh5kRVnUJ+oOKH/AvK+
LscQ2gYwpN0mnIIvNNssIrQG19Nh/eFO7dsygjlje3ygaNelV4MgENNKin99xt4wx1rYeXWaICUO
2MKir6tb34qDZfeEcY2lZnc/TiC6wtVFAa0wckyrSuMwsEdBl2uziLeeHULUDjqcSH06PUHJQg+2
e7Md3YSAWH3NZLfZoGxZ4VfDzVO2FyqB6oZllEbE0RYurMtt2r54H/rS3+SBdMWR/rTy6l24COXy
DYuQ6OTy9j5tOeagOY/+K/l6hoQHwlB74QUyGj5J33e5XT6RCMazYxwUFfhefnx9yjuORxqlRNYK
29cIgZSvENIUOZNKvoROhI8CADmMNXpvAf1CoUydMv9EtrLba7bnnEpmDTRzGPlPH/TxjbEHOjZS
BUibEnYm4TLojAKt4xnMogkI3CSoSaZKHAt+/RpSNdp61ZW6tkdAy6wt1P7i+fa8XSvlR+55RMrW
7/gpJ5T7O79OlkvL7FBbnGPD/gHiyBFf5kenlBfh29BOsxitz+vZdB3GifuChOQPa9sgeGwWVGui
Cz39Kg1iOOxY3QlJD88ynYcZZOf7iO1v3HorAIlYhsFXKBS/569JnH5SjHaD9ZcF16lWWF/J2igu
V3VWw664lK5ueQhy18EpRTnZLWwLE5dPociNbh/0ySfuMLqlcSyoLhpe2s66hLKK+CZixa4pevvO
8PgWZXupyz/0GtwDuLfmMQOImwCLSCbd+sJQyhtyzricX5o59Qj+ap43JluLEA3pt2qwscV+aT4o
o0kEGvvwA6AWVtw35jmjrG0kEG4hfStr4bEyEW7is/5ubepcPj34QLf648EZ8nZ/R16Lvboq0B5j
balErtuTb8aDAkpdtiXm0VkGf+6AB2tm6Yy8WUXs308KCLodvYtvUofl/A8/rAVKIywjMyUeN9px
MUhSx+YcuhBggOq8GbsRPfPLcTRbE4rAqJggaD5FEXUw+wG96aNtyF7R+sKBOO9mgnMYMcrFgLNi
nhiKmkKyrJi4ta4HamYrHh3bubcov5DjEnIreK4vvIeCifYgF4UvGgLRYM7X1UljSfbzNo8gHFpC
0pXf1almbrJQ6QddSXXIqBXSSG9/ZHJLANQnXhSHvlPxszVp/6sJIO86ZRa/m0fBE6QN5ZJ3F8G9
YGeZejH55qXFmgh6BXiPFGK+i7QH97O9bgGnKFZ3CXthpz6Dealo1qYA42nAmOeBntuY9Nqd76c9
w0GgMTHacl+I8KywODs37waoddS0195V5SwVWYL8OtDJj2wUiLb2hHzaMJIban6/zeXA6GS6Rv3q
uwsD1Ty6fTQv9r8HMYNPRhIKs+BpBWtpIgHTwphWYck70LvIJRT9jqw5O40N8833X0LOwEdl2xXX
wyeDoAYxEOHiyGcWdNPfTj6yzJaC2FlXJRFVGO5JmBpgX8L1fub+taSZrkpwqdDlwSeTsyZ4yTxE
DjgIi5sMoXNfoF6jn6tDjb6GNvgYjUtcPyzpFxSYSzybDCfp6aFjie0pgTYp8MEUmQy1V+9HBV1Z
Iz61WDy7gGyzXtUFFsGst4KjNvSGfhwmH8s1WLsMA3sQv+kUlVLk2QUDiO44UFAs2ZiWoSKngW1H
YLZuBSjVfhCALNuSEp/dHiA8K1Dx4vIWr4vv6Mr/liMHFySs0MFfAdzHmVR1Kb5dkvSUFMcRwxTj
ICx+DwFIAXr10CmAf/T5YN0vIrqnRU7IoNbskgZJ2h121DLuG+mbjGHT+Fcg5p2V6/QT4unbGlMB
zjAclYA3po3b4++tPwHZweh8FbLY7vewpjh5Zo8W5ru11Hcm5MaAzxuyCGwIWfC6FDhwrUAOodWS
2jmOD6qPmfNPgFz0NCvCMNKq9lpUEuhli5vNikDsU+1VcPNYSiSxD4EbU9aXb/y54rbxOxzXgVeX
hKT36s6Zcsrc0YZQOYBelsPzOkttDpwjROY3W+k7Hi7rIcqF1V8ON7RR2YPu+xgWD7ZIwoXatBX5
8k+x9E95WuKg8HdFXTPOWdNIs7+0RKbBpw6/gdy/qSRGsqrjAYA4tEtl7VU22pSXC2uwgg9mgeYu
zJcH5yxgOmUttpr4VEdsEh9FZOtUEe88gnm0FR9soqrDBjNkm36w0cLPw1jfWzsdusB65v4bL+e0
ebRweQuRT87QyKmq5R2uYVYdi8th4aH5k5xX34k9efCph+Gky/+IxhKOcFYxXMj0UTfpcx1ttRul
ZAoxmzBmiOZGSGZTIjdRi7wunOIjXmwvcRBtBfG0cmeSdpBETvuHj+v8NqeBi5Lk+d06c8lbmih2
fYX5HZhBDaf/RwmlN2dCrXF8JoBKa/cviIysjffFyc4JzDTOZQqYXL7SZ0FnxoAY64n5fYUndWpQ
wPtWzZ9eA7rv1vVNTi7zRWQzPcus47ZLlb6pSchnv74atDFKCE086JUkg8LTVbtBSawYAZKIxKue
MqeeOLO4u3PYHsvoVDUOf+yY3HfnSEpEiKucK5ocXRiHwr8NYH5aJw9lw6Ai+3eiWvmyyraqQCCY
nkrNSiUAI1IpnUvoFh35eSfnrb+wyP0l9kcHf5orZtlXZtmRWNWKNT0RNatxu5PDmN/I9iMVaHA1
EuSsWaA00hHtH5rG2Q0YltK2mN5K0p7iFk4AZXXONJIwaaX3f5r+BW2uVHzDPgURQr6QzFLJPx5l
DJpkpc1Wk3Dwtx1x1LJ1gcQIClmjTE6sCM3Jpg0RFjL/fGr5e545z2Z2IVD9LV6pVK+mDqnoyCwg
NnXsPbwup6sel6hIg2VUMZoi9c++dTeZGyVkSlzNEeQsrgSWL6u+pVHPvr8sw9/d5dl1qhqH5pqg
8RZwJj9fmJ1pQH38cJfyRneU43Zbvgt+Xz9vam9d1TbvcY5l6H261LOZoVmUAFKMATMn4Lmgt8ri
ACt+WdwNCAppEPYg+4pdKA1Oi4LzwWXpZdkMy3gaDJTMbvpJIV9V/OpKQI73pG7i+Z+0qlEYif0M
tHVmXaPjT+z3Tks7UL6xXa94BWCAyTwr0eJzario4J+Z6+LEdlJ1L2rYOd0nGM/Sge/nXzjvaBV2
7Ygvf9XnVVURfRIGATf5hpe22k68dqq4aNeC7+rT/MoST1V3OqzFUJLjPf3D02Z3zeJG3MQNY3sI
dtHopMdcrCQxKTthNSJcwm/h1qskYzz+pzR56D+Rpj23mQP3TUJ7BTfmUXIwaHlxG22MuxnfN6WW
jlcq7oRZDlPGHaB0nkLOrqMtb8vdr7PaB/p11WYnyjakvHsPtn3006DP1bdWqMXBnppTdZ7LzM4u
8x3NdnCIdNsG80eIsk5mGXyutg5RnZcPIdQVg8wY/iwLQOuBFh4kZDyc5lsHxpFNhx29ni8LJlN2
M0MMNcUS6kgzEAooiptdz1knlMUA+DcyFGSkp5+91hhW8W9GiR68Br3Ed6NWCOFCiwMG80tWjnA/
L8oJ3JyjgffJTWGyYjnVuHDKbK2JfRcAwUeDbTm+MrQ9njjdMf7RB1RtGFOeol3t4xHV46yfP8Ms
B15wPb0Xzb14LFbjWm+vuRB6YwA4sz85BfPrlgMkHr4brEuZD3lpvHQaUbGqXyfaOqJnqsT7u+Ex
PGk6yZoOMWNR/1whoAACGNjbxN0E+nLLD3LjbtLFASAtWQIkoQ4DB/DGAJbMSWBTPWWgcMRGiFQF
xQoz2ZtE0FY6Wgm1TKNong+35RHfqj8xZp2s4WhtxEAGbKae0fPqe75vYHBZCoLY200z/RI8q+zv
lnZSVEW658Alhf69hymsbzoUKH/2d3LIgpnM5dI/9kviRfnNEtADXLwnrcUoG8y1TIW0iHKUahOZ
HkQ8j0zkFQoCEl41oO8F9XuXQ4Nv9dFDvE43w53HYlWxqojzXWqoDBF/ZivdVYT9MEgv1DhX0O3c
9qcePZhRquCFZ3fJwzBlhWqRBbI5ugndCrZIYhDAntW3kUcNDMJrr9JEwk7VlskhBDoMPMuTab1x
j9ORw594Jzi/o9B//EvCrGH1t8nrBlVTctdVrpgwOmc3j07/8Eg1C0CUPOYUubqJ+L/zMV63Ijlj
tnBlPNdUZ2mTajj2mQwjjaND3aiwOSjtwXo41W2tPALPGZkeaPh2RzUPP2/hYEZV1CoLVCwTli4I
8SCgYiaZEgB79NZc2mRD6EJWtEXi/vCHrzGyMqkBi3PEKQiU1KajY8YiIYVL6rP0gFLOT0ppo3m4
LbgQVfe7d3KyNhlAx3jpWGsmuDIjY6ZG/+BKWVfqT5ySFN5nzYXGlC29rnPETnhls1n++VU3FQGB
Ml3K5TCUTBgiK6Plx6pYgGhDyMy+ObvDyf9Ua6dDdaTLSgqpj0Sc94PKD/k48pffvpl/nIpBE6CH
n7gbYtWfJ5WnitLrt1EjDq/ggCC5cfwwMKCk0StOls2LpdEBxUIErrBDsaNHoUva33OTHdC8bFwE
KUlDQDAxU5tDHhLSEPuZznVodbAavfn1w699RPmejjsF0j//4c/MZxTrQzpVpBCm8/JFRLZqJvSY
z/p7mQr12JEujGgAv8ZwI/T03QsJlNpfB0/hjRWuPsivnYq0XmdzEOPSYHl7imJ3uYixWFh/kPak
Bo+60q+CffTUkVnof20M4qYbd/fakj61MgbNHZcC9HtOGxzsYZJhbsqn3hVybtrARGilcn6eeoyR
FZIuIDY15x39xNB5VPVMBZ6jF5zbo4p/2ONsp10tOEBxI3WNMXE7EoWSr/2rshZpvYbBG+yFAAtE
FDbUMRWWguSOIUGcj7AplH0moeFo2b+G7AfJQad+R2AI9nw37dRVKDOQomzK8CvY7RTVSf+ZptrO
jGqmNzbTyIVKisAZzUZhxIu3+7XTJEwOVOBMVJnYe7HLl9isMr11WKHFwrwBFrNv1uSgRtyHnDkl
aSxFnIrtiOAzgjLruhpFo7TeIjUmBYPCi/mRz8lejYzTpM85cDzuFbnyZoPr9WiuNsYwACXMjxCR
j8tZbALeGcNz88jLEO/ygQ4PeY5LNNDWp+WuPCArxVPBky3b+ALEnjhPEiBOMbfq2DD+bSDO5z4E
OicSamuuTC9poE0X40V+HxCye54GgJTS9pLSuQIsKMqIYLyKpKAVSG1Q1mEUI/O3Hm5EoK6T/k9d
Q41sdsZ1O82BApPFIS5132K5RC9SH6q9nl4SkmeWWyKw+9Kmeg+vKbCthsKd0Ia0GMbqt+2KDoHO
EJodZhBtanARn+9c8rerxke8D0RyRQJzwrZHsCxEnwt/Xa6GxKUT2xkZemkN+Ntp1IFHpU8pO68c
Imv7uOyaW+jiin5Lxrpx/SY13sehH6G9aCZ3pZDY2mDqa2HxlSGs16xHjZIE5W3G/VTghR8zvB5Y
K8lYwyRYv/qRdS+jLhw69AgDhCUMciV4WGfxPBnIPvKgyzHeujnL6qxjipibdza6ZB9+TZG0aVcZ
mFnO5lXQLQUUKxfbyMepUi5v14Ut/GDMSkFAPKU9JMzNLsTPmPbTJeuga/xyXoVA4ffkEG5yhMPO
9RQSQy9KcwQqm1uxHZDKq84n7obN3TbYvgG2wRpK7nIceUhhC76ZF1iuY+4s1rCIOnUJMaCBubLe
IvEMRl9Hkl4HS0Wy2+ANu2VfjHN60XKM9SwIjhzxrmDpvqWfa2j4FipCgDh4BNjb0fEEXXlFLldt
kw6debjg+Z76XTDAex82GmclG0LUR9BMVYjf/Dx+Ngp3Dc4qWG8lLe1HD5nxkeB1QrxWGoCbEcjC
PiqydoiWj4hIjzqyew6WbDV5KIwIn47xKOb658dxOqCfHOV3xIxE/4+ptloq+4j5Id2jZfSRgQJE
xV3XlCkjcSKPcpJrEb0nXSV+P+Q/KTzYfmdlGJXrvG7xdrLMhh3awUeCYpJhAtnyy9Xcw6cdBIPb
GxVtjDyrdUg8kLSrwtr+MYNgPRJPSt09O00okG4rX7VZXfsFt1t7087syHgjxEErTohsG7drQ+sv
u5JJxKMJrdSFPytymiOF+oWGHVx7G2F7xV2FTda2I9fncEY4XyguHUFseL+MkuNYxt+dyOdLHZRZ
+XjR0Mc4bQH3sSnlQ9+9PWIomv2Q81zDtjrHDBmaB8/XukJbSwp01ToXn18U4cMDehPVHPbI6tnB
dByQJsETxYQ6EbBBXsFskyWnZR+q1bF1ME/jX0AVU8oFF45gOtzSKerlduhTpXk1ZDJwzEZaKD5E
OtwaXMnUAi93UejDYmtbgSZFZzEv1rxfuzuSO0kHD9APO1cfGD8L1AVcn8QcXNCOQmAwjeLZVikH
kqgpL4NJ3Y/6VCTX86UcH0Og/6B8QN+vD5d7wHDk7CaFoaMFpdwUd9QBt3F9yyfhVT5BPmKktIeY
Id0m4w528Th2pK8K6ixYYV/ohN7BjF27cO3ear3sfVzEUfbfB1befmqNxM099sq0JT4HWWD6zd5c
5NZwnlI0D0s6cKet2crTTgUeqyALMAIQBk8PkH0ySN9aXWfRnnPbI8xb2IGR5CvNshaComdsuZ2X
hLh0XxYLfNGvrfHo2XXFEoAe1kJflZ/qZdr38YQo5reSGuWAu4lcji6TM2MIpmRMN3LRPwWmGZdm
Bg07HyrZEcflULMtxLFvWFp69fQ6O4fL3cTHcAEouApP9h+zncwuLlTjjyjGI2M1wJWboGcaMkDh
g8wlAgutDQava1Z4ntJbwLhplvk4TzDrD7yLr5osKI8e+4QvtEkeYX2fKh1HdKdKm6EtIfpKrMoB
WJoicxhdrFo3NjI4t0Bkzv7SnlfsiT7E8DorwwnwtwCggExFNm1/utOsY3TBw8VqHzp3KShF+Ba2
sy7fYWA7UDW3RKyFb9d5Uo0ASK8tHdFvRRdmt7t6yv+btu0nP10y1U2NswSDrwK94cYRwTnwf4bz
y+MwAW9FdlXKTuAgl6SFD040i61r9k8RAAZ09e2UIwoUJboS0Lhd23uVXHJbAVDw3rYoTckkzDiq
3ji8/l9WWSBCmrLfJuTx54eZoIxEcYhABV+rxSe2eU3xw8AmQDS8CXoyDsAYOjVJVxtjXnK5m+TQ
TMaUNGEVdx8A9UL9yPcKsdke5ou4jopMZ0k8O665Pj0HRlVHZFsZCuVBz5I52kwTQj5+d0bVuYKX
EEfiey8xUkdN0aXoswizdGS8u3WQSRfVVZAilaY23zCUeyZoJNv0DDxm1QGlIFDPlSRo9Lx5TRe6
7diIcjB6bnNv07l7TIdhDSS/Rlva6Vr2Pw/Q7f5b7idoXwk+LeQXAKLh7fJRP7Ckix0im4kERbR2
WtNK4FNb4Bv8iWa6PM0gTtA2kyLBV9fYR75RmYcSFI8n2PrBnazd2XNniCtbBRDhyuGPj5CATXoX
yrd9JJGwADAb9ZsvJnYGhBKwIffW8Kn4j6llTZznR1Mfpd5Fy0M/1qfpbCsE1Yzh8l3CMch0Dr8c
Ybo6NzQ+BUl54Fskhk/ykrQThANyh9CaOldJa7ePN7Seb3BSFDvgOpJb3XqMnXlxmxghypHaRCfQ
aSvM3hlhuIfRZoKokSjHb91e3h14jAuptJqPiCGVwFLFe93JmotW1oqY24yxCWIWc1h+QXtYOkdg
+vv1v1H+9WwFli/GBGkk1tvzgNkykOS4NzEpodOvBN8MLsdt6da+teQcykD0lqSoYZkmqjM5wC/h
mLg+6I8u1KsuOy3cYpglPMV39I07ezHHe2Q29hH7sEv/sqLaWfG+CshVJt5ktB7MBPuA8EMQZmcb
Vlu1Jcsm4CNg/5RqUCsGq5stX1O1YtWCoeCpMKhlsdoz9U+pMVMVg9SYv5VIZzGH2C0jhteMRqut
/6nMUFOfjzco21QDMWMjHITsFTzDBbWF2CyoprYXjqgGh81D51uQfe0JDeYDK09uVjUpoqMF1d1Z
pjySgwU6eHIsFT8LkPEKGxZJkGpn2OfAqfhTYggUxHoPlyZtlbXPvjzbqwsL+e1+o+xde8nEw75U
uIrcPn0r1cpi+kqoSsdGJOhNuqqMFQByWmIr4jXVyewCV0bQngdY5+DZI04IIIwG6bWIdGBVe4fS
3RkTWhb7nIFoMMw0QUcOcs/HnAYhnUffcUEH9Q3dMEK7LxqgkKpkSTGacew3lRA1w8/rlV7ckRUa
wCDaAoUMxMnYGD/aD+Aozp2pGSYwM+5JXviNL7I/3E3QBZ5qyxMu3Lsl7HPAeO3ZL0cewST8Kfx9
r5WMhHR4k5DlMPvyMvNLFkuIp83+ryr4oX1ji0R1yemnP7MtLmkS3UDZi8i/EQpNcVzVtmNeIFbf
gmML4th4ygVD2t/1BZoTb1PPK1xz1X/QVFZi8tSmVTXwS5Zm5J9c0yExKDvfoGZQ+7DEOfUM/iBZ
x6HZK66PBLbad+JPSo7mGmBxQJn8rej8qTtA4jd8KMuJN1thWRRsOoz2MmbRA/ikV8Wg6PUfG2aO
m/4KPOH0sw7FAAq4Iva7CHV6TmcPLI38VDqPUM2jKt0WaohIBZo/urvjo1VKF0m+/Lb40Nhi/TmP
mw5HmdAXjKY3m0kadmzS1tqApcaLjWgs/Q8QvD1MvewQfy92kt9wQCvlX5o97f0Di/Nz6XcX6RA0
Qa85uYSqCBBaFhMc9GrA52zWqzNCeDrF2XLytZ/4lZ+eviHR5vJrt6zdoOQTrSOhjhDfs+izS7j4
Yd3hLE3Fd6zoUh+VwXFQGpZ/J4wmZHlF3YSrn0EfE0fLcW/KsSlJSjYgmnRTND4YXzC/97FtUfj1
bpg7GYAt+U/a+SSXF7wwk6IiQa5qO7mJSedql/6VCwMQGiTMMJMDkPC0h+LaIry0IxUWRrMRphyh
KeDa1mpXoRB5GL1jlfIATbo/CUhltePtpqbPSoRC/BPHCh+YeDU+0SwUqXJihtFw13a9RDUA/t/j
d+N7vlvqqOMH8eequGc6yoR2cz4xhXC8dh/dvWjapKOj8EG2RGVqK1dVLT+n3xlYoZVP8o9uRKlY
VuoU95yaiZforT9ZCt7WxeHImZuejNGaea8/sQwWtUW8KPteSYlcJJuZbgO6wO0nfOJwIuKNkITW
iT/XqYawUE607khGy5QfLvKGQFs8//14UhPVARScU5Ed5MmMsI1g0PpTxaWO8INjXE/P2juiGHFm
aT7FGts7imuJDFonqA8hpp6eSR7m7RCE2KeX6oxsdw47OU2KlXf5gsImTobuKk2dhB/k0s62DUIz
kojOC6Y9LqKqyZMzFnNKEKYm4G/OVwy2jbrOKRYiFh4oyjukmMm2weU7FAQATY08KrJSXuWlv0DV
l+ME/XuxrUzqhCpxkfniGOcWHO8TuAWL02QDAEPMNQzk2RmG2V0Pcz2/NX8lK3ReVHRgtrI2/i/f
GI7jjVF7g7C9xWcVPTxf4VNrUVyvt1N++ce31RtILpN6EWVr8YuVXTv5MCQkGT9v9boI3GYitW0h
WJrJpighcUnQGDR4M79O8sTk4Saku+L9tkZ5saL+gu1FWMSj802l3PwIz6aBUmbFy918PF3thHfd
+4u32ZwuRLGpFDgY4q+3LUbK5bu43zf2z5TLGtQ1YE1X/dzOFPW000xvE7TIaOEQGz0nHFNCbhDl
doTgUryQiJfGHfj04pWZkbGSlow7fChVV3wmwc/Eqzc6AeEWAyBF02aaoK25IgUwk0QQviLcFVC+
4OiLQv1daDe4miJglhexjO/OUPZRNJ6jfvCDt/AzQw3sPnMpwIc34KxGzPXMxx9UZwyPXrOfkmIo
0JOez57h7i2S+0fDBjwqIoXQcgOg6Av2QvjKzLdb2um+5Vo7jeKSD1RvCxj37Ndci0gEkqPQNpb9
hWiq8icejh2wAaqvJR9iQYT+frrQOOuw1Fnm8Kat24x8MBilIwR83VOjcQBXTM10YTfjQrqjDQW+
4RcRF68YPGv8ZHzv6tB48ba/vjMd8k0tNiTB+6ZzyKN77QoCDJC89SZeu14do2vJMP+ZpcV12DgO
qp7xvASsOGJFt1TOELdnMse1r0V4cx85Uivo0X3E/u714XAERz3ML8P94CuXMKbs1n0LLvPrZrhi
9RDc/Qi9vq7348U9TldFT4ECErLAYPhaI6MYqjrz1IAg1ljtd1wKuJ22MXKKQOGhGMNcNx8Dc2KU
9zb1jcNBv+ZwOM7qJF/Uimv1vsbScXWSNyTIdhdiVD5LuWIqcuu8pinTnqdEhgTL02W3UmFZjA+X
j1Yj1ti73lt/TZSewDMtHWu7rtjmMZ53eXzAlJv5C2pNSG5arImIbplsMlFZf0zsCQuwkj5Uf9NB
kRqduyTau28b5H2mEf0rFvtR4u7DDYyUortZelhY/qE/4uNg/cwJNspxBoDu/OCzVWsCC6Xj7SCi
S2OziA0hJqlxvnvuxaZ7qYubA8VeG1YVinh44K5TPGF9DNysgTESAqLleZSFmA9NrvoXgY2MTnRo
ap2AUbdSFmGeXcDiM0naZX5YAsHkFu0zlmYzMYbah+FVfFQvMDin7hyilOZBOpm/fBZl0JsWz07s
Txoecf0eUFRy9eOcDwnyF1IHhWUXst8sI3OEsNsfwzLJIso3fteJpPQa0Ij7DUvME+Z8ojrqhUIx
lqJmRVlYjwwCDXpiA7MRZXH7TnX7og7TFM1LIoJdp0vhchtBN6256tJnZCTUOuYae2mTYngf7eVb
TFDQZ26fcsMGXA+eI4WJoseGVOk+8lpqeHfhdX43Uy0fgoRO8WRcq/1f5czlymyCUGRttO659mmb
uzenB/PqNRO6EcLe3ZbX16+EZFfx7qukFekTHOAoqt6P2Hbh4Xg36xytDwPinwWBzs0MVuzXxBt9
xCekubb3+df/TsvVdNAFYfnEEIw54Q3cuJzhFqXHM0Pj9f+vvRVoLB1bg9Vp9eBlgH/wObj4DdmD
bHnkcqrCRHOHHiv5OAeYp7iMgP5TPnkIECB4GI1KrO0C5oxX+XiMiB5Pj3grB0/63SEwBR42Wrte
fgWYANL7zeGuNNvPfqDSnjedG0RtaBv1FGvjtfMfhgYRv/ZRrCuW0QLtYcHhiHQWN0pR6VfOhOnd
4PyV3hOOYfl+fqyjq7H5IAPZbdNncYRvItyzkyeoczztGbRgtylRl4u1GErlcl6fT7xz4iMW7XhI
177fAxGkJ4RxeDimr0qdH1BGHTVG28asK8R5EDA7V9/xeU/X8N1rwwR7FE1T8btymzoRrb+qbTje
dvK3bcN12uRgxmWwwzb29dvhO6dT34t0EsN3y4hF3V3F5s0yIIk058qjMjRvz6wciioa5BfXfrsd
T/9gM5SeEIgnWwRe2sbbVTHCBwkUrt5bkraW4Yh88NPceZAMpaTkDW5imSIq3HwwjfP8f5BOaUZy
3cddRzdWUqxzuOZy7BIb+qxtUjvOVgOBoztVV1EqtriYJlU6VRIgtqkLOgtxx951/hOmb34N1E9R
2iE77ACfk1GYckxIeai6RkGFpIowdiEJaz/etE+LRrvhXD64ebt02QzpVyL1jXFqM6kA9Q2Oz2Bu
zpC6+a3WWs+TXWGjc7+R2m/GoXBSJr0I6A4WO70K4Wg0kgnRQjfhItR4enEykL1XvyAuWU5HoZTg
j4VQykYJ2xCsxrLtVS1s42cOm+q1N8iZBTxyqUuGiOgY8R1Lgh8uIYnIrvCk1I/+qoygtbDqLCLb
Xk0TwuooONJwGoqD/au+tAzwbBgvIXaXUEpGBm6cyffx1tX+NaGW/SgE6D7c8Jju5irrV+p6WA8R
i0HJ0IFnrI3Cy49Z1XJmJjIWdX3os7OyjEf7x9NmS2yiN98AAX6ZCYqWRfn38qz/9zJPCZK/uDjq
uIKlbDm762neJhOuEWxXVi3U21jjOLXWOwEoq5POsDMmGjoAdEGjpbeX+joIkBKV3w3bksRx0LL5
tDUceV027q38fcTs4QUx+UaX9vT3rDRAPhe8Wa0WCt6tmGaKkOXQHYF1VCp1AAtCSRXT/lB4Q4St
erWrtJUpqvKCgWggrIh874a0Cn6JjRCvyLes5iMsIT8o1oN5Qfz9tBnjf5JyHpjwY+ssIw5jj+pW
BIu3NJjVJkRQLKgVMDmgb1JDSK7vbrZ48VGjfceMiCOIC04568GYcJj7MgTI/RLbi6Zi5q4L2JZO
6azLSzZFs3wwr69Q8rQlD4WGWRcCkq/YntlC+512gLZYar+lziRLaStZ14jdmgC86GJZmPGulL11
OS+bDY3X52V8muZM9atz6Ab74wPRmk3SaCHpsfJ24gyuQK3Z/w1yGtRrWERBZdtPdvz8oHhye1b1
HdEijNY0hARnBvT4FGH7vWgBc4oA+nGLJVDLqDhcSHnaPniCX/Ey6LyX8l5529P19vI1POnwU5tL
7SkWsqhSY+o1R2Nar1RMj/XB9Z5doiTZehZ4+B5+VKcYVekNShwcPUlUynGzW0i7Ph2wyVFW94Vi
td/EbS1Y68Cv9yRAg1/r03Zlq+J9RxnXjKewU2TK3GZu4O9k3S/ZUWB0vlXl+TtVoZYO9L+MKoMd
3IKI057wnoXn5RuC+xgt0fTH52Uat5Jqvu3CuQN+uA2LEw6eMplFqcEIzFPgLA6C277YuUumLevl
OUk2GbF6gqYwzosi6wTmkpqtQsxg3OZZ6b8vaRD6xDz1ByQtKcURNIXvZhrFrHwd05JzH9tgDr0d
DgI3c7rey/YgR79x9oP7YQsr4i1RAEwf/72c3kPmEoAiGu8N9j0oEBs+c4Hp5sqdYvZqLmifjNLe
XAjT4Z5ZGnO+WCpLtrso2YvFi3tKZzIc0IK4/cQJ0btahlUKVlFsUs9c+WSkLbjzW5rkpavrBnp6
+A+5zphBmdlqsYZ2C/4ooJPRvYU4oksZ3x7trdOzhxI+Wb5bP+ETATeFKKQoFKQxINJSJBRaYVzG
UrQ1uarsp4WHyEbHyTDnC6ld0QittJ38AQDsWc5UrWUgbTOVlDUHn8WH5zQ9QRHveUMOqdzwjz6p
0vnMtJmaQJQ3RI1LW1Jxt6qU9vyVm09AgfvRC8NSg4K2e9yeaEScoY+5ADUiHTzmOHcZVeEd2TAV
qDDkJmjQ+8cviiSuf8EZUlaZ2D5V4wRdA9PsS7yfudKe5myW/1u2VPhiOeeILP/cyMoAZEFeciXm
fZtS+4S9QbF4ZUw1h8q9Tqqs9Weh7fw2DrzPekK4Mh2QEzPL9NxBtiiyNrTUBTlMRrgdMibiY3A5
s15VPXMx+UL69duHn+ePua2uBOuAUzUs0gJy8Y7/PYrkoHx131JLuQY20NvYIf/mJU+tWdUc1VmB
JXTTFTjJNRx1lUgZPo7ef2LOELQUG3P5KcAD5YYJvDDCw5HtZQlWXs+oJd4im+5ZOr8u1QWKt65F
G5D2/g4y5qPkDZJLRZGhfWh2DLZPWRgTEs2DP9x96mVOIkfJvMJA2waVEvnu8uzs1G87se+ma9XY
Bp/swVYCL1rUyWsYx8QUT5RS4n+PF2ELG8uCBSOp6mVBzSQf6g13aDn3r9UoVqb6Q2fZ594rp0n1
/kpkaBHw61cIykEqSRtvRPwCqJX30q25Sf0ksjepGrNkGEmgbLoZ0CIUCVr+gmX4lA0L9MaaE+o7
g+UwEOIK+ALydPsCoeCqjzj+uGMxx/2WnXGIAKPBejfwb+iHw/7MAJtpsW5TrNj11SmAFKbNrfnq
emffpEzNnXy5yWjsJ+Qmd+5rskdLHNuZo23KtZRACVeL6or5Mwl7Uy9j05ehKcWS3aLTlFx/I1JB
eS/WcUA2mJVWjKEa1dXtxdndrGd4CNhjLe4hmEVYfpYNedJWDjRDECuZc+RYUWPKjnfMKqbvgkoF
4RYgcXCJvLmMwnRlNYuyM7x2pU1LDgmpgROrSEdM/ofmZ20O5tQABnLsg0LHTHVTdX1JN4pnCAuz
1D33+xOkMbIBSQNIAc9y80SA4Py8lAZNYgX0s61CVuW3UIRAOfsAFC6exqzW9/sOECVJPfiRMGbq
Z4M8K/FK7g6dFLAE1A/Qh3AVM7QwuJfUCZCR3MARAKLM01y+1jcKFsbJkq4vtUU6RkdLQs1SNfpL
lct2QNPwTOE9zetiP3bP6QjviZoYk4V4EkWQ56MhaeAC9N/TpFsAbVPWOwZYUKDsP0p6rNJjC8OT
1x7bvP4LHr7z7dbNNPk4W4CzdnoIr/YZ6jFIsYnwr5qXNLpKp55pwoJTZunm5uxXva7PN3jFPgJC
fGG6GGIh412b7+6DJv9SFM0AZUb/MjfHC4IBCOmcIRUoSVM6ATqno5a0z8KSX4FqUzDe0tUgqRAX
/fE3LwXO54ZaeXnbuauMdwqO3Qry17BCJdE2k8g65RHFXQHGyyc2pU5Pefci0SAGFf2NDm4fdb56
1wCFydNiLIE+EtcDO3Srj/trCHpYFustCzsO2Ha0bEJP10tYufDOKw9xJshsUKvhj8idZncBSXMa
2ocBQV7819ICKvaD5m2AfeOOXiZxJ7xo3msG3uXEJo8v0mPBHssMWGWYWHG5jg/FxVUSqZzEd5+I
UY0pIcADm5xGg2oAY4Szoavzf2oeyOVCbs3SOZUFZhXsiGVA6PETTV5+O/A499kmzhjgtHyLDNHJ
M6CCO2Cbff1/a+kbgIQcyYjt4Ayds1LDW8FGYkDPZX7iVZHVgCYRQoKOf9FgLHmNB49lDQMF4gtJ
4l3GZsMgM5NeHEqVfw+mcyBvSdZ579/8/lZ3FR4aAvkkGMjZZkdEqIGzOq/L/YltK9fDLHm05NzF
ifGvZC1cyidopO6SOkeUdiIsTc4duXLhJp/Sp7SxsYWMkj9kvHbsSMWzyH/a5r3xpJaPRQdKUUuG
zZXFoqeGa3i2kyUtQJpTrNrhBMCcH7vsPpPj16fV6zfE+Pn0VHM4EfrmmjWPCdpOrC8bzGbHa3Qm
TLLZtz1zE+S5B4aU66gpf2K5PBUFJ+MdVsvSwtRD3NcERBjekLKIf0NRiSQQXwOnrnn7vlTIhGwE
Z3NuHLCUbjqMguVeXIeVduo9HSuJbmJCaEym7BcZPzvle1eTZqlCQidh+kxqzIM+9qwK0n8XhFbU
nIO9yIEB68Z8iGtSr36tJXfbxRk54LQ3MrWrR75ZJfIB3Kl3iDbN9TtLoVfzBzxZAtiW6/RTQBMY
8LSS9a/oJDyNLn3FC3xBDyDo8ZD8fCCKSpSY1X2eTESpJKMQJZ0PpS18vE9ruN0L4uJvGEbNwuMg
EOEfjxuCV/+cfWIC182pkRuTmtVfBEN4QIOL50VMwWpzyTuCqazZ5PuS+qn5+CPmKeDMY+36hNJt
ZbjH5odZEPb+Djjs3zXHdyQgUQpO/32IUAvZDTqjOHt1khWnIZGacXzJOhj5bG4i7BBKXZ9ypHux
eHnzDeyYmIsPNRw+QWT7UGMB6zndxBf/0BQtouODU+Ihu6LRUyy0JrwcygsE1WGioO9UPdwADSyZ
K39/IiSDfPiaVoSyrgYoX7mnrD127IwB7TtahRzaeUsG0UvNjchUTq1slm7ho+nDZGy4U/l2puyD
DI4mcDvC/NsniTzQsxAfswvg76oupKbbR6yi2ktgUhx4VZg0Wf9QD6i8cWzWoHFg0LhHewP1SVsU
SfOM4UDNEmd209DdnMsNiQhmv/GNzcHGElpk2Gjg88Xaqq+BvF50nZERgUxBeg6hzpo92W/aBNqN
zwprVQeQiTy3otwmR/xqo1q7ClCow2UDFmcNb0hKjGO3qu5CApTi+BycKyasnUz5mTT+RM/xbwAU
Eq8fU+7tZOmxSig0cUXwDIuZi+OMK8irY0Ly9FvBKlnQTwBGJaZ+E+Z5rE/n/AfUEGrtUbkW2r9V
newy5BDUeP2HAJSofP8LR+d1iJDy44J7pGYa58E25eKHBdbj1L9gXxGuppNOO3vHlShMN2YOmBk7
5QIPm+FCXHgPqevB5BbW8hYsLPe7/CRE+n1TPfn2WANYgnNRhU1gTp6WUIb/1mTVwyV1/XD4iVJa
OP2NLRJRpdIqJ3JnekQ+JUANldKaEcTmMebp/DWGZzNt5cVOFJA/0KkUgozi/UK98374dPn5hA5p
IIb9qlfBdUQpqWEoESMq15xw1YglIZ8Cvthoja+YkvgVXuPLhaqRs0wG6MJXgXzI2ZWc9KJJ26gN
YMv67O+RheXKDmCk0/A0M5quDMfqDLppjuROiZZ0XFCq3Su6SK7EIURtdEMG+1BaS3u/nfkQadkb
ENQTLlnniS5bha9TdJRhNkyzKrWODxXzB79qqC5muqAk4S+czYEQofMcKJwJjBxpaNmsDxKP59vZ
shBKyVGoOwUs49I1GMV3vUo83fK7xVYdDz0Oa89p0vhw777gORdUJ3hmtEN6LzHIpGzqYh4a68ZV
oGA6lTUdvScdDm9HPOxgdcDJRHA473FkDW4qvVdwp8XGBAlAh2rgvJy5sxmICCVfqkJwrzxlA7VR
4uB58yGwVOeiyOwlx2pIPPautPgppEARf/2BepJQEsW03DuWhtI8R+htxgboLpkDGT42rPWpYiLE
CGIPeRFJ98bOpBtHKorQ9ckgPs7BXyR/O0It3o8WcJDl8/UH92fkLrk0ZK3LROJA/MLTvbTxA5IO
gICRshfB1nJNDdRAHSmt4jbQub2djXtxkaRi4Sub2E/TN0rCbIEYRAA8h2/rhadXjrvc3LnD78l2
t6iP8c0+xDGuKNm8BsDyEE2lU0MiYrFsgJoY4NbjacZaXusseZboV4qaj6iXphJ6kZhyXXiKGdsa
qPszpT5LMcQ8rXlztESumDRxQPzkIm1wv+PRyAdEMnt8eWl7vqPBYCUWAHdRyUnJ656xONFqXPua
ybmtOVVF0jTCxKGfdBtzExK3bra/uJ106trwd/643PESoEJgIhiBXt9FeL8bD4NlOo0KI35kSO42
mQ3ZjkndPw8c7I+XeQ2z5qSaeOirStlcjANXwNC5g9s/GMNlNxKaaYwIvojgTQAAWAzIN4EW+C5q
Bz5a6rqZ7nWzYScpOcXmfYjAfRDfFNcPHWVRPXOXmfI36klLzpSqE3p3yFPa2Oc9nrh3JR+CHwxq
DfSMYFyyTN+2CeQ7tAO7shsGpQmSdg7P5/WFZ/oLRUFojTTDFx1Eq2VnXP6BgSYxLsKVz9bSoWEa
4+27VC5EjaFJP99soycGFRKVlgM/ca2nJLcIpksE5dpNjzdCvox+wkRONn1e+OJySdKc8IpjKQN5
2QY10w5RzPLL1RMFNQzjJMD7MpMJ2STk/aSRtz5xQe9SdiJ/+lhxY2q9PMsfrlizIWI8D7TKM+JD
HnyFRmnFtiKNVck1brSk97W60yJoFsthROX1KGHC0ReDRqcXE8hVvbQ8SOk3VtpzsVuvjhi8zffw
re/hBpysAXtQ/i7qYn1Av76C3R59Eaa52rHvKxnyQi/QHnw3KBQPasYo/ZqQMudpb/CSXm5Z+eM9
ptZvKuATAGwTD6Uvje8f6AVpYVeyCaupGQV1P9wepZS2DR69pJtP6SVP38NQEGhNsL6QgPiCz+jg
iUVtOTiNrfxm08DJ+NgHi4F0aOmMZ30fjYcQUHq9I8pHmiSVOXVcK7sMe2gxU+2JAgjufWsCATuD
YBTGvb+qQ7pG8o7iqEsP9fpYhxDOOgaUCAULOMd00nYXaTWy6ioYNG81jLxlWZJBc5twdQxZ0fO9
R26VvioWWpBKuhyI/uHDZA4Fh3994W2uKiQumky9uvmtID+aJkzND7QEF8+jJT1BlROwEPT2iQk4
Lju4mInLrEd7G886WAag5oIAwvr8dJlOH1uiWakuw1Cu6/nxArn4gAh9InDFwfTFuKzjo6Y6FY5k
LAo0y6KXLL6YpIc7jyT8QnXMiCNXgPEglkiJjzbSppk8Dte83Ut1oFm1xNXDrC0om3bm3pHVUeBC
1eSQLKFRVZxi2eV0yzT7gNPhmfo3u5wBU9C7e26DUGsHoMKsTr4n1sp1XER7eMeArN1vCvrKC3Qd
6Z1KnJORM7/qydXpySpL59I0tHLlYWC0ayYgoFpMh1RqnM4+EMExAd/bm9d66+KL2ZQJ3w6LTDjB
lC0GZQNekyHFPjM7Gz2OguGuTLHBfXnHw27OMNZfDtMbKpSkDMJNvrn0vBsuKYvsOtzHP5FdTD2J
p8L0c1nZ/ZAqjTZuqOhsHLqszutUkitxVZDxfN7Ms0rTpWgc2WpcnvNp3bcF4qwdEb3vguwBpx1N
MGU41wlFjiS1ek9ZLp4o9FPo+TI/G5tEcxsZ8BKulqvBzBGAs9sVJgbi2fKSYLB1bq5HBexlKfHW
ear9tyRMS/yuNhJH3JMVUjSgIuvTBQaSXoFVyWCxhTIFyhuLii2XXKZadpV3tMu3jl+Va/lm/xU1
ZoJqZwoEhgTEl6hdrWgsl0HYOPfbr2RYMqlmRG852FfMzlBIclzzWAYZ5YqmeGkW0RSlR+8b/hlh
oxzN9NZ1O+R+8OiPkezmiUyr21lEix4bPDeUQkadkfNXlyWpRTcPkhHL3JPQTZlU5iSumHjiXus8
YNJkEadmElu56meUSOOEYvo2HeuFGI4yA0SGpGPQ+fd7bYJJaQROc4W5kQyYrELrtNMRIJ4Nm9Em
m5SDlRbQ/dWTrzxxck7wp+GTKYW5wB7q9vycfQYxUvpLHkzL3DdduCXbpMaZO95OcOIi2H++0K9s
2E20OwWRQKXqr13YCsAixA3fXKRlxtN6fZA24Fy3iLmkCS1/dw7T2iXzGp8NVaM24QDz3yLebpHr
6XIarRYEryQXMO50VOAzOVGdjBJdumAhPu9GFCxfwECPU7qwtDv3aWSZZWFIU1AlE784+0oi5wzH
ADtpf5p8OBnP96zcOC4XD0+ZnbSnfwAmIzkCRWQD1BX/vnYgcgjDzG2SiH7QgDa05S1+0DngjPEz
IU6WuQXaum4U9FaE8KQKInl+jhnHYCzGKtseWVKtEL/TINYvEUTl7eM3Qiel91gB7z7ImSVHd4IM
h41iX3BY0P7peWeOaYtCs/IEI7t+CdBDXJj0budM/FwfNs/AHWThunXQIxmL1C2cfcfRiELfzPi7
Dyw72RJkODFGlVNvsAdJg4bd4CPUOf/u5N4jUjRZpRC17cNyFIvD/J+Gan2wG0nzb9+pYYJSHKab
8CfBFrUEdjzgckf687r72r9Y5WHEKRz1XIArUPU00MED18EDzO2e2DE2rZyyDWrf5Q8gF7BqoUd6
QbZbMq6VsI+wwu1+aZzRDV0ppHtJ55W9b+pQwRl5bpjVmEw6cVggtaDpyIswHWVA2KgHnFckGvk6
B9s1ax4GiNV9PDYe6GYRps5GaKPPAgWifd6y0rkOYtMLSlQlJQmtvSnUifAEJtV+KdXJ0C40XQFX
toFA3B71oK7TgP+XpJ4ZtS46/3fmVNDO2A+t8giNweST8jDpACRSiwziFKdSt/bpaRX+2hwBRRFR
rvbvSpJ5TwkxCdTBB0kAcxxJ5ctM/bXG+roKP/kXXhhdOcSTUGX/j2nFpT86Ag0WvyLJDm/jx4rR
HNzPCqWnzu+xJWqS+MB7kjjMif2Mi2hhoIck7O/aIdUH1EoJ6cvzff5Y75C8HdAPHA1ZrEGVadOx
fSCM5d93R6ku7sliPriKFmDmXBTAjROyUHO/3LQpQ20dpl/4C3HeTWl/4NQdcJImKCnYuTnXRuSj
f7UEQXIwh9p7283iV78peYcyoO7MSN6VB2CsS1ki25y72h8uxRmWUXdpcTZjPJRZpnI/BtVwqgiF
hFr3xylLmRP7zskby8bdhswq3U9Ph6LEX0ZR1+y22ZBkuDU24iiT9Tq9eN9v+46/mQKVGR7L+X/b
l20hGlKlvR/foR076sYX4wXbdaqQWm9Mo2W4QaTGgeZRQuDRst3ZsIRLA1kU1KTUXcA/25wblBkd
+eUcVNacqPuJfbsGiGS2DeVUPu+Ex3pA3dX11II5ujEM3VUCa3mt0OvSiWWfcnukDeRWUm3AQ9JI
0wIKb363E2Oj3SDHEU852fJnTJ8PoNQa+9f40kb++5Vh5jjeZRVHJWEyCwMuelOJ3wXCfs697GRa
kqlgfBYGoFL01+c3QizVLkNpjhy3w+RwyQ0q6nApVsngbDyEGhqcvHmaT41iqKZjhqV7gA9HMQCH
N6y56yp3cnUzWfZgGDXOIcUpcp8VtKgoR34fxQ0DColgs1Xcob6bXDXQlOnK7KZAUbbghX4aagLM
cRukF59S07J/yIlCWpT8zQGHLhTZwWSFIMFcdF4ZI3bMjCoW7BpvbYHBxcKBlHKwjaCjMQnfWWSZ
VYYLRwpA1FJxRkKuC9m+PFHBRZGaxn7deKpSFfvHJLSEvQuMgAn7ZSGmZCnQ6OOQs3ldCOSlN60B
5R26vNjQbHVJ9H9gjkkmdJvlLBOHUaqsu09ofjxoJ2BL04DahOmwmh+x937K9Q6hvEfsSdYhz+WC
1AAeg3rllMGM8ht2FXqz8FbBtGyVkYLX9V+BkEF2t/QIzirtRUKIyrhmYmYeSpm04w3WeEmLWUUq
1i6MKJlxNGVhSgztGBfiYlDGMrrmYNRdSW6WOybTAbfph6t9VMtAFYVpWrwHbPOddyIr4kTLBGFd
D9TWUUQ7FdunhROOX5dCuDqZ69Iq4c42TOWhB3EIU00uoaLUvN2GO4dxnVEUeNxoc8il6g8vC1I7
SEQ82df9Iqv2A5tbiioEGDkOagzH7zjVqrXuV8aJe0MmqnTqjIWBkCqDiWID0ncMP0fe5ks0MeSa
Kocz58pUWuSQajx+ki1CRBVyrkhZqQKj3ebgQdvqJAg5RhoAU65rdE6QSiVcEKbG83+wJ9J2czfU
T5jtXGc6e5LxrW4QYzQ6djUVMDqqK7lllwTBW+ehZzqLsMH2DxYq8BcgVR4N+lr+d1tpNXZGNRiq
bO8djdTH6YmdtvxgFSgTwqLzJTR4RRa3IWTcrpakPjzfXXZ5dbrQ4FYve1YrHlco673+k7p4dam5
HcJx0nIvBlHg46xFjQQdhYJfahbC53nWgcCOCiXlWnceS+ddzu70+RuPCLcdbH5cxzhHuXeH7QEP
Vmiz/ZEVUP9tWxSH6CWNeix2fQVjgQA9q44SlTc4cnVWJvipvUdOstyEKygF9nJTy3lafpXp/ERM
eXE3qwZw+A/v6lVYeOw0rNaxWpM/22FeYfJASQHtudmxN8f1FXgMbaCaqSkIKM+jE5BtqnF+EvJA
L58QwYsq2k8pMZY4BEYJ1innHmRjCuTWY5QBBhNgKeQSMkwb4YjPK/ZaD/WPHIeraVLrIzxNqfao
IFeSBwQhTGnsyC1NZThp3ZFvUB1Ih5FDhV/PYZn+fDxmr9b25N1Udn8zxLWo0owsV6iINXxDREV0
UrQOja5IEOzsUcODJqzxS4EJClqyT5AkjtLoytQ1EHDOvdLklHe0k+HPH0tXSMUwmGy9lR/11+f7
PN5Lz/Kni+TzzT2yDQBEYLZwFI0cTLSPoujX7UbOwRbHrwEDjmotpUzIsJeC3PqPRXBNGHe8zP2o
I5yU6ddPU5R3YmihCMT83iyl9SQ39LGQU2spq5TVjqauwCVjHkem8B3jlXxicf2K8rv5UdOek4pF
+hf7fD6G4h0gYcUEDbu/oHpXVuEQKLJ4jFsLNv34qqngsKh8A65Om1hbPqXVJoXG6fZxzMt6bu9b
LHvN+3HI+5bnRixPFLRKr15kCYGvZBGsFYxQib+HBnvEcjUF6zIVKYy7Kgs9pOz+4SOZGrmMAhaH
IjKhX+MYK1sfxH0hAo/wBQPYwAwcUmxwDhSYpJ/6tuOlaAWUzzZPU4hUTchdHQBIi8KkahS2/qZN
JyutFF03hi01m+R8ckhTSZcmii+0w8VO4v5aq7vYHk/cWbGr7mw9rHCAgwq+Z/3EN4lT8JF9OOpN
zx5RRz1TPBOb4+ggu1zqJv/UFPKhhfgysHy90bQ75jja4Rhqqhiv/vA4a+vk6BByNV7KVHcpqtv8
sPk8O/fDaqOcqs9E35BzF0bIV4XITvw0yaBCBykMkm8LQyxsLHG7463qsrBEU8Pa5kx7yDeKz96r
B473MOF+RzuXAkhsTRzbI/xGrBTzh/PcQXMr/ymcCj36qSP2gSN6OGzjkgeIn8hSLCLZ75gA30kw
U4VN5+aM5gsKf4bZVXKPnBc1FKytObslaprLITccm2e/hgKnNXyyufVGm766EHVjrJ5V7rjGcd1p
KBSxS4cU8sc955c7kiewGjdGzr74DXNcJ3w8dGxvxcaoOPsF+eECCVh6olQg8Bi5Q83TO/3gh/VM
fQyrZoYg2z/153SRFHDXAusGjPV0+PCPHOlW/zrPo/5SHuoCxoKGS/f+4iSVvjKyoSadPJcyXawH
/x0gGMY/mNSjJXETNkFbCRUA0sWpCe5pmJEFcMl4CVDHXyI3IMEFRgrxJWj3MBhheuICVtuN0Luy
X87Bvnk4PPw+GIKXNEpuX0FmwxJ8BihhzvAvuC8XgaVWih8yAFjV5QLRHLybz0vAG8iMwVB8lK+N
xarjfKR5LwAsUx/94nFG36j8dodMxvNE5z7FTeHW5xR/OiRMqsOpeUOIC3x1tbA7zjVm2MWOk/fZ
xa8PvVccId/GSVGu4+e7tatUEYwKDLlNO2gvyyGsbaZJrvCqGEs6+lzdtgvmNyDEJYaVR9jvceAc
b3C7XLMcF/yUfbHpwBgOfW1BXd5YGAyc1wq3JDLsSNEyA1It9uINRmKDZZ+NYPBZisBXT6HqqwYO
mRiJFJ3f4G7Dc6NlOPzHZDMnYgTpEZ05vqUkS5h+zuWIbi6LekkBqOv7+G1EzOO8LFe/JTv/uvan
uAYlKsSmjZnFxantWR0/JEFo4Q00baI/V/dUx0/NFipJUp3pcARyD56I1rOpODdGrG99Xx1+l2SW
qHuaI7/UmSNM0nlvy5bN6Q1kam0dlqJ9TLGOcVORVUP2181RHLYKADEv6yDbp+So/1apwVt1xtSe
8+2C9Htg6rR/Nx6e1Xuy/Bru5OxUYnYMqpkG4txq3yuXHT52fC3FWJW1TMvshCzkypgBFyCigEJo
aSPbpN/GUn5ssj//t1pxJSWrvCDXhhV+21NqHPaEfSZCYZ5V421En/7MkW0xb7+LDzJkw/mjCGgr
if0p+4wV9AVn5Ez+JCXGp+IRL3RPJ20uJYK2F8Np/vCXhuiW/3OlAVgVYglsHTJywrq/rcFv01br
exqJe6R+EmbN2EYlE4P0bukZ1nKvyE678mJMKkXHOOeK+AkwoopvG+On8FQWpOdwPJdkOx/a2RiH
EEqr8JY9eS12jpZHKGiMhqiBlc6Wy2NeIqbBGc2e0tI3xM759eCEzINj/deDi/1Qur9untJ7WePg
1kPvSwNq3/gLvoTC6D+EIPEdXdXLudjuYNp06TMP7JP6P+IMFQh4YOrsTxyJ4vZZt/DhdxelYRXU
iaBThQdN7yRbYIf3dWrIqEUtBNC6vwXAnpv3Ro1RIOP9QODx3Ojcjv9JRayU5Q2Yy2dkFloBhtab
/uN6bYDt8dUCOzKjTFCjxTnIz8qr5YerO8q292tm0OhGu9Aq2KdIHq/yWVFjmwWHDSpgNWMDZv1e
zX3Pp0U6a0puqy4R96zV7eO3efv0Dn4b9YpYRPPSRbYYZFvleBR7QDHh964BLXOT4DR0WSBd1SEN
0l4lxvmL2Y50Mi6mCzG+D0juSunun2Qig93f4MCGYjhpUbGLQXnQPXsgQiGxiiCENJQy/AoOxVMy
1pGkS4OEEr3TD5J1MmlANDD5/qNLXaHaABQgmfOdxS1kIy4t9HRNE/JpUmhOgoCgr/j0jU5ca8aX
VMk2BIoE2r34FJgEuHY3hxnzkKcSFKjNzuSxCEmstf8dOIIu2KLr0DBsQCc5oDJHAJ7FLURrmZ4n
eOPGr6qr5m9Dc8UzSPpdAhk33lSMS0N13Hph6E+TJCYcQ0jxmrWWsa9Uf7C+tLDD0bCOpr2Z32SF
YQxd2SegWUHyaFmVKTOUA39pRx73hj7hoLzTCDOTGAm58bqX4ayyZ5BCvvSrXs3oNqwBRNeBaYVK
eCBXrsG5NwLimjNgyWcxAZdUSgZPkIxe00AC3VdIQc2IAjVeweuT+Ix7Ox5gjmuoNzwuexdJfUtZ
smlfpJpuuLvIqjI2ZVrkUHpnU3B+bVGwHiAHqX2aW1uFdHQ16yPHZEpvukXGPxdmSQJWAxatinKM
EQyn43Eev+Not5xPNGVbqSbJGif/McotZH8hXCkNR4aLStpzVO1OYA5BddS4WPL0MhX3JTjYnf9C
ATI3SBzQlZQY9pu7aIRilLgRrKkecMSiQYqy9Sbi4ajXyNzNlcBSbDvIkfJKG1zzqfuGZ6vRjDRh
zVHheRZvB520SXLcpYoX2eRXtgLg1j12K7J8aP/NcbCFq1AAnbFI5iFPrkwgoVPDV8POg9NP535o
EPIQwnYA6IQXifO9D0EuoPTBpfz28rR1sgr3CF6EsoZWJHyCS3pUvdQnCzID6cxEO6dSlgVu4Ze0
tQAHWmfjOIulXceCYtn2phkVKLZNkHqugWWIkbmuk2mj7w7nPndEZan3kKE+TB9O/XXtXUlMU4Ne
aBKr6/QhtOddrsO/s7X9AhOqr46h89FLUxGOWbPA3MzuTn9pfgRz5alcDArFF0AKCDYw5dxIxyBT
0597TkIrWSdAt05L0TZH8u5/1hGyKo1APOgzN2495I94XChTplMXnWwcvNuKmTuoXUDt2GY30YA4
trB2O5D7WxQeHNKJQHw8XJvK2OekSh9b+AkBMSup/5VPw5c/x1u1QAD4jlJaqQYeYvXgflHBk6rt
jL//cedbHWtZ5FK30/Vgx8WdaeKZ0nVG6Z0UnwXBr3baGpBoEfNDdhzYiIiAs2WoS1z8Gs9HjHSz
m7VHjq6GJsXNhKX+nKOGLZzfh7LSFTZEz//TTCmoH8KWpz403Qq7UcH/b46k0du9PBMqdw/eRkdi
jd0mKHmftX9BJklwX43j80rG62pfN1MBS0fA3eZgF0Q5JmoylN6UQMNN6cMfOdimaFwYiwjE8B7l
SjnJmF1FOzM+le9Zmyz+R2CkFHQArA1nMko1nYfP3EnQAcJGq6KORomISmXSE5KrwR43262K44Fc
bZ0EQCNEVFSdMbJB7XnEnGc2Y+hcESFVqfvipMr5ZydOPDMWBRtvh/z1O2G8fxDl9xq8H/1cdWao
oQ65jshqe1IuWjDLfwdTQrjbgIj3R4/3w+uFHycpOkySBp235LD18x8ZjKbwJrJC7xogVC0CAI/8
PeQwCf6H7Q3hcLHP3kVStfn/c4ok67NwhTqdONdDQXXnm6keDsu0XnAUCaFxpK3X9OTiVVoLcjJ1
YY2F/QGP8B/d08+BTapBEaW1IznLi/MJx8bqPG90+tVIYmckW/mbVKdWNWLCkmT7ZK2/ySv7ljC3
yRbVaDHGarE59jGzGEOLUqaefQk6mJnMrQzu4QsK6+fEgdUcRHSY9EejLEQqkI9VGnbxU+ONPVJa
J7IW2CF73X6L1EXd2kaMEAeMnyRqE/7sMll96PnGrN1ut6vMm8qJJPyjWnlUuRD5hhxVgoFxvD5Z
RHRGWVrp7YDER+iYfQJqqjHL1AoQue0yWOUlujlbTuKgJVTaqFSLSG0n3mf/FH86vQUvB+iZCpjQ
YStw1te8pZTMGL+gMlrJtJyJsNVYmYg7D+N2xVy1YpipvWgMFte9g4P81FtX4blsqCiL5CUNaIrh
7C8S0WpK91l7ATZxCKzzsRq0Mpkwb0N+e8lpInhqCxpjvYTVjXIJjcEif/27XCF1X98i8z/nwzWh
24xkJlQkv9wn0BlNRz4sjBoUKCvYjJP5yPNXkc+iBHUexCwaGwHGquKtJwCLWsNOcrdOFoS3oV5H
hVga3uxsY9O5Bu7/cTWB8I3yPTGOx0t1PYeeLEvqQrEhvsVXnBleGmTb1htFrRsXi8nr6Mtcx/jT
dLpOhFwhQY6lQnErlqnJM/UnuJ16NNyX5tzw4yy2ZL4YpJvMkvZmTuO2ZExRaixV1pukNIkc0RM+
HAPymuzE3WxZqZNdX9+pMRC5V9eEBPqkmgLcZiTitO4+ejNtY18U0kK8SVfNCvpCKidFO7xo3KZm
4A+7ZUujhPjgOI+fzbv0IovIYQE6vzPoGgD+YIYSEOLPM9htciBr2HVrBZM+zozZ0le3ZePYUt3v
GLcfl/0Rh40ihCrYR78PDVNGETy+6Euf75/kKUd5Ft268FkYX12gDbUAVk5Vt0zJrixBsoKc8q3B
Wn054nXe1repG8dhcxwMqfdvWoAgcOrEmDczP4ztjyYzB7T8NZ9YXPLHsKDD1hQxHmpx8h1MypJQ
yVv7UKCiQylupKlDE2rTQ9btPBbLK5Jfl/WHNg+ovLtsGmrPoqVwdqC5FnIYmmryc/Ci8l6NiFyS
gYYVtkAWYGQGSx+sDN/+ZgzOdOVZyQfnk0H9BAKYRACad1q+rMwxw9rvwgDcIZUx3LjLSUGwgHTm
nTiRf21v0xYNvd42PbrEjkI5SZ69U9hDwjqyIuE2/epERXpVPryVO85a7m5WftW8xRCU2W7XrKFO
A0LvWBzvgpajzyBB5ZUCHFEu7Ii9W+s9a6DUDzHpYH1KZuIfudPlpREfUQU6oJGRs9n0g2+0EADf
6Zt8hgOAZvUMJecM5XUsBkZHTKpDxj+hQU5IRdM9m0G7R0M+dj90AAtNOJ2OYgm23lFCehVAvHhd
XzWF4fPSORnA9aMZx6FMaen/kCM6hqlBAbug0y2TVOc0EIArV5wa8HqyJ7NQkTXeWPrNWedXUdjH
rHOrK3qiGq2hOQDX+8FpMwA29H7K/0UK0bxOvmt4OFniPNlAiDn+ExScrcn5rY8u3eYX6lXOXqaz
loFJENU4hR8pLHowvHyzLuhiTAXnMJkzPLACsNewp2ydDTno9hmlfcAfuE8OQ3DlqXbsIg5LO4uo
DIvdNk0gYfdUvtAWYqNPE6owmHQxjz9X91I50FSE+e0y8UscgD1xSWqnU5kVpuvialD52KNSoEO+
6ze6xhJuCVmlhOhkCzvOW3wnMK0YWKH5arPcRQmLo806XEOS1/lz4NlSUkCD+PRyMl0lw8R/RCYO
v81jX+MjhgYO0HXG5sy0RSFoCsjvefbeRwrffqa1Oz62wvkKMm93uH9U2aEgZ+3hF593pS4DhPr4
faD1M7IvOsU/4tJnj5j3WxiK05GrzekQPCIcNoLudsEV1bxDD07qiHyIlRaZtGiNZVui/1YbIrb3
NHZoNTAGNXiYPiGmVimLvP1f3FtbbgfMh+979e+0NQYAv9uxG8G7YeNnYygA4krNNgADOs/12Xg3
u31GjTHBbEGYAwk/VTVsDJCyLQEAgsuR57OguilGZ2PDalZzmRnJIHQk6RA9yf9m/CZV8dbekABG
lCHkwn/oOVtQF4uAikqRiTFelb+Ccipt6UdJXYFzI9VuZzAwwLp2ZszDkVa1GHGSlalrguMQ6L9g
zArxeJ1PggXiRJTa1aDoygpHkUGwJIb97FA6c9//JxVcEampumUCMsd6jnxvRFGRtThTwoVUMYQf
SsBb934Cw0E/bGvV2UQ+GnCRH4Lfk2BB7EFEtfwgKjMGhntkl+VjBJnD0H+svU1zYH/2C4hHWJ/u
ejjFOVfE5APEqJStIyHTWYzuRs+/S0JuXJQHH/lJAIL/HAjYiBxLNBMvC8LnG25tB/EGyKSDR6mH
FnA+I/r/OTXjtSoxUYQimP7kQojDx5rQEATLeCFAr+7UqB8HVD/iAa4hgLKlfXoyM22UCTs7Jl6F
JeVk+s5d9M3rPI1a64AWEbB+u9uxR0tVUdZmP+YHDq+ieSU4BrJSRFK8PO9XNlvWAumAQ0A3AAgG
w4ucCAZTr9J+IoqjMXtCCWFnBWvY5Y1zNBc3uDte7F6eXwRR8bYLK8/Mz8wk7afSOIlNFk735xkF
XxG2eSL/80Om3hShHuChaY75Azaa4/fXbBA9TNb/s9DP77bktRXTic/U4l6+6HZ/ujAVY+60pC5u
D7L0Yw9m9YCAum9mkinPJ+RemYzXIoX2zwUD5oVu1Pra4/JfiIoZDcSzOC97/uDLQVlwSsxhB6eR
rbSLFEubX9XMU32rJS/3To1Y8P62uE8Zxs62FsV+zzr4VTp9IYj+RnHU1vWPbQXhwfY4+OsPrLMd
BwvBPXoh4eX8hW+6/iRCoYiehgcJh3MgO9xwonfXQgtmKTAIKCoxR2CF0uqn2dZfb3p02yMmxjt/
L3T2R6XE3YqEjMiHBJViZgdYIZWjnrsLfA4POdJgV6A1b38wLG6H3FrZzFXv1M3DIityKfBq+HU6
e961G5Z/1N9UbUkpmaxTf7uuqxssmEqFFLWvIFvq8HnzqDSlDX3XAev1N+BMjzSz2YuhI1p//IVG
k0E/1rnICagHh55lyHZ2tmmq7AFVj+kJ+XBg36D4hw8JngbVmQhCVZgMFvCjcHg6Qieb32zpA/sk
8GkDCCoBQzkjuS2loCNhTtTGB1GZhGEBvBG0/oePlF4bidyKhxME+8Hy4Vkti8oiq8d0P+MTiGt5
OnZ6HtkVSJnXQXzhWH0svE8mgr84QQIoOELVC2lQv4YjDutiYNXiEjuN1qwVSYx49eIx8xOlKxX5
M5ACRXVPLcCeH6w101g7019FoFuElo2SdsiFUGCWhOPMoed7yv5n9MvOy9ANtbHXnB68DYD5LKQy
QMkUf031FnIdaIim5M6bfdGd0bIfbBPYCejRItVy5jy0XrcD6LVJrNV5WdWLU2sl6vRddfRUNxLp
XbPFBsa1bOrhza55jhaNTdljyhFfJmJ+UtGjhupNG9y3dotsHS6iELbxngBbgx/K0Z75E5vzym6m
ZEGrNBP4f2PCmUDZgABJNjarU1gaakzkWrbcX2Yg8APbd50Coh0z
`pragma protect end_protected
