`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C0DRmsC282LWzIFXIJ7hlMJHvzpI2dGTdrwEMNozVYJ2oAcbbHjg01jG1Kg+6Uk8
5VPFaGc4pIjDf5jHCqEzO3ChBPINNTKWeeh/QSaAlaLW9uOGvZDNoEr15YXMCxJP
aCWSG9spMFDDIotOpITJ1ErrrSAJ93IywRooj1hSCEc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
dS4fSynd0Q18odj66kNWzu4hc8yg3xr5plCkYL4vtxFf0FXWi85954YWFZah3Mdf
2OPvbiH2romjsN2vzQ1wItHaVLxyGwCp8xv+wTjncv4R6h7dZf36qxR9ujqzsWs5
38NuYPOCxa69UOyaOrYf8T5sTfamOOC8dBJ2DsCPj+10+JR1J9noNcnIV6dRc678
V8z/CYEMDf6ulA3999m3MbkB7bov6YDjyvhcib/oju0SS1xQujW+sS4p1VtZJpxn
aBXWFIMffiSjUUcCevav4Am12WzjNXWCOgQG2LWP1yYnVfvNlFpwy5yOU2JOhJqR
LZqCsqiEsQ5Sn8nS03yfCYRGqA5tC8glV8+cdeitQVSyVq9xPkmcX6QA6BzCcaVC
2o7r2WGr83EB38zRDRExX5lHUay7TYS5dk5GndjXvsnnx3mBzkR0wu2EyDKsobcy
3JT/GZkbtNb+MYj7xCVJOJt6Lyf3viYhFqGmcmaB5s8ULYLGpyJoT0K8D8Ysa5zn
K4dUec9Bw3hG37ibPuibDWW8gmh6YRcPg4X+ol2j5VLI1Z/BVr/XuhEb3yihCBEx
OHKaatYgQlfab1IB3rUGHyRUuLe42qwlpIvSOuBHDQZKwaMl2lkeX7K8Xy7GDNpz
E1rsLyTLo09Kfl669/wnxJ95N2KjuhixX7HwYZ8noXJ6T9RLsQcX/dkvpgiITL3M
x5BrJYL4k6zBJLVi8YAZHbeF2MkfyKXqs18xNcpEh7jw2rEvn4GXfGHzuGgDTje9
rEA1valjEiwdRbV29st/sBh+/fmS4815gxeTsp+goivnOoaR9JSSXYZx8PvYXZ6r
EWjPonxNJkX/gaoh0XFCjZLFfWpBOuqsO6dSGdD8IzUMN4HUL+c5zVQZuaNs/rNk
C4Kl4PtZkKeHm5WbYBxJv56dRkM8oDpBu/vb2h6PT4sjNq6ZCO+pdhGhtGxyINxU
pCrPALZ8SDqiC373y9T+CXPsIizGCMk1G//HJff+lFDcbsw6Ir6hhmURQFMuDRw4
+yRntoqEDCtjgxHdTQ96llStF0CIMBOo6XBgo7mtBMpWFzYj1X8pAc4ZanyyHQaA
02fYNYChWV7diIEswB7/iY/fwJg8jioPBXrQqDbmVMKOd7wUOIYJbfzOBth3FIGq
rowh70wp/UPWMoJDyfdFiqw9hGTuqOpRIgn30QYJraI7dPNZmGAbh8vDXM0GklKX
gaEMc3lOeBTNcvEDPpRVri65IVwdRZ2amjlD0TnrKj0N1Z1T9GT9fXlVDmqP69lC
czxMOaijVAA49gcsa3ilCo122cWkUVcjSo4ZzcawH6qK7Z+lNt65d84FISGhWbwJ
/5TH+LzU9ZY8dv1cHv8pxf5qi8ww9IQTIewBH5/AeUkiMGRcP0Qc6Q6Kgsdl+Z6s
7odioZtburudqPr0lduXi5rW+WsyYQnPqvp5R3279id5E7DiXMxOHl+OJpajJxSC
ykKILagstqElRxp3AQE11ITA5rlxqXG/a6oB9N3qAB/qOsxB4VteMd4XDfbPc/UH
KKljtQKLfxHWY0bqR3RRAgEeQM52zpH+FbBwgIEZVergXJXdlsu70lSrRakurDB9
d1A+R1QbGSIOAp7s9U4rXVmja0kENPqDqDyELY9MgQxkYQMrIyr7EtiFCMjfZBDL
zWki443RvYBzgyYrChO2i9EBzymHXY2HmDLB5E2skcAO829KUrpLJPMPbRYsmVUB
Yk3f3xv1KEFHSuemYu5OxpHoc7snufOzYcQXogxdTK/e+MGpLTtfY1wfuDj3vkzc
zD1NMuTSVHQYd6+RhqlBltVeXDHIDdc4lol90ETZpvyvM77c1g7xVePjtcljD9Pq
CqKUaAgPxBITNL3AYaUutmzl5BJe5/8eEBh1MQu23vhB3F+ldM47tZhRDIZqrNkt
cY/g0Uw9LtsMRoyKQZ+AyJ6H49QrS8DVA35yrIXkzkwPDJSZESRCYdirQ4rSFARD
v16ShR6ISzpZRW23iz6UkU8CDdWW3kMQ/JHBNfNMmHOTAdKm5h2eXYGc1dUKa0A4
nRyud14ZPL0ou+EH6CsuMc3nlLlfrUabfXRr3p6vH8F148h7Q8shnMvgmw5Sqy3z
jhYy/+tyhx0Twlz8JP/TVOWoafRZ/4Xt8wrj4XQ1f5nCD71463T8/L3m2AmiAu1k
+5/ykTt+WIMpzdmiXLFeA8atrBvvDp6ABu0pMO//EyRP7J7WbV0zxi3SPvOYac1s
o+mMhdGUTV0+xpmrrleHvZjUe1/gdU6MGdAhUdDZZwG4DZvbLMQz3igsqlkFPayG
1R6ScOH3vLT0WM0gx/oHtt8/o2VeutnOSAflcakPW+hvwi4r2lq7p23J0i8IPiPl
p/Y29hj7HXr3wS8wMb9hIH57/lRd55UcT9iX1ni9Z9R9fPORQtpoEjMnNCw2dGAx
UyOrzPeL8N6J5Cga6+IrYRM7ExRUVBwST7E1ieYI3alOgeR99R5OypwhdHOHk5+3
ZGN7UQ24hl7n4AUoXDF/C0IcINtN07b9CWE6pYIxMIeGndnSvrpe9twORJaOoq/D
GyKNdEx7Pf0O0Nm2lSEezKXUSN0WtVrhJsnqmunrSmcBInko83knSvs6drO0IPSI
VqMZnq9Deyt+UvSwy02jVOcbcD6vjHjam9K/B3E1qvlabaVfSl4/14hN+k+8TXHS
4KQ9dYKSg1lEJ5eDIH5B4Mw6xN0JVl2NUcS5H+uLLsGugaLi7sEqNgucbZJfk8O9
+UX7rKM+mKbKTxkHA41iJfxoMvy7jepK4MdW0nqqQCqoLVWHKtg+WOVdx9FNOUM0
t84TsFSy0wbfVZTc8o6VDDSOIvTTKgIRPs+EJfLDf/oaWya/XZymZjox6tl3O8Hq
GoIbrus4Uqk7WRtWp3NB3EFuNquIvxG/meYs6gzzQo/iIIU2YU6zcWZjAiWTH8Bg
Q6dt2PBIU37+g4WC+ENUbnG01Qn7gsGR1EN3Hlm4Qu+litVUFXYLmIEkmaXccwg8
9PJ32Gl9mjc2CRh6Oesy+LAAaFyLRlwJDiskR4Bf9cSI0knCnmLfjWNcFdi6X9Sf
RQIpD16kBVvXRECnZGsAUD8VjpI/0e2KWilgs1jPW9vuNYhNvE8kxFRI0SdQ/UVe
Vi7z3M2OcDm2SzbVDo+hmR1uB9TfeUrQphhBKy+1dED+obyvi23V1f9c24dWY+n5
GMeCnSpVF09cVP7zeouUy5ty0kS1av3mSAxOcnI95PujBQDXSuRHr1uYHVgo/P4T
dklVKhzjzz8sMA5wk9ahVVrqsls8eAX7MSo8oyvXzgEI/iphqeILPxe1DUo7JSHg
vFq5Zwxk4pPpQFsHInG8ZARuvy2joKU8ij2d5CN7j5UG6JxhJueBAEa08Is3N4Bg
pFP91NRIIpgTrpTW+QZyhN6uMuXvoZBKq9JnJWKPjx+7E4u8qMxZl+z9fxXbdllu
2SBjepjeHSN2ZfIr+HHGLT5AVJEWmxrCLyAThz7OEeaJXeO4nC86sZLyA6YYd4GI
kQBDFj6wLgfB4hBTaQaS64Xl5R3xa1GqPSGivoJ0SDpw1me0ppwXeWTkeDctKeN2
jWPJ5wXeO0X5KXf9x6K1HxtCDp9FJswLk3x5Bz5lZCLCT1tO1Jz8TSOzLacLuo8V
2XVNWggYrIvRQQ0Bg46w0TUOs9Hzm/k790iN9dZFzbbJC/FwTzchCxVSMZq+1qTT
bGXbeL+igd97Ydfi41ClgxlV4U1Q1WAHqui6vxP4/ZwCB4tlCDwmBzoYx09oabYK
ZMtUA4UQ9nw0wFz+rI7wU77BH0Mg2s1+CXkZvHr4+Bic8J3kHioJbKQxBNqCXpNG
/uG7uvi/5HlK2r4xA6ecUmlbxsGBvOq0vEfPo6lI7S73FkFo+Bwg78ByyrjPdlgl
0cmVHpzxArTA5c0jSQAHhsyIs5xT7e8PC3etGCHc6C8NxRz4RzOJesTaxGkZQI31
aLgBsCsG10n6zefm5/6BAfzzPe6f+njApUb+awnUH/VxCk2XHIRuv8v1Z2RYNZ9e
VFVxRRt6JQdkAl3taUxpWL7wCgtyOLkvYgE/PhroOXbGscmTUmoBL8E0078tVOE1
YdL1CeNTxRd0HmWtGaMUOEPztGEy2IZgVKFnjVJz6zS1GfZb2CACLbEAlB++8PK3
GgdbNzrxu3qSd2RWme9TUQ9fYeifEbYS9oluP5r7P1mL+PNCdzY8jb3vbsg+UAjR
a5RTGoMmR3J6ncB2Uu+/aPeojQMeSRB/T1Wkp2HJVUWZSeItd2MizvcOH09US/go
bSDmj88cqI81JW7a19HTOPvepTbKGWh0H5BJQAX9jbK/0Un3pEmere7M35/g7Phq
q31CjJBF0ysuKPrViwPjAkfL89QNOnvz8hHLKRyYshXh2D9976nwpj0VwAZX3f2J
lWDEqJHZYIzfgVAIPh9yiSMr576u4o5xcPdUhkJOBQIoUzlw37f91kn3QSg3arKb
dGR0n74P6BfJ95MaE5mWAtwPjQJxuEGpivxd6xBtqM8CYefW4Q+m1OOxnYG4z97c
IieLPO4EBEcCkgMg+XSouN9SQ18c9Fz+RgQJZn1i+khwCtDZovSv8iDQA3+Ehgtl
BDZxxMXB3v0+rB1Wr9+EBvtM/Zn24gdF9aTU4fj/SMi/ob/kwHE4dV0EX41dcmWK
3niVSJM9+p6GpczQYOUBbjNxARyMBSj+bqkZJ3pVPUVxW/SyosE6ILmqBiPtCL9M
0tOVkLdRAmMgggbvO4ETzwB02jtA33deYGWkkBwXF33JYaFN7gxtyFGPTQyqPTPP
GVODKkAh9qtvOKU1pSYC0u+qTUP3CgMgvN786dmv6ooj79OfxRLgsR7L7sbTDivu
keYApezZZ5r9+bapnbm8pia3xzNC+LtJJNMRNaRyZbFTta7XpXJ8ewThQniFqwax
g+C84igBLNXAo1qgMQw0YSxzzBZrGQmVVKQLD1ZxUQ8R9pf1VngBojyASlQ9SW7O
1x9EDe7LVQqMHbZOy3QH70FOD44ht9iTBzAnkqZLwU68UobKOf2H9JP1pnGaUDhW
RxmI3D2eX9auupbQmXN/uYglAnIj5Sk/YBkG2t6bF0Cy2TGM/mEGaC48HrXr5AcV
IOw3xa1BmQ8J1z33PpRPbd7cOvnkrAXnIX4yawFgq44cyn66wbII2u86ERSE9d5W
VP59bhFoyGTzEUflFbknpV1TcRzbR4MxPeOVKNehPLjAo0/WOfSW4I5h+Lv232A7
l0atA/7sBixBaNFZtUtLG1DOkdWAf6WBG7wHUKgWb0cBPFU25Gmf7aNVQ997tsa3
m0lwPIpdhX+Jyp8RCoaNAUV+woOiHUeg8HQHw0P+nUpqHN6tPV+y31SO+hUmg66Z
lrseKeo/36c96/lTco+eRByOszXQJUnS0spsUi4vMbAZ0uKAPvs1H+obIoe0DrDy
YGjIWez2OHU2chbUWCqflVgTlPurAt3Wa1lM4CSLLsQDFNk2JfWc/RIUtLSWbmnC
5ldGNQJ6409w3Kg2/WwIYMZa8hb0zusEWD0UzGH0RwPrjHUTJOdYS9La2xx1bE/E
KvHydMu0epW5HnFa96rWxJEo1IGe8L/ktp7epZfS38TPAH7K9Y42e8e9kyDYSBbb
ikYgrPpCkndolbkxHrTkPJZivLw4aaqKZj/jjbLQGjOISnBGmbr8ulTyuqlhSX+o
ypdoioKWHiSaSdukAbQfWWwDmqLEIQym6gytFUokv8ENBieOTa9gZYjN/yCgR/1b
7sDeEUZeLF3nEbGDouoQvQuU+U6YDguAarlPIjaeJHkjBF7LsFhez+hvrlf9Y1g5
PhM/01urz9CgRxGisoKA1i5QRFneaAf9cjBhvrDBXqc42NzSJoryD1lnpyjnYNTD
mbtZbM1zBPItWEafrg8f25TME9v8e/My+kABw2P7DgIBpfR5q5wQBn+jLzP3krk/
pgEbYMItyvdmXGMDA9sDbVS23lcRC/EGCe8v+CrhksyBGXHcsh/2HQH72+D7k33y
k4pfK3Z9xOLdCnT3lZKViLOrkEuliC+EPGTjNmxyRo51Xp8w9RLsD3p7oPHACdZ3
JvcI3Wuez9J17wTxTUjL797p8hXNohDPy8YvKSoElCZvYnk3lULfnoGvx6mWKc5e
phoOiiRui5WrXXKPVRTxRxG0wfjhUdFm2COiwjYAfZ6ZTVSlwee5a2tBEH6EKXXj
b3jiR7a6YaYOmmmWxnE0BjOG0fAbZXm2daP3btJDkJ7XKXB2nu6Hf7EAIZglXeBn
uABSYo2O3voye5ugtK5rbOUUn5/lvLqwJWEKwOaFdV4lA8ymSTtunrjxziihZV5M
xxgAddZJKKXoVfT3hR4ICPOI2Xe5Wed8OORxZcalvK5le3IP/mmQAdIDnbZn1PFo
5Z3Taix1FSqRT+kptUdp0XHpg/pO8fYfO1Z0wZm3Q9sImoRjox/g+hrNacgWxgcr
Vg1jbB7UJ8oUYuRgEnNWaQ9dyUnP33rWRrhShk5lJ9bhYmp4VHGfLlZEiZfX9REv
cNI3NTzMk47meFvjxsTxWkzLyL9L/fTHi5WBeMh7lrZFru6UawRKAGZJKJXSBUnO
tl+XKBXQByfE3AyLWVnL85n6cYt7zUFjZWrpkBc/alKV7kFnsxThwssxvnKMROwH
9Pjzsoh4M3bbRhqyiOQCaO7PavJYpKT/PADQnlmfmDUiLQfplfuSOxqzVKkbyA15
AV8W/fidZWoLQGBRw8VsVP8hW+Ryo+EU0Yo/8TH4ZQM+H2WqJ3sIIW5rKgqi51er
4p7vZYtrFlONF0AY3CjVRchmX1e03uDBe6HKqTqRGcqtemLOsNI6jygkB47vNv5f
cJc/Yl92xLWZyCFNESqJqnSMh8Z61i6QkE/9pbryrKIBhyEqvT2V773Lq/0S0GJS
Lj42H0gsY/ssLtG3rYrZlraR6m3irMR3PnIj4431q08=
`pragma protect end_protected
