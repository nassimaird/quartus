// niosvprocessor_tb.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module niosvprocessor_tb (
	);

	wire    niosvprocessor_inst_clk_bfm_clk_clk; // niosvprocessor_inst_clk_bfm:clk -> niosvprocessor_inst:clk_clk

	niosvprocessor niosvprocessor_inst (
		.clk_clk (niosvprocessor_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) niosvprocessor_inst_clk_bfm (
		.clk (niosvprocessor_inst_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
