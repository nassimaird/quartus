��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG�V�����3͠l!I>v��c������{�^���o���S,�}��I�Y�k��������]:yɉ\hH(�oю�l\�CE�a3~#@E�j#�ED�H��� �daE��z.Z����B�5`��fd�UsGp��e�H�Ef��sr"��j~?�ᝯ>�#B�y}��R����>�N�9�@̘����Z�ȼ�H:�XƺP�:Ԗ��'b��X4�Æ�3��̟�Q��݌�X�R�$��N��K7]Bƒ�Δ/�!l�`}�;~+Uw�rV'�Vu	zČ���tH��.,X^����Ԣ�_P���CB�(d�`	�6�;�I�$mG-P�!L����(V�cs,;12|S��(�g���?H�y�����~�%�lJ���¸�]�5blQ�����J7s���Baݪ�������zrŇƲ�J��m��s�#�Hc�����-����'�{�'ŵ���W� 4���ZUrW��Yl׶�OU≼��(z����[pB��ᐣ�uz��j>SGc��I��V~�+9��B��Mp����;�&����.|#�N���EX{y�3Z���^Y��I��c���J�s�֠~��J��Y���;;����F� w?2�V��˞Ok��%���G��
EZ�����M��4P��&.�=�M�.k�p��?�_�KT���|��|��2'<8X�y�^aLjJ9���g%�P�΍}�H��֜���M��_đ��)�V$_�i۲"������/���X���s=�T��x'���z{���+�Xt4T�7f4N��������2�K̅@+�1=�&P����%�
c2��zL����/�Ҙ5�R�5M�p��q��Oz/wA�J�<�ż���h��Ϗ�}�"�S;l<󍏸��&O��~�AX��gpa<$R�i�����$�g��o�_�˻�u{��}Vӛ�*��4wZ#i�m�Q}�nq�����w�Qp��xː��}����7��/F�2}v�XB%*45�L�Q�M���Y�
���lFS��xϏ��#NW�M�q>�S�sF��.ӑg�\M�<� t(�#|�F�r&��|d�>Ϙ¯ �q=R��M7�2���ϴ2z�0�G���|�S�j �{��.l���
��/�Rѵ����������#��~�rQ*RN�ɚ������3`�V+ZZywi��U����z-ر�ͧU�W�4�ذ𭫓�2n�~�/_Y����W� [�}s%�|��F�e���6��ꓚ{;p{�D^� QiK���z���`[��cy��N�SV�K$����>��`�&Ͻh�n\;�6�G��Li��T-�y˳c^�T'���?(J��B,��1e��l1~�8|f�,��8��i�����2�~�FJ��udt�k?�pW�b��<=h�h�3kuYX%;�&Q��~��?�)�
0�����+�c/�ٵQ�k�.v��h��T�0���$%��/_�7�Ok)�rݛ8�;5%�W�j�)x����17:򭸳�I�� f�S����
9�c��X�R�OGb��՘����6�R�K�Q�o.�ԗw({���%ک��?W�Վ�є���j*XV`�P�Ȩ���a"*P緼6��//�Re���
��F���V��q��i�E��r��+<$x�â� |p_v����R���4�C�m4���� �,K{�������c�d�[�E��B�͆7W���b4>����biF]�s��c0M�Q�)���+y�t,{��롱HoY��ǏgT�Ax�L)�W��3y5���E�_�����bP�`(uZ����#}��ms����A5I&l�a5��}e�i�S�Ջ�?��)���h��.u��[8Z����=�/`^�*�EU��HW�oB�����nz��+9���i�.+v�+�躐�!=^A�G1��YeޙX�\��*-�f�)��8���=_C[ `���rmf��P�Szΰ��`빖N���ю֍V`u���כ��(A��!f�54�ނ�!�M\H")���w�|=����*��h����q����*����Ť��hx|��ba,�o�j
"�b�.��� ��(���2()����Mj��h�.0q5���jz�=3���g��n�k�����;�2��DA�8�܇�,��@܍�8�����2�S�Q�$J����7aDr�<=D� ��~r8�V�J�!-����&��=������+�)0��}�y�'-p��{�N0��y�Gvo�+��R��C䡈�`v��lg¤q�������c��:;�!nu�
[ȟ�d�n�oO����
U�/{�NլU�p��USwܽ��ꚦF���2�L���C��w@ļ��{�	�����ٚtp��ᾧa$v��0,	�fe+��c�����V+��~,�)��������m� }�^�g��<�k5���i�%eZU�S˵�Bf�� (xar�%6�ͣ������a���Q�)/��`�C��*�����q�-�9�w��iwF\�d�S���Z2��"k=�G�:��97�F��O�f6J����Jf�s{^����;x������^�����1��S1L��}d���%�G�Ww�z;g����DA����zlJ�(;M��t�MJ�o~YbeӴp7��1���9��e�~�����&�1��j'.�Z��I�Y����~��Brb�>R�~̀�d`:�6[���>�w�w��= ��(�r $2����՘��QB���
���\j���Q����C�+�(�ӒH��Z�r��� 8��w��^�G�6�n��A&��0'j�1y��C��r�F�UG��K/w��<���U�Q�����n�~�ZJU��i&�K�{�p����s��=WL5�2Jk\!/.��Y�K�Ȗ9c�c��Vf�_a�|�^�[�$Gr�iWՇh��&�Њ�݁�g�\ŀ��R�>t�/�r�Y�f���mM7���E]�67G�T�c�
�@Ѷ@�*�I�$�E�O{��7���q7|��
�ܼId��%��o�/IQ�f�'���f��� Q�8..+vr�[!9%c�m��z7��	���aVS��9�ىS@8��m���(���J�vr1��R�,!Y?�I5���m)N	?��Q���(��ﯧ�DX�y���#/ G����?�(��SRv��=�?'�Dϟt�޺u����n"�$GW�5���;���l�I������2ͱ2T���az>)�Cey�K*��9Z�?�@�M�1���Q�OwE�?�6p"��g>�5_��� R	i������i�>S(V7��Ɗ�[��W8b.2���U��
�bnĎyu�����[Z���K�$ߠ$��L��)�A�����Qi���@U0!͝�Nq~ q)}��	���Q���z �T�L�k'����L?���l� �8e���Ԉ2��Õ|��\m��	���/�x
O�q�~r���7��t��o7�� r&���ik�'X�r��bC=IQ9��v��f����c�R�ʠ(ԟ�~HiPvUϊ�����&d�vX��#/
$}�����^f}�=F��Bw��ZR<�3�乽�(n�Zt����0q[@Y]q?	P�ׁ���nk):����KE���l!w���_�R#t\�9��~40���6�J��X��-`Z>J��ʏ�Ĉ-\t�P��	�//k8u�㊀�B�Y�a.�����	�����Y�
�E���@���SMd��\tқ-U��H=|���ϫgKC/�|F;�r��!T��lk%��@T26B��]��K�؃�����L�iaTEʛ���rzMbU9G,��X��퉮T�>���Oi_�ϛ���}_j�n)S�9��k%�W/��\�2���^Н��i,9$;J(?��o�`3ǩQLw|V�RP�l�ya3�Q�QP��D��K�|�0��L��6TB�G�	�xm�le��9�XW;@�Xg����O@2x3x?D�!$r-��ԧ,���k@U�A:)J� {�!��A��EZXE��rL"��������iWoC�R�"��bTf�4�o�_�w!����B�p��?�8�n�0��� �jZ�q�.�A��&]>ҳ5�=�/�<��ޝy����JfJ��}�\9�V�㜾���` m7�j�H�2(g��3W5do��$H��T�-6�s�%@X�NP=A31
�q3K�uCz�9j�t��nG���A�O\9�@���Q���Ij�/���g��F���9�]'�9JNӐc+�(�d4�{���+�	w,TH>Iҭ?3�X-[�,;�S�֐��2���'O�/��z�.w+. !�d��˔45[9�2��k�<�������L�Cp�9S%�3Ȥ����WT�S��vj�a�q����sV`.8�$�UZ?���}e��P�aŉ��v�!��1v�B�Q�݊xݦg�@CUZ����C�7�
/�`}�f��w��6��|�
ۿ��	�������9���/�`���lڔP��������aȳ �������{�.r5LW��l��\}��Q��E�r����~P��Ц-��m.˖�f8��>L����_��1�ot&����:��չ�*}���H���].��]�$�I}���V���#���
�D[?&���C�:�*d��kU�D�C�����J �������!Xb&��Z�.���\
bo�S�=|LP�Y�~ޣ���^���(��5mBH���$/��,~ �������l��\����֛����ǀcg�xS��j�j�*I�;X���߷�h��Y
��h���q z�[v��klh4��Õ6�K���qk/<�=nu99�'���ȃ�-��x�A��ɑ��:�Ӟz�P�h��w]8�D��K�����iP9J�:����82���N��8t���:M�1�>�?䅬Y�_��U{���0�9NA��{�NS���?hѠh��0Ӧ��*pFʟR����p~d\W�K��5�yTr��k�iWp~Z<���Ol��d�	cO������ �L�-b��'�B�G��v��!�u��+�|{���,.p܈W$,R��T�������[����E�BUj3���JQa�Nx4?�J�����3��p��l��q������M�<"H�E�~�i�i �kߚ�#5��iSv�1t����ց`�s՗��1�)��fn[j�z!�g�ۿxr���R����:M�^|����뒺p�k�\�B�~�l�����h��$�.-Q&�X�����+�(?�%i��O�KH=á$��W9�
�y؉���I5�ypg�8�?-��v��ӆco�i%(�"�A�ۖ�Gd��f�7��~�-F���B�dT7\qI��N�F�Q�P�t"D'��!\�� a!޵�$�$�[���Dt�R���vup�����4wh����w�+\m#�n�����Nu�8��3P�K
f<����?�I�DcR��e@euﴙ�˺
1l)�����RC�
e�JDS pcQ�āA��@F����F�g��QX��.��}T}�[�هZĠ�9V)��\�l�1w<%o������	I�D~�Sw�.�u��fS�j�y��rP�Ϣ��X����򴎈��U�[�seo������.���b繛�;�� V�Z>�:�-�}��2����Ț��2g�R�� �.'$/�<�W[-��	x@"[����ԓ���V��=p��`�@�Uk��ȿz��#������d��������fTV�R�fn��߬�!�x�%�>Ȭ�2R}k�����3�T#���w�1ó@l�@���]��Y�-1R��R\^��tܡ'�qTibg�Ǖ�����Q���Ӂ���D��?�V��BVf��}&�w���Mޙ��`c6�Ʋ#�X��*���D��0�ХE/ K�3D���k�c��Ȳ�,��#��,\����Q�N�g
��%��|a�2П_s���(L����藴"���}AK��ɿU�H4��b�s]��m�D���w%�.�#��$0)� �X�Sط��]k�}�(�Ӈb�f�A��E/�Jd�ǅ�"=ߜ։�Ey�e�ڿKW�N��!_�P�f����9��Q�D���x3 �2MS	,+{W�{^��e�8��������2�<��2�{<��Z����D�h%&��0��i�w��j�[�7`v��>�Q��t��;����]S�^��63�$0#�==���c�l�&@Nj7{@c����6 ��X=9��Y'�����|AL��
Fh4��|���U��wļ��y���;?�y�u�K}�f�6k�2����%�m鋃��V���+��Թ6+��n&��]&y\����Ũ3vN����l�E��;iH�T��޲އZ�` ��Z`�A���(��*qd�����-��z�>D�C ���'�9aP�N����������+W1��M�F��kp��v� 7���
!l�,��β�hd���X����0S� �G��!F�ڦ��
�r��l�ɜڷm�5_�d��iW䘺�2�Z�y���Y�L!�bWAW�;j��{(����S� ACS���)��2��n'�Ib�����$,"�¡A&h�%E�$/Vb.z�J#�~yɿ���+T�׆��G>�U)L����߀�>�1ń%�P�?󛭚��+�:�AO��X��qZ'ǣk#m�꾯G��22?�L���u��%�L��?3��@\+M8����B����[��	��rLis�fQd�����,�ƍ%��P
�X��!3���q6=4��*eI�cװ����y�x��@:����೵1]�%��JfQ���A���4_Ѭi���VB��qH��Є��|����Y$�|��Е)��E���6�FF��'�
ǋ�KH�'����q��PuA|Q����ަ^G���|���+�D�M���<֊�c���N�<	%��P|R��e����O $�|=`��gK�U%��A���1<d���f
u�В��WEQ�̍�h?4���������MŢ�s#��4N���h��&ӏ��g}��b|78p�1\��!-�����/C�6���9�u(R=������4)��vL,u���,t��oS����v (aʣ�Q�I��bR��5Ɍ��FJ@
c.yX�WQ�(l�B�XT�A��bՕ	��{���g�I�Uh���=�Gsb�ߐ�1�>cZ]ZJ�m�q��)�=qL�6b�����vZ��N�F�>���ih�3Mʵ
���� -���������&��;�3��kU���$�I+��1.l������|�QV�o��5�I��J4ŧ�d��n��g�[uX��6ĥ��y-p�DxS�uНy��;J�����;�'CT�H�_kF�M�o|J:��l0��)���F�LG���~��0�5�O��7�I�I��<�n�"��puK�#��	�)Y&����C1��Y�DI���
���mz/��ֆ��V���ɳ[:%�%�u�˟���AK��k��J��y�`��F@=W���UB��C7*�hQb��z�ε�]�H��C6Ih�`��.�B�Z��>�ܾe�Y�?�B�"���R����45\l:oJ���!R�uf�T>��M���]�!{5�*!�3��R刺���� �+�$8�V3���_�dy���=�Ռi���R(�w�BS��L�����z�w���E�.ZU�X�V^�!o٦&Fs���Uv9�߸���a��2��1r�uw+J�������j�0�w%���K�F�ʀoE�s��S��,PoL�o���y�?
�#�g:�=1�s!�!�Q�d�3�X� ��MMܸ@�t
��w���'k��|�jLuܨ�w���q���@�U�w��Hl ��ȸ���Q�n� �w-z���
����ˢӳ���е�!:��A�����a���9��s-u��Z��r���F�ֻ�5i?!r�.�,�(��R��=�5���2���fg�T�O�f���OgjkgdCS�2����o�'�>d�W;�,h�V2��Oz���oC�o��omU#�;�wP}��	��n�W���`�J ��պ�&/C]�?�?)��H��<��i�K|��P�X���h�������fӈ pK���V�b��K����*�qaN�i�� ��PGł�2�ˑ�/��fΟ�A�~8���*��$j�ԺȺ�e�9�٦����1�H�"���_P�,��+�[蔶j2���	WQ׋8�Z�m[7VZDZk^�Bn&JU������aQ��,�||(�����Z�i�̴���Yި��"q�����P������zO`꒟)zx�{�%[�=,����-��C�&�離���J��!�� ���#VR��+'O+;��O�yt�R�~��,�3/���A"8�ܒ�P���ED�/*�"��&QB{s���i���@��xo��2�_�r��z�11���Q�
�@b!e1���fdѧx�Ht��;����	��\�VP��D�s�D�Ug�ǯ�&�� ǜ\�3�T��P�~}{�[��C)���p�O�x�n�%]v���.��
�2"cj�Z"pL̠T1��(��H����і�����N�7���e��b�j[j�Z1N##8Z�J�� ���HT���6&`&�>�
�\%4���E�[�h3�W���>4�qoV�S������#�q��QO��)���ye'ԉS���	ͭO�./|Nev�O�SH<y��XZ�
�39��
����]����:@��vq�������j��Zo9����m1�������r��(;^���T+�o�\L,ue�t�t��AP)b���<��vj^�7h��d�Ig�߷�����q�ge-L�ރy��ަ�9�c*�e�wx>}��0�A"E��&�+v,�*7j��d�@&f����0���̂�������G��D���; &#	�TPA�ȧ m��*
x>��RLugH�k@[3��犯�XI�]�j�n�|��ݮO������|�`o��lG~h����|�!s'��>���:x0$�Y����XZ=��42��ð�o�;��ZnN/@����3�Z��쑵�MS8��fU�ځW״����G�����<�?�Fcf<"-p�J�n2��]�z�7jLx^U�+���H��D��}$$q,�.�����,���]T�Z��ˍH�0���2�ca�XRP�n�~ӭۍƖ��_QE������e@dr?���t�]�F�1�\Ua�/W���VϮ"^�1��~��U�����Di�W��OD��\�`x���`�W|�%ޓ)�PƢ��G�ri�x��˽؎��׈Ƀ->�#���r"�P��Ƨ�v�w��������$1;��A���$���`��cM�k���\�ˤ���RS�1\�a���f��B�Ǫ���Tho�b����D����~F������D�G�����ᦫ��6�J��Rd�ڛly-�uX�ɰjS�:�m�x|	�G`��י���"����0ǀ�M���G��J6 &�8�2�>�F�b�`XI����*ew�A_��37�~�y�T+�vH���k�p�M4��v8
�7�o��9|r�H�v�&�JAW�UH`i���k�N���߱��C\�Ru&�E?2�i�|gSs-�"�]C�����>Db˥tD��N�:����A4G�����M ���X�
h�Ӡ*��^#|"�`~���>�<��g�����H6�C��k��/���"���1Ų���!%K�%��!�����Zg3���?�igpB�\C���^�]���k;�)�ؠ5�YJkuu
2�;��w�N]���@���[n���zۺ$�3�/���O>��g'�
a�G{t!�l������]��~�o"Ď�����3���A�3*���Z�)	��D�f�˲��T��]'5�}N? �4���e>o���0ـo�/+o�~SvKʖ)evFF�X+�3he��FgE�zY�Y.�����/�}�
AO�E��� ���M�ޚ1�0;b�g(�x�^y���PB3��|I;�u����VL�{���.�O�/(���?y{`��	�h1�D�l�"�sUu��i���|=:�-{X�o5q�"����	pgV�_��2M^$|[M2mǃ��<1�"��*۲�nĦc7�+�g��4�z��3� �Q�7���C��؜��#�;�&��j��+�H�겎Q��A��j��o ҵ���z��w�����6px�NA��9�O���@"C6F@Hm4��9�x �E֛�w�_1���K�|+]Vךވ�#r��O�BxD'w�lc��*/?^��!q� �$�09�C �_���������f���{�q�y֋/���G�C'wV0�ƒ2F�1,�*㹩���Q�E��;#ߍ�V�Eq����Xe�����}��/��Y�aԃ� ��A�?��)���ED��\��b��^R�M�z���7l�{ކ�V�m�2%i�7g"绍3�E[����kB�M���!��ؗo[N{���!4��?���g��]6s��e�䨽����X�1�����,�3�ٝ-�������,���Ћ`KUy���)�,��S?�ָ�v�ͥ�})7�[>7��{�gZ��,��I7MnU�a%�8��"�q�S����O����)C��T^����[-�F�t��LX�-���WpK�xfŕ�3���B�4*S�G��QJF�驛.�.d@�l�U��%_)�-с���% !����X�ɗ�5c��P�GI�$a�%��L䁋e��y�U`�p^v&��K����� �ƨ_u�S�o�ג)����?(�����O��@0��ۅj7n�-��!T_ �7X�V�4M�#�H8y�e�"�C?�Q �T܌�1n������D�]-���@�U�g�}F�?n*Id�]}�-8|���|qcn>�q])�W�i�t����q`���\�𕷪��Bz�*;�v��Z=FM���f<��ͷ�g�5%_ic��8�����Rp%>"�rf��D�	�T�Ҏ,�xv�?ҳ�|�S:�g9�/J|���􎙮�3��y4R��(-)�ѓA��J�\����0+y�grGh���JA��/�m���0��k��f�O50tz�F�������O�=����B&%:�#�+��W�{߳q4�X�L����MwMF 3l����Ր�EoU5�P-J��/v���N� �6�uI\<�(X���Qk?#��n,��SbX��M�ύֹ����?���)q����tyuZ�4���u�DOOO���΄�'F�:���[Sm�*k�9d�m�w4)(P�l~m>U(q��h�`��\1�^ԭK���v�je��3���g(b
x���xgm��}Ȼ�-�7�"%S�K�}|G�ۜR����+.��]�b���9������l�1f�X�Հt�D���2_����Vii�s��4e�qA�O������nu��.���h��gi^��¼� ����*쎦#�͘t�,T[�����Z �����\Q���IӁ� |"�2c+aWj��M������*����k*tA~yC{�[�-�KL�j�p4�[�D��)!�5#Q?�y����},`��Ks��]h���=���gyj�n�aw5��w8#�~������:�A�l�eX ��&`��a�pڋ�n8��TG<?�f�$��7�CycG�DJ^6��ǵ�M)��ո)��	m���/�kX�&*6�;眢a�^��j��V�#�I�{Q��O�R
��ߌ�;iE�N���/����t�Lֳ��;,2��k�-$t��vs��G-����=�q�Ԇ{g����:������Z��G|ZS��}?����4�#KH��oC�)V�^q�b�F�+�Aa�d)2-��a�		{W�eM�n�׼?���;��u9����n��@���Z���xh�b�!��K��g���p��"X�&)-��;�%I?���
���3�w�G_}��c<ǽ��g���溠G��g�1�aVҍ\��9�%�`M���:�ߎA]���C���=��y��E0"�l����?�C�qr�[�n���u��,��Ag�ؚ#U���]�$5\?�+�C֘� g���'�@Rk���L������޷�v�+	�5~���������o����R�b��_Sy������*y%���<-�&���%�;�J_u�a^�	�p8�$��ty���]�� 34���/3;n�o�DZ�����G����D|�!�nJ��P��ۤ3��|pY��҃Sl*j�]F�1aKD��\O=�8�I�� ���7�G���W���?�i���[�)#(�B�_L$Dk&WBd���_OKi�]j8��P����L.!>F�mXeP��M(nc4�?9��߳:�/2�.�WC��=)PB���f��p�)ۿ{�Ib�a���Y���D�,�c���On���t���+�\�С|ш?���]4�M�K9��yӯw%ļ,[��B�[q����&�Pپ���s��dq��S��;=��b]���;�R���C��p0V4��M؈�	�S7憧��X��q	�scQJp�ʙ�HK��O�q�&��!z(cX����'�����'�Ϟ�I��%��,�fm����ń�W��Qԏ1���}�p�|.������;e�zw��*�{(��Uha�l���r���'&v��>�3�pI>��ig�xR"��/h�ug��=yi���Toۑ1����kR �TIb�� �ܼ'H�Qដw�G?W5f㞄���l�[+7O�����j�?݁����s���]��Va�:����W�0�Zw/��7Y�B&��������� 8�W�e��c
�[8Y�ǵhz�ݲ{�a�E�Es�߄�O�A:S>��� �-g��6���-x�Jr���.�>�C�V�6_�4�U�M���jF@�V���U9�sTv�}k��}����E�'�Mf�����dR���-�L��Fp�\.�0�a�h��SQ�Ǳ%��5_��%���$!�, ���ԕ7�r����u��PTr	L0x���EiqS}h�r&����5K���v{�v7�P5M6(Ru�~\Z\���t`��D�����47����3s嗷=�иj� �4�K$ǒ�"�
��JP���D9R�b�y�gy�Oo��K�Â9�#��JnߞO�����I��ô�!�6���������i+�8a���3�p�������R��F~b+�+��zŞ|��y�c�@�U6��4���?�U�V����?���gz�[��_%�8o�΅�8	[�t�L��\w����!��^a�$�㓙8G>��|c��Q���5So��XX�U�����~�LL@��YO��R}�v'��>���:<s�?�������6�����\���r�b�d���#�x#���]׊r3��x�����)n�[a�u�9L�3�B|5|��-�h��	&�3��_�^�b�CIJY��O��?�X�W2��:�@J咓�`'�Ҿ���`�$��eUV�B����1�n�F�{���[u*Lt���cn'���Ή��Z9s���>��HA��ĥ ����`��R���x�$���}���l�MJ�p�r�զ*����ߓ���=+k���4 .j-N��+]��H+�2���P�r|�e��J׏?��������n�.)�L�SHԞ��Z�<M=�E��nT���m�,���dO:�G9�4 d$��Z}�:6����Z�A�U���F�94w��ģK{�d�_�h���L7L�$.>�l&�v�"��3�=�=M���3EW,㹧[NA�0���mb�PuFO�CSq)��-;�/#6")�}2l�2�vc�C���ƺց̲Y�ݦ�f
Ķv����#�x�']��f�$�E���'��BO��
�B6�ή��ᏛaSbQ���u*<k�u��8J�Ӳ�]I��(5F�O9Q�����VDϖ�IMv��q�	�bew�o=Y^�����⻿e�����H�`"�Ų\"G�?����t��ԇ�n� �:����[:�u�%S�=�z���ݣ@�R�r�j�/(z�NXu��=��^�Zb$�,����_���r�;wڱ&�g_ ��L��s^/��(�bp{�!%��{���
� @Via�P>~�n���UM�T"y���O�g�MC��\��,�D���C7��IY�7$WߐY��kq+#M�Pj���Q�]�O^ܙ
��g���D��'��#�q[����b����x�6J��`�O�Ԭza�a���Wt��~�ש�3�,����j�M�K)��k?��Y�0tٝ�N~��
�x8��P.cb{#��>SϽ�N=�H�4z]�"���R��	@g���UjJM��u��<ޤ�z�O���L�r�DO�\2&~6�gru3s]�X��M*�������"�q@B�jFp5vh���J=]ޖ>#s�-����H����a��'�n�;A�.�keLY:�x��AȽjDGۛ��T�^�N�������pZ��\ڀ8�Îw�"HK����{��H2N��V�(�T�"��y��P�6�z[�.�r3�&���2<��%�#�ws��[�<cZP����X��݁����j՟r��V@���ls�נ�v��2��mB]�Y@�>�LQyGG�|(���M1�d�蹠T�"a�f��.`�%G<�D[�n�9�t�3aT�:�����n�;�f���v��ϫ��[;q%hp�S��)VT�dv W���,d�F.���e9���7%I�iqv�V�k..#����O����FY���>���<)T��3�<f��YK���*h���e6r�����g�PnV~��3���H� �Zw��j5G�4��C�2���[C�]`t�����@���'�^��H&ZB����wW�P�P��
Թpo=bsE!]7��8�j�k�e3���q�еLsg�?����.:��vc�&�)%ho���S�0t�yf ৻ƒiѻ�0�pc`Nӎ�q��H���"ds���)����B�n&v~��ߺ���ĄӔX�Xc�t��&p�&���f8�)��aRǿMӑý�uҚC.ݲь
'$���f�@,k4�puL�옲�;�>��t��f�z�<(�@��{KѣTF��$�b��<���k�k�l�)��9���́�U��ĩwƷr����k�Q��,Prq�)����#o�i��q܁$8w�6	n�ի�8S��X�v�dv��2�QU�.�	_����X�tl=k�K�+Jr���Ug����lyQ,�MD�ތ�8���6clR��t�kʡ�hJ�Ŗ<��v�"�BjB�R;�2����ɤ��Ώ���zm����h?!I_�X(x��l�Z5}F<��("}H<.B�+$2HSSL�xF����G�sG���h�'dKF>���Ҡ��	�����P>�C
�r����JԢ�d���,���ap���g�>�:`�M����d�
�͚Lz��uK2!�y;�6�#t"9�k��!��|�I�v���8_��	:d�57��I|^;��r�w.��~xA"9;�\%�#��������iќ}�lY�-��d�C�#���{I�k�$A*�������l�P���r�=�7�aRÂ�B5�TS�Ƣ��Q��������~��ߌM���r�)m��̠�\+��{-%�N�����Z�mp�,��݂���_v7�)�������Nb��W��`���T萩���BfhWkK�3�*3�XF�q����CK͖�FA�L����	�U���eŇ���Q�3���m���J"M�L�ta�M"7�����YN��`TlX�h��S�,�.ge#�v����{*�T��7s:�;����yc��?ܼ!�x�j$^�Ā_f�����Ў�2�a7�	���3���J��)� �r m��(H��ݜJL��َ�CVG�є�̀�E����g��q�7\�~�1�qb��/�C�זIMד�EjsnL�*`�6��OK�cz��3~�h�"p�F�6��:'�y�m���p}���Lü��{g��i�S�@_IѾ�㡭0�8��<��H`�dc'�ó�V%�m�_��R��^��@<������S(ó�O�t}�u����LY*^6�K�k�
ע���XA��)t����)AJ��j[�U#�/?C������K��}9�p3Lȉ
Iy��b`�8!]�'����-}Mn�����j��j��}+f'SJ3��s u�v��0<'�T�T�{��N�f:�q67{�'t�Hmh4�CoБFQ��I`��ڹ�XJ�؟�X�b��uHdv�;,=��Si"�X��D�r�`�	���F��:�h�i0��˞0�1�� �0�]p,����&ꕹ���#8�jʓ���F����Ӑ�n��G�?�Iugc�,�M��uϐsC�/�o���a�h0r`=Wi���<���B�u���u.󳛩��*�ƬW��p�Bu�����w�P�)��Y��M|l<(�x8����k���srU�c*B�L�{Q���3�%-{:�Wǹ/��%��1����*��Sם�o(.�B8\��m�����:���EQ$#|��R�2@����.���"-�4Η���~5B���98�L�����Ŭ�w�[��ǁ���g�f!τ@�7G�����S�|�](������/Q�gI���{Ѣe� gL�ۨ� J�p�a!#��	�/��՘ɇ������o/7��3��Q�D��h�M+Ɉ�p�nՓ�xf��h|�0�����ϖ�G����E�J)?����2�y�Ѓy��)0,L�*�vP���s�4�}Z���"���`�}����=o��/"uD�Qd����j�f��BY��Y�ڜ��"X���b^p�X��v��Lw.J{��5����5�]/�9���v�Xߊ|���1<�{�à�/r�U�� @�f�q7x�y���d�|ĵ��^ji't�8��"�;�)�<�x����ɓ�ؘ�d���Q�x迦�E:� �N� px�o������
��R�͒�F�<����'ٝ0�v�;b,�g��D^��|�<�mM#Mu��}�����H��*9Y��ו�g_V�?��.��P�kU=�c��JE��;j6��,~�>��|I��iF�e��
у�f���`B��s��:��U]0=#��!	d� ��ܖ@sG(��
�_P�*��h�H�n"��d��σ鸣Q}��m�ͪ�|$�~��/	'�n��𘡓�4����#د��+�]��xB�>����ۢ�6R=�}(���6�S�bTQH�U��(��f9�=@m9e��\�C=����0a�ݏcgV��-����u숫���e��؆r�v;Hx�>���ɪo��>b�GM�-��Grq�t[{�'�%��jDȀh� l�'�fE�W�D��'��9��˭������n�%����=U����g����cJ�ghJ6�>Ftݡ���cg2�H��PVt�L�ͻ'�
~ۭW(z�� �W�bu���9}'y�H�ss�|2pDx�8#6�6�ײYg�]s�_!��W������D��l��Z٬�F�V�90���I*�h��{�uL@$͉0	���i23c����?�b��N��%�}���):�@�{��?mXF��S6�����+���0Q���p�F	y���,�[t�:�t%8@+�~c�&]L���r��r���k���y�*nkU�+A�[�� ]����'���l�D���i��s��l>R�KEU]�z�u��t��2\٢��[�1��Ƀ4�t�P����ŏ����|����R��e��Ȥ��ϱ]������!����Y�,V~�T��|!�1���E+,i�usE�]G�V��``;�M%D�ୡWAQ�(��X���p�z6�� �ۤ��8���W{r2eUa�@˒�(�ŧ_M����2��G����?sw�)>ju�N�.�i�X{&ZD5�y�u�}5Y2�4���>�ِ\�{��!���n��]Ვ�j���8ȐR�zUd�a�[�l�;
�J�W5�L�#�-�t�-/�4t�.�#%���'�'���Ep� �@��r��7��%��m
�ꭹe� �d��+6�w��8��e�y�����暾�/Q%-�d3�����,��C凜f�"!H(�G�(��%�������#2q�#N'���^T%�2���Au@<w�v61��f 7��Ͷ��/��z�DysQ�#Õ����Nd��G�oٯ����|��f�5�D[`Us��u�`�~f����T{��`��f|�Rh��%�3���q����1�g�!�"�B��H�&V��=�@w3��2�����-r,�B�� ���9��*�ٚ'4c�����TK�u�1����o��f7���}DUnd�'Z=�D`�[x	�N�'N�"L���1��w��{�C���!)��[_�7]Y�,8���DPm����~��S���F�D`��c��9~�����J�r�x�e���~�%�&f�G�S��^+�Z�)�*0�Z�W�I;xa7j��k��O�>�/x�y���7m�i���P����b��i�T���>G�!������~�mO�f��u�^.��@/l��c�*�����$�x�T��,�%�������H�w^V����/}N���~�T�����D8�s�xx��(�U����4j���͹��Y:$��h[��-^�|�<�P�Q��2���;�|BI��v>ߌQ^&L�<����:1�(�$X���J̡C�!���'�9�O�8^Cy<�E��%pI����g&Zl�aG%�k�d
+f쮁龱4�W��KM��)�$�bJ|7*��f������\�㎞�]��ٝ�o���S���j��q��7��$��W_+T$5�(�Nݮ��o���Fa�y'�J�
ܐ5����s@��/��;Љ�bXu����ˡ4Y����/��8��2���>�~U�>�ŖZ/���%�C�h�C�C����~�	k�����1�G-�J5�6�BKk�M�G�22O��Qƥ@��D85�)�F�m�b�c��*�d邆W��)�ۃ�&̄z�x��}��g�.�g���o���=�2W�9%!'��S	A�Y7_]����ɩۭ9�k�Ήz��'�!H@���-F���u-�K�d�=�Mk ������;�X��fB��|�٪�$w���~zp��<�z�C�xdۑ��QP�����Zƈtڧ��X�2��0��SF��e���S��G�&��<�{���Jl��ќ`xI�w.>z�f�P��޿c��<�a�=,���c*P��G����#��lF[��Q�m��@��D)"�5�v�������?�?�)/.RVp��)ɳ�ķ=�r�2�M�����A�M2!եk�V8Lqk��&1c��yY��.�J���� 3�~'�tnN��ɸ�tKM�̧�w �s �x�eX���0�*��_5n���,��VD �3�Ɓ��7��p:e����G&�թ�m�4.�k�,�\��!�>i "�A�p��b�ڎ;�v��@�"�����F�H�C�ЈL���a�̚T*���v���|�Ɛ-ʯ�/�$��C4���V��I���+ߩ藘C�x������|"^��R�����sS��oMwK��&���@�u�u5pp�@.��� �!O_�1��yf��p��o\�6����!�̒����ĭ��!�UEzwǰ��ԣ"�<�(�ws�A ��@�@��(���*I��`�4c}u���� <c\qkc_�����Q��K�]xV?�X;0�Ѓ�1f*�Bv(��y4���$e�y��K_�̊�R*��w�5��f��f@P�.�LQځ��=gfŪ�~�}�C=n��D����F��1}��>,�l�V�[Ŋ�K��`�H;A����wk���` P��T�I҂Ud�m�����ڕYO�.;�p�3�lv+K���!Oݠ�H��Z��TW��m��=�o;�C�c�Z�S�-ͥ�cT����%��79�(��ʍ����T�������Zٝ4-\�����Zۈ�5e�s�����=�ع�	�q�km<�Uj���B��`�qg@ئ���%L�0������p(�����l���>;Hե��tTF��6��c7�ܹ���1�
�w�nJ�Å�{���q��3��DK�c 	K8��"�	?D�O���|[�2qܳ��A�?��踋Q���w� ��$J����\�]i��m�!������_JAPV D�܀Etݯ��!L��`�Y��(k� q+.}]�E��/�$8ha�x+-8m��=F�`r#L�D��RR>���`����W�6z�$«U���%``g�(q�m\�_~rXO�T���]r� �-�
 K���ʏ��#�"�/�����u�d����[d\F\%ϡа��&����K{���H��4�k;�PƓ���9T������x$���c� ]I�yV�"N,U��*��S���z�:E��wdN��H�|���}�Yɳr�3sћsf��3���n3�$���(7s2":TIw�[F��ݱ�F��y=����4g;)� :g#�\U,��:]��f�1��X.h֯�>(k��m"�x	�P|f1j��V��[��B_~���?x��s�{��o��C?�&JɆ�4]7��٣N��L��;y�-N8I���tS��z��*�,���!�X�Mə
�#�4D���Z�x�.�}4ܖ����!� ��p�o.�#(x��/��%�~Q3�p�?�+��4��x��$�+�	s8�����91H!'_��!�I.�cO*�a�/�3��-������$�p�R��Z���)Q��"��f���8:�4R�\^�N��f��Z�䅵�u"4��Qc�k;.FS���`nӇ���i.V� ���s�:B����Վ��*s��o��{���t"�C����*�S����g�x}�����;ʩ@����wj��p�����43�*��_��bz��0��U]/���U����՛���?Y��Q�w'��b-;�ש�t�ZO��'V}���x$�E�!���S����-��B}9��kX<���pO����OYQ/�q
�Y���[�	Ά�[gB|u��		�[�?P��y�ѧ�NE���hl��az�lLQŲ� �O��.��Y��1-/0�P
;?��'�K�I����@��j(`�EBr���L��	����iE�G���ӱ���z䕟��Ќ0�󢚬G�kUhɫ�Pq:Y��|����DE�!v:Bj�D��ă�M�;]�5GexRǋ�T}^;w#]N#i�����y;W�Տ��)�J�G��l�e��۶^��B�M�b,�ͼL�]� ��d���Eó��B��P��ۇ�v�D�Yi���	�ǑR������>��t����!���4W]!�A;��0c?Q�ڜtW]?8�?���r�Fu`���1��R�9'�}~f��S�C��ߧ��c�W�LA�aPMKm�8�M�J*I���]h�?qnn^;�.��������<��u��w h�hD��1C1�x��Q�6���~Ozߝ��}w��WDO.�3 ���@&Q{D�w�[��E2E�����؇Q
�o��"�P�+1��)�*�èQt���/���S@/n�!�={H���'���F�♃��'�ǭqD>�tL0�Yq�O����+54�������Јq^=`����v��5�A���C
k�[\N��̼%���V�N!z�*ө>N�t�7v���*v�I$�sqQbC����1��n��	v�\��Hi���%�v�Ļ瞱���ߖ"����ɼ��q�񼸣��f��N�`�X��H�?q��"�+9T��
�ώ��by�� F{Q�8��'#}�Z�poI�	�H���;���ˍ������O�!7.�s�I9Rk��Ϭ�[90��0�/�[l#�8�KL�d�W�Յn�4����/�terӧ!��>��zF�*��J�κO�R�J��Iddj �ܓP���B�|�����z��e��e���V�*��پ'K)����L�D�v�ȇ�h)�ч칏C.�c��+�֪��K:v(��Y�߯�p�<	ߞ*TRC��c�'�*�)�@Ԙ���2������#S�Zr��9t˸��NU�����K#����z�E�>S������c索�`ԝ0�������}�(An�qU���+OІ���U%�O���&�|����S�()Ơ�n�S��͂b���	���T����BF���4G$�"��m��+I��L��ɸv�����G�Uh�.D(!ۊ!���m���j�VOD�W��;ȷޭ�Dq�����X��^,���azP� sa�ɋI�i���G�m�{V��1�X�$�UrK��4���XT��`a��ԧ���K�ޘ ۜ�dNYB`�����1s�ixܐd*i��9cG�5u�9���J�6�&�w�Zg��bb��A/*�YZ$SN� ,��j��QU���n&TO�+��Z�N]��?�,x�bs�8^O��T�ҏ|�-�� Ɛ�a�����ܝ�?5�޶1�l�D��nS�g�Q�1�캒\s�4���R�&�a�D���0e�7QӾ���c��7��Qy����l��/6���XL�;)/T���SX���C��n�O�^�_U��_*G�5��'����Ϛ�x��3ڎδ���K�����p)R�lȉ��AT�騯U�l/
VSBEW�`�$u�Q���I�����S����HL1�w�
�r��^U�o�3�<�B2ؙ|���L�!J�{T.�Q_;<� Ì:����:޻�
�� �AU�	�XC�Xt�i>7���5f�R[���f�ǷF&��h�_�N�g�3��_ŧ���(�@�pA�4�̎Z͐�Y�.r5E�-�DI�'��;������2�`(C�hg�X����'��@��AP?�Ԍ�S�
7���H]T��K瓖�ju0���&�8ʬ�*����*{��A��p>8N�a%��F��e[d\W�+�!S��Kn-�;]��Q���� L�3|�NzA�e/����7���8��*�x�Q���rƋl/bW��scx���L������t���,yͰz�,�G�ىV�\+X ���:�m6���^��u*9F����|�"u�lKW�v@�mWT{����.�*�&H!�gI�!�kfz�T�,��n-`��O����.�펑bQ�tn�:j�N����u�}7fwt�s�gbI�O9lw�d�+��R�V���.���#A,%�݈!��wQ[�o��Pԩ������y$]��d�f�im���IXصo��|bf9�>�;7��-ga֏4@f,?�����a:�tr%In��ٽ�h"�����rSM�?m��1��s�������Ս��lS{w?ʘ����Cz��y��!��a��
E�&%h�P�X����dﲱ�{v[C-uL@n���5�bw��#mޝ�t�K�ש8�y�~B��	 *�8����Z�d��VZ��b�-T0B���,�C�.��:�=���O[/�jˢS`ׂ�=2~tH)�!���k��@l�W��|��AykWjo�X���M鳨c�K6cQ
:�ܲ�e�����Tc�#��Q�KЬզ�|�:�KR6k�4�6xE�[M�}er���h��v�u�5Ⱦ�9R]����t�U��X}@xH_v �!�>�--���e�Jf�9��(���ͨͮfo�$�k'��%#� �3*��WI�{y��8�"E�#�T���Tk�Q��i�*b��K�e�s��"8!+�;����LV`���sj=�e�X��d�!�й�7�o`%�V3� {+վ@�-��83����� �B�+wG.� �SiN �$�����'�Mŏ��������<�O��FL/�kdF�����e����]��Ȩ"�p{��H��"̔�
fnz��4�
g���-���D��<��r��3�0�y�*}�D���3��xk�fi�&�~+����^7=���AhX������b�?��;T���l�v������aG�����e�]������H��$f���(鰴f���+J>���SLz��U:pIцա�A�M��M�Q�0�1[�O&h��ΐV��˜w1�eC���u{�囷�ާ�����nY�����ݚ��i<���	S;QS#���N�Ϯ:�I�KǊ�-�"c%���1�(��e�5V�?k��h)uSJOPo���'T�#b��}�Ŋ�~� *jš�G1ڂ�L4#��]�V�:�q�K9�$(��`��oWm��΢@�_�P�t~���#�IkW��.�0�P�e��?��톯Ci���'�E�F��M���Aϕ���U�6����U�O*�^�`x\�>I)���xX�Wнg9x[~�����o�����{ރ�[W�~s��g7����ω')�)s�Ԕ��e=�h�����xa\�!����<��7B���'R&�_ɘv9f����w�w(@��E����de���(� �����ܗ ��Vo,t#���0��]=J�'�[���n�v��%Ok��)����F.��;�ig����28��xԩ��5��@Z"�	b{��M⻗���L��9�a{�A;�C���3��yn��4;�y[A<����	uΚa|\.ZARYyJ��K0�	$�߇O�fe]A<�y2A���/0��
�L�ˉ0��	�� �ٴ�&��~��S�(s�@�)��f�
�On{X��il}d��q34o삨�L]i�qvC�݇"����푟[@L��e���2�.�X8�A��Z���s��Y��"��Y']�+(�T�gF(mg�[���85?.���˴X��/�<:D4�+E��� !C���1�K�q�77����
����5+�k��ưEU"m0y#�~����T�y�s�m3%Z|�G�[cI)ָB!q�v3O0Rأ ���}�#�s�3��&ErL{�c�'���y�@�|��\�̺�&.���g~���gb�����M��p��Y^�I�������b�Cl�/�6w��["�V#�����4A�|#�����ō%�b�&������2 �So_2�N/���D6��
GQ@Vʋ�ВA�>�~�@� �!3\���h5��$TDvoY'��4��Eu��Aj�t_���)&�Sm\]�Y{��B�P��k��)�:Xk-wr�߭3�����o�C+@j��F���҆e������V~{����_��Y��	���^Ap}U�8�V�<�i��mf�H���(-��>,�tQ�v����j�R>B��m�?�q�eݿ�ÿ�@�a.j�\qx�},��nLys16 �"�-LAʭia�?G^���\�?� ��Z�̭]��A��۵>�@a�;�ަ4�_�N���l{�'��&@��	u��
�@��k��msQc�Ŵ�� �qV7ץZY�z{%*�b�5����*��;��x�&��̀���%���H����9�q�IO! j��_j�$��;E$90=���U����:7�����%��fPu�9;������:�㤟�TR�bS���H�I� j�|�_���}G���1 {� ƿ��	�C�wc�p��8̍�W�L��r����_�_�,��|�oe��#��L,�q���j�M]��r�F��x�Տ[l��"�ko�vޟz���f��/����[�� �R.�`oV�UkU9B��qy7����y���
���X�0�;��(��,���Z���
)o��w���M��vR������I��Ǩ�����p�� ��*�����܌K��\�*ODi~g�eQ�}R2ձ��Ģ�q"�a���V"\�1����C�YO*��?ʸ���*V�9��BФF��$�����;e�q���N��9<�R���!�\5@w�I*Ez�LуUZTR�Kf@B\n
����`������*E�*�<��uGBMi��&���(�����3��E("/��ɜ��A�1�4�f���$oѡ�\Oи|bp�	.��䷆+Mp��������`�%�o�lC0��drw���.�ʕ$k7���(E�ت�e`�I���F�=�~�^�2�F�\,6�<��\�b�m	O̬<���ڜ]�o���X�X^����ڳ=��}������ЗfE's��=��R���À��lo��-?��
mB�gD��(��LQ�P�q�,`ۧf��Q@�?�[�u;�q�<4�mGM6�Q½<�; �{go�Ʀ
m���>5���#��<��=�(.�a�d���m������>����M�ЫĊ���q���$Rt��M7�_�v;T������� �B��Eؾ�w$���&�h��0�U�;�b�]��L��ɴLr9���� �ky���!�m�G�ڈY?�"��~�l�_�O&���d�TV���LF�g����Nj�E�I�vREQ�����Hq����:�כ���Ë�Ȋ��jj�*U>:8]G�K�ƍ �Ln4���]��dP�5I�����/)�K�"�����2�3GB� B ��+!!F�M�LX�j�~�N��T����a#����I���1�!��r+����ה,%s5�Ы��ͺW�}��@0=+m�x`ާFeK�����u	,�p�Kq�n�/���Td��a�jP`�P������珵����;C���=�ݍ;�q',ΥÞ7$�f� �L(���]ܼ�q�܆�>I���������^����B8��L4T*)V��iD����*#S<�hȕS�n���n�=�N^*&J^t�7[��y%����ah�R��Gr���AB��ں�6��L�/�ּ��Pv�Aq����X��y~���ʯ%c��0�ۑ����2_�/��h׹�;JQV�6�G���&�.�<�B(��aʥ4Ba�-��ۂ䷖���V���8�X��,҅fm*��	�+�1k�sҸ�����B�YF��G4!��θ�;�i W��D~N�p}�M>�1�昊̢0@��2Р��6�%O����na��~φ 6T�w���~��{��)���9��pt;
Y;�us�kq���?&������)9����<�'sɁ`�c��{��p�h�Y{@ރ+lTD�Ɱ��6���n��$�)1!4��,�\���
�N3�:�7J��T|0�72:l*/F?̀[9�n���~ٯL�y�F@�� V/@En�m3@G�Ery.�d�t�����)�T�>�o�Rh��=��3O�U��F�1 DY�5��cT"��q��,J�����qܱ�8J��i*Or&��˨����!�IQrW���듄0?�T$�K\h9����d��'Q���F����7mQ��=٠'�\��e��R�;8v�p�<�a}_��"Ez�<��C�]Uʆl&�A��^0�0WI)�Y37���\�-���nQ��]4w�)jrZkX�0��(K��*�h�W�e�k8�Cpӂ�5.������~��� ���AeE��á�<�����Ha-�W:'Ym�PLHg�y|>����z
�؆Pda����\LA�$O� 7M@�'n���:H3�*{j�v_'u�F;��[ a�r�IȜƲ��95�:��(̕���;�B;��9��̅뙲�ԫ�SR�?�Yx2�b�>%'Y<P��˪��S�]�y��_��Q
�K��0B8�&F�L͹��E�b����$�:~��l,���-��J���ݿ�;A�L�L_��O�@p���R�1�
C�*�/b.�A�����F���#�#�Ώ=�+f���|ȶ1�������5�tF��j<��ȟ�'����{�
�AP����r�8�L�ݲ����_|�>x��X�%(=Z���7��CS�ʫ�>�Z�,8��w�	���9$T�"�uo�����q�i��Т�S3kX���h9�S�<��I�J���o�)h}���F����d���ħ��B���5D�f$�`v��g�����,��c�=SDaW��QMm��jf��G�n��voh(�G�$��'������V��t!��K#�����l>U#���/{{��@���~��Rm7`��^���xGP�;L�T�J�*14�ҝ�A>��m|���Q�n$�I;��XApf
���݁�\�X%.�c�����FP�c��.��5X�mPx �;X�aՇ���ʊ��Aɝ����=�,'�G�Q�U�b�+��c<;��h!�GC��B0t<6%!{��hvۋ7-s�w�k}��OҴ���L:ܜ9��#SC�~���ȏ�+���Bt�I�.�����SC�N��*�Kx�ȳn ��EI/��#;M�%,�Y
4���/%7�ݺ��E��>c�쟑��}mΐ
9m]�2r��3�[�k"�-D=�k> ޲:\r�R�ni�u�7�y����_}ٲZ�����p�375�r����"	���-\��� #�L����n�yr~��IURM��:d�5�V�)~���O�ǎ�J4i�"���s^��Ă�r���r�H`Β��EF��g��}�ɍT'Z��IJ�7\�@wB�I%��L���O$@^�*��\R�zG-�S��6&r/%X�������Xɂ����U������,�Q1+��~�C��)5z��b��b�P�m��LY��l��w�;$4R7�S�%���מQ�s@j�$���-:�l�+h�j��b�0h�!����`�".��Kd�|��ާz<�	j.��^֚�C���pg_��FßDİ��#��V�Mq,�b*�@g����G������␲��-RF�p	��BR�+&�I���(�S����������M�R㉇tPmr9��ד��#�-0>-&="x�"�t�"O��/�~�CI5�Q<YT�,}���V�ܗo��xG;��O���AӜU
Dq�NF� ����'����P6	����=;�De�-�p¦��}U J%�	+��A����WV����Z��fn�Q��F�t��(#�N���A��7w\�NAm��� *%��-�La	e�ϛ�=3a��b�,�;���zR3�a(Y��1[c�7}��__�<-��}��&WN���3��T=}3�[����	ɠt�͊�w�cF�n|�R������쾘�^*����;�Saj�^G��s8���]�a�����w���>lnD,�}�z�N�����+Zm�.z������pXs�b�d�%��h�5cZ�X1/�mѽ�88���]	�,�1�2��{�@�=���"qZ;[w�N��oZ��I�5��)�2A��7�o..���y��|�q�����hD0h7�p��ġ�R;D�Y�a|Ҭ`&�f?��9(�n<1Op��ZZB"3��}P,��̼�.���g����!KQ��|ى�QJ�Y܄0���*�k74RVK$Dٳmή��:�pc�r��V��Ad�t'i�06����*^qًb��ɴ��fQ��+!hlb%�E�U�Ī�hF��#Ѭ"�ZJM���k��|�,�O��W��a�&$+�G�O�O����GI�v�@o}JT]�66������74�^%�F����$#5q�,t�g�-���p�s�
��JS���=���h����m��P��g���8�7�VH�X�r 閾~o%ڙ�h\��n�rl[���;�=-�<M>��������D��޻���?����8�ڜ'�ZS���޿A
�e�?�4.7����9��FP�M�?b �X$3�����s�Zqb�?�2�V����q�|!�G��&������%�SE����?`e��c���hR�h%��u`?��A��)XWL��1�3�*�75��K��d~�g%���S,M8^�D���x��p�)RU�t��,�Z*��l�NbH��r����޽����P�o�+ϕ�V�1_�o.E��C���/�H�{}9H��CN�|�ZC3*�2d<=
�P�!����d�Yk8�߂�A��eY��y����M��_�o#�*�hŧ��N�\7gk�ҟUJ�M#a��}J�H���Je���m���2��Z�]� O���P�j��)7_z9`B��sP�,d$G��9�dQK�w��i�с���e\��w".=P�N;�|����_VEM�3B��_����Vr�֒sqF�/�8yop*E
t��x/���3q���9��H=�ߨ��gTnI��̋�#��- ��H�e�!�
L�b��rp�s��'���񥖡k��皝��	'`صχ��{|a���y����(���c86xe-9Gb�W��~� ��,nXj��ݘR��S>�PH�#��8��h�(8*��*W,�IV��Dy��q�E���j�����$�*���Ԏ�8�[hF��G®�ʷǅ���.�ןt�mKh��B��:N�v���/h͛�����lʨq�6�Q��X�T�e��AW<x�T�!����*7$�}�K,'2��0��sY��`��X�H,˥�;R/�wou�MB�N�������_v��Q�=tDJ�F`��*��(��'r�G����+bN��p��f�9d������'��I��}��������}�׫��+`\�t���|l�G�=�,�8X�e蟜���ugD��.w���2.H��E?Il�����^�c[r�������O�j���z}'�B"�b56s���UE����WN��p�dE��tW׋�92����X���F�����<ko��
85�r�zM/��8�N��h��VcNӚ?cZ[7Q�B5/k"����R���u����!��G��5�����gyuu3h���2^`e7a���И'�ףO;l�oob�zt10Uל�q�R�]��Xl���:����A��F )� ��9�bxQ�;��?�u�Q[a>�l(�G6��.��'�N?�z�H3#�������o��b�.0��Q��En	��ӄ]�3% �m��Pz��Jx{v��`�4�ء��g�^Qu�����2=�NT�P=0<hk�ѼU�����P?��{<��Z��]���R��''��SYR�ɲg�w����Ƃ��
�������²��7	�S�aY'��X(Dˇ�_��
��T��u�P���#҄��óg�z�#��U@<��q�wq���F����'��{&��y�M�C}�R����ਕ?0N�qԳ)?mM�D7$�N
�Om��ɃV]���J��@��rI��ۗ+��B�Ꟙb����bW�t�Bn��u[U����yҲ)�uT R�W��*)x�1����&�.�o���{�j�����;>fm\as
�"����	�U�`B� ˽Ȱ˶�ւ���pw��͎�ُ��.�)�>���:.����y�apq�5����Qy���v���o�[=�`*�Y��%f���i�	����qW�n�͑+3'��Lsm���sw�Cѿߌ��	:��\FCڷ>ޡԞ����s=�����>ʋD�Xޫ-B�C�����I�j�sa�Fk����q#'TPE�?5��5�x}��t�-c6~�m 5"c浿v_�����x�8�zz�����5�ͪ���@��f�]#��<�[[	W�ig���>�"���������w���O,��o�}dq�֡��"��K�����0�@s�m�a&�t�^���@C��ڡ���bb
�:� l>�p�Q��#�5E�)�5�k�([,�qe	���'��*>��g�ul�{W��F���΄E{���ּDlO��l�,�Z��Rx�+Ԡ���c����SEEy����L�����S&�sZD�j����b������EA���v���*[�8X�8F(O9��go�+�䱼���e-�,���|`{d�R��j���KF���e�y�PV:,�R/�_�N1JħQ�WY�'>"����my ~��vQ�٥C�Z2P�ό��z��Y(0
�� $������y,w���O�er�֒I!��N��S�.���"���:k�.�ǡ�����uy��r'��Ys݄��������������a�yŜ6 "yw�5&�18 ���;'H�Ѫ�X�Z+�S(����o޲Zl�u���4�zbW��'�.ބ���Ǧ��Kj����A赉2
��)D�u���&��c��ٲ���:���C����A�X/��4�8�z�ɲbY�|���^Cc��#���/�����{T0�lWҀ����d����z�`_Q6��w�(�AbẔ=�f8=8SK�R
>�c��H{ςJ��	BTa"ɟ�͠X~�C�N
��v��qx�hu�F��S/�O�c�|{�|n����dz=�F���S��� I�Ihm2v���4�J\����F�?�R�<U9,��:
��U[EQ]1��y<�����Uĝ1E����"�,�d�z!"J෶�Ę�����/K�oa��o��c�HIz!e�G�7Q�<ъ��h�mֺ��?�f�p9�����i?�07uF�g�2�
�>��EFH���E���ʐ�^�5�f_�~*�b�<ص���OR/9���@q��\A *�:r�.M�n��4��&q�������Jn��K�����ҞL�/�N�1u�Ν�;��x���T�T{�d� ��=|����8��ֆ��w���ޗg|�{���=�m��^�/a	`G?��"0j��* ��;>�0Ek���Y8�L�����ޜ�
-d{���>��k�oTKN��bͺ�y�c^]�ץQ%�����3�MfL�5��
�?N�h�1�<�Uah�ߒ+��Sƪ�ݷ�e���=�׶����^C���V0cG�2e���yp��S������%��������E���/��VO�v$L�^��l�N����)�i��Q����˘����c`�?XwL5Y,� ��uލ�"ѫGpϜ�s&՟�9xJ���?��86�5'���X3Sx�-�,`�6N���j�:l���]̈́4o�p^��137|M��]jV��P��ҽ%�
kՓq�0�c}��*;8J!��喵:=pJF7����x0n�C6�����G^qp�ط8ݳ����,;}�	ÍOD璲qP��y�q˄�`���R����V�݄�'Ԧ���K�S�r(v��Z���W�(k���r%x�` _��U}۰�Iș�gu�[�R�X�!�3A�,j4�D�������̏Q`ųs�1��XBWv4�"G� u=����>�� c{���W���@ڔ"�e��E�m�<��0���ZԜ2Z�ϳg[wm ۿ�>��Q�BD�{�J�r�ے��zny��˜+�0��i�a��d�S��'�f9�����Lı�\;]�@�RI�1³�Q��0����W25��w�خT�G�v���cal@�"_���#p#
FzM��*AT�p�.W������=^�u"m����8�I	���X�n��q�V�������6�-�#�{ ��+>���vơ���F-HYԘ�>nJO�����0wM1�ERG:f��sr9�������e�ܦ�d�4��:�L��x� �=�;݌0��������+��"IS����bI�a'�59�.�	����R=�~$�C^a�{�gN���x;�B2(>�ař`�0X���c�FR֬�&��(�2u�
����.�X���d޲�?8�q���~��(���1� Y�:Z��-���c69ׂ�Կ̏�	�}z�f�!���s����|bۦ�x��=k
�Q�(���bEWΣh<$9�'i��|P	��"����F��
��m��8��'1��-#��67E/�f�y'�b�&#Tx��~�!��AXy��۴N�*�[}-�������\xji��C�㢘�.�r@�N�\�k�'m�7���4������P�����ꇁ�ηyY�Qɢ����E7�8��P��1%	)�T����@\8JF7��K��|f`bge6���\z��y�}��g�%1����_>�"�)�<���\���M�����˦:T�?��Y�b?{����"�j�E���0����Dm�	<�'g��w��"���{v�7L��F?��,B�N)�	�a�����C	Ie�,݂^T��}��U'Z˂��d���S�pg�3�GW�n9�Z��Q�^��>�\c'w���ӳ�d��X�x�� ��w�k������ qt}#r9d�F��r��0�
K��Q�����LL�hLI�@k@U���D1�̙��{�Hk��V̥��2<�0�ha�c�"�s���V�����:�4=�s�~͵���"m[|��:����z�ӊ��z�<@ie�&�������D�q>�����e�&�̎��+<[�b1�����ey��#5�ɠfǆCW�� ��<����c�4�����^xp������ݸ)���yɗ�IO�tof� )�WG<�d'5�/�༶{&R�p��Z�'��,D�9M�ѥf�����d���s�]��Zާ;ϡJ�n:T.j}5\�C�`r�7T`B�c�\G���c�U�����0�k��u���-�A� E$���,���ߡ�+*���_o�H	xy��}��H۹/kߖD.얅D��'c�:��Ez�~v..�Ƴ�ݹ�2K+�H�m�+^��L'����*�J�o:/���)z�T��������r%�W�y�d*���9��޸n�T�m<������M�Rr����5L���]�Դ7El��9:Ƃ7�c�.��������[ꉋy'f���.��ʣ��(��Mr[�V�cJ��ry"h~8���7T4 s��Ԉ�;Jz]5u��@@;�u��UM�х�܉� 1�3�&����zP���&Tl�g��]�����_��^�{�G@.'�?���*t�ۃ��,�^K�g�i�"� ��u3�L��x�9���14�\?D;ڎ������L���G=�w�0]~U�L;�����l���x�v�@~'Y.�G�����z'j�\���5�c@?������H�)�2-���O|RJ�:��KZq޵��w�l�䋒9����B�a�'~����W��מ����O#bӥ�$2���y� ���,�YJg^����p��A�S�Ϟ]��\N�E��޸�]ܤ·Zr�ʈK?�� l��Mo,Y�¸� N�۔sh�8P�,�x�AY�_U�����@ >�����ow.�I��;�P�0U||Nl=�T���ɔ�Z%k�4�3��el���&��m���?�Ao��n����WKd�q@�"�x��z]��QǦ�,��ݛ~<�j�vKF%�����{Jȥ�4F2�:�d>�ȏUnȌJsϾvP�S�(F��X	��ps	9��T�;��������j2���I���EJ�4�m�stufQl.Y�;j��X��'�M��8�W�|{�蓑���;#��C�E�,����ml)23��7Ak��w�wcj�����$��eQ�z�m��-����f��:�����}��\��Gy�'��	��gZl9{�yڰ��q���m؉��*�O��)��[,b�ՠ��������$t��܃_-T;�\�����?[����1j�r�$��s3��ˆ������;��0��n�RNN|����9@*�&���,/7��RI�s�L����ݲ����hC�(��,|��>%���/Up�A�������	��͇���h�S�:#ŨY��
��!��Ej\g�p/������U�PT�p����<��L�,�y5�I�Hȏ�!g�~)�|G`�j�ځa����!��M�E�`�<=�����j�KB>|>�^��k>|�\�*&f����y��FR�>k�,��/m̾��~��d����y5W>�+UxY���'�)�a�=��{��w�~����;�������ӧ�;�3���g���I!��`�'1�\AZ���!��X��Ț-Jr�7��`��a���^N�*9��R�J��L^�ЕS���2T]XδV�t�a
eڡ�+�S�|s��Ձԭb��a�oк_�=�u(�py�eqG��(b�C�m��ou	�9�vچ|�ʟ����z��h�L�:���)�-|i���>Ƶi#�l�8KE
/�\�N[d�^�Ǩ�Aʯ�I�{�w?�+D�+/��;����7��pՑM�� %����������>�
%Mp�Zt4�H6�Ct��Q0��Nu �G(ut���;��;��=r�z�x4�ص���ҊX< 1h$!&�׮�g���8���!��B'�N�,	b�Хx��k%X˛��� d���C��.������8��eA���V�<_�rَ����C��x�#x�"�?�}E$_�T�%q-���ӳX��s��˟�m�g��B����&`�l<�����I&��牄[�<���^���
;9׶�[�k����;�%�X�>�b��������kV�vwD�-�M��Wp�sb0!\�+��;��'o#��	t���R�|��]��*7B�d��]�ߧVh�^�d�d�I��~_�P�X������j:��Iܺi��IW��R�h����|��Q3�J����H��8�F6��Q��v�G+��[�\�Ǣ^�&B���ƻ	^d���;oX�`-�����3�� ��
��@��{�E��)(�?ٙP�&��ˬ��OK��r�셂�x�%�W���,�^K\8����/��7�f��۫�P4=ܘ����O.�k�>e�z�>.���c2'q���*0��X�>��HW��k[�^�H���'�����^��፾�搾�&�������bePV�Rs倪�(�QK�����l�޶X	�ҝD.ϓe-2doA�D_�e���1Kb~�u*�Qly�
�.2YB��9D��	���_����������_�폹�q���~I*^W$�&^[��#��I.�Y�q�}p<���`�]��;���# 
`Q�tG��p]d��|(�:}��&�n	�0ՋW{5=~�uW{��7qb+[���1��z�S?��48�\�/������ϳV\�9n��Gy��%�t�坴�h�Z}<D-/b�r���0"gZ,�(0W y�v�AlimI�q�O�C2<��l������Yp��ȧ� ���9����F	T^�uT�ЍZ Q�/u��!E��� ��0��ؕ���udc�����%3c4�@Dj�+�nt�C��:iyտ��Z1�;��{c��B>�p��t��.~@bhr<���b|�D*J�!<8֓�D@&�a1��d_��H""B��ITA�7h�s����@^W�)��:����U������<���=�@h]��bn��eT�e��9�w��m�떎���oa�a�'6�k6ѵV��ro;3S�$����a�CH�w��x	��+ԓלdfݳ��]t�(nj��$�e�%+��� >m���6���А5(�S�Qܟ��k��6�m�[V��$ȁш���ƇE������N�(b�xXp)u�L��Qv����G$�?Ue�#��3S^�ks�	C�M,�c��2��C������S	o&E��i��T0�<"{x��9F�~J�g9+$k9�C�� �v�n䍒#"ڪ��X��t��$�iJ�	���G��ܖx㶔&�C,�I&��\�:Yr�^Q�d��j	s`]�a�i/Y~i~tkcK����~���ʣ�AYλ||���$��]H��D������F%���Tv����7�9|�k�)I�g.����$l���(T����T���X�)�����d`�L����~��F��YEՅ�K_��MC^�������Sܳ�F�]є=��p���D ��2ڀA@=	w�*V�=4(ۗ�����ǟ�L��_F�Ѱ*��+�!l<��Qb����չ�K����1��1�cCCF�Z�WmǇ��p6��_�K�a�)�@xo�s=\��<�6���ijk��^ ̽����ڤ��������݄㩯�������ۼB���_�u�l���ٮ(ݥ�gw��%.T:�;�<�ȇt�b�s��/��H,�һ�� ���z�g��L)v���k�9X��z��Cm���hz�	��ݰ$2�����^d̆K��� mA��B�����m�&�?�FmK�t�6����=.�̀�ua�:J���DÀ.��[Q�7��b�R��L �緮 |����\0X?$H�%ڄ�%!���Q Vxk����G��pU/�Ú98<�3z�X9.���'� sh-2&�}'��n�X�m�D��� ݃�@���BV��`��T!�G���?�Ǿ���q���&�O}y[o%�uJ�X��ސ��·ڂe���a����K:��P�}ܖ�fg6ZQ�Z�"�W�8��!�<�⏌�R�_����y�z�j5%�b>N��	��z,X��U��k���A���T���գ��{P4�[�+�r��9�M�ϸb����`�����s��
�\g3nG"��jt�e�D'��"�"��=x��Z�W��YSg������C�J���h:�|��WW�cr�(a�J/H�=i�.���.�C��pbC��7VV���[(Nל�q�������R�zᭉ�eR�9��4=2,
RȦv������;vQr�-�쁙�F��/9�P�?�w*�t�OP<��}��n���0$Թ�z��T�1�h�f�
� Y���m���aU�Z�M$�E��������
�M柃i�Z'v�����+�b�)�l@0XX8�A��*�0�j�K�fe�j(���4/�T~�M����/��ɶ*@�(��<��߅���N���bA^�����a�S�[L����xp(�-MC}�_�E� ��[X9��^E>�?n���d��c�\X7O��a[F{y;����|Ri��_M�����:I1��/�����;�������)�}�Rl+Gz�^)�&��Ik0�loOV�Js^��Vx���O3�x��%6�%�S����ȦMt�h��f�M��z�D�ZtMY�^wt�绿}�ˀ�+�8�,��%x@���zG��.b#�%�b�TWR�:�ީ
�5����qﴪu����o)b�J
����s���ѓj3B�5��8z�u��ab�6=E�����$2��u��\E�D�W�Y�	Ik})�q�����Ŝ_�����$��]ы���#e;#�CY�w���/��6L��yoɊ�Ey���]9Z��c���L��K�}p�>֡W&L�z$�"�M�M.G	�{���@��:=Q[ˑ�+KS�'���=�:\���w�E`P��Xļ�=��D�"���v
c� ����]�`��C>N�H���y����u��!=�.�o�e�i�Y@�x莴 ��ڗ��h��Hy�:"�n]?"n����8���ږ��Q�Үj�%<��k/�^�&^c�<�)���4��fzVa���sU�=�RPZ��'�R��0 B��(d�-����ۥ�:P��Q���}��q�Z�b3���~�����'I�� z��;*w�X3�������s��B<QLC�0:�%[\���ŋ:A�nKJ�����
��c��92R1�u�F�2�	b\���t����X{:&"[�f꺤�F�5�f��G���B�f���"y�
��`��2�A�r�O�H��vW5I�4�7��qH�[a!��l������1�O
A���h�U��c����z�H"�	P]٦7!��A�	'־��z�^�>�՝�*#6 ������7�:2Qgg$�d����?�K�[M��3ƾ�E�G�A�Z!�(B8@�w0��v�^�4�Q���G�V=ZE���m����yu��ྯ]�ț�s^��&$�|����܂14$%!�,)��A=34�̃r�"�؞�5�l��B�2yM?!Qڿ���0�{��ѐwյ`0 �3c~R�������ىsx�'�^>Wd�A����;&�rk/���2J4_�W�js�L����q�a9� X\h/o:u�V(��>%hhN3mXl6j���%�׀u��|����Xʎ����@��LS����^t-�&��6�Aޭ5wft]��TUO[���]�GJ��26\/FMGU-Q$a�ݵ�$?�Jc���L������vc�2�� ˗��	7�
R���	u�=�vk&�fC�?8�Տډ��7Ɔ�&����.�˅���7���Ev��l�#-u�a�>�u�k��a�L���7�t4ܖc�jrM�N"�GA8J��~a�� ƪVK�����x�|���<��\r-��S8K'Wb��zvr44�T���X�z���d�h��B���&LN�5 ڬֺ��G-z���#�"O����D��o�vU߼��"��7���Ng�m��rtV�����E��z�4F�%��t�O
V��WsA����C�y�Z�g ��eL�ݼv��u��a���u��醐���VGY!X���H�G���#,���/�M"�ӗ�侀5G�������0!�f������;pP-�<�_�1�1H�<�k�J1�. �:H��9�d�زbiu2䊗�uJ�(�D�d��&�},-B�nڣ����FO��ۥp#i��aU�[��p���
@�>^���Z�9=0k�7Y�auR��6�sڬ�}G5,�.�sh��0/������&���f?
��e��,�?�Ɖ:�Qҋs��۞��Լ��oS�	��8�tE����Ң�Q�zU3q$��Bz4�R�k9�����f9��l�H��0�������تY38��k'~+�K�"wި��aڎxC�C��7��o���`O�2VDI�C��Y6��Z� p|�Ⳃ�{Ewd4��Fkbi;�9�UZ ����q�oY�dp��!lP�iH�1�vz>H�)��<�1F^��pH�x,��8�'
�PE��m�>¾��rsyp-��'u�a�ʫb�6�����