��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�APq�lG!���h��2�&�M�N�5�cµ&�z[հp�F�/s��2���, ټc4[Ӭ���c'r+�f���W�fo�N�?�z;��O�UP�D����#�3�R"��Y1e�!����W����T\�ۥ����-��5CGLI]����S
��oz��~�d韲T8O�Ç��Y�ld�k<q���4��TR���۫,�P����Z�`��xb�X�J��`�㱻\�����4X�����rl���sM�D��ߍ[��Òv ΐ����s�}׀�G14�J�9�@��Ӣ-C�ʖ���siT~�@�6WJѩY�|mCC�ϙ}]G�N$�e�,Uc�7�H����S_��i��:��G�}p�.5�OQ�&��lao �D�3�e[b�����U?+2r�`�د˴%����9$e�4ƻ���Q�ZI�ڹ")�s��2y�=��f�h.�!TR�X�佔Z�Vp�S�r�)4� �&����{�b����H��vc5�T��u\��9�E�ڝO"�:���^HGM��o��@!?7-�"��oˮUǙv5�|�&�4�c򪲤73�Ɖ��BT�V�������`1<����M��z΢,Q�-K��?���2�=!=�;�()�7ig�1]�4L�h'���-����㱮�
	�w�� ���V��
��Hf���*�XN
��g�]ʩ?�m�;��,.�(����'�Ө�_�p�j�5S��:���l-�+�+UY<a��s��`��Ҙ����̗/?0>�[��!�2 tv������L}�+_�WܔD����.���)��X����*�yW>�����\G�<�d�����k��%���>����2]��"ka���c�yOܪ7�$���E^ !�s�����B��#i~^:R\��ޕ�л�3��D����P�����D�v�$�~�I���
�wo��l%�z�*6k)+��
&�F��H�$y<�6~���Rs�Bl��K�ӣ�\i���\�Z��{��+!�F�0+��Hֆ�o�C�������!H�/��Ӵ^ji����OJ;�5����HL�k5ړ���*5�-�杀���:��\[h{�W��,�ɱZ8v�zf��M0W�ɞ�)��T鉭e����c�ׇ�#f���+�rȀ�a�]�H�k� аL L��V���զ'.ؼ`%%�e(Hfod!�?z�i�˫S(������ "G)��q��[=���(��o�\�d��|�թ����	/	�l4B�Nw�,1���i}� T���Z,`iAj'���u +H�SG�5̱�>Z�w�?!#j�ǚG�pj���v�e2���xC�������j?!�`ݏ�E�@�U��i ���B릆�1��R%�\�,W	wL�HH���V��|���m�P�`;{x�l,}6�(A��Ń�Ƭ�)�A�]Ba�?Ʉ�b$�/���O�y��h謗��1�!��`�L�b�Ё(2+�mL�>5,>s��tKzFGY�*�4>���ƙ�	`�ؾBQt�<JMc��#��kɌ��扫�z4�(*Ϡ|\��y�����Igq����I�?�.���'>��p�@��}g���N� �%�(S�؆s��b��%��+���/ ��_��I�v輕!��3' G�F�k��l���O?�Π4Ψ3��~���1bU_�We����9��D���KU-/�M�����}%�X8T"����!ݤQ7\Bո y��Hq�������dAI�Mě@��g���@��^�;22c_ �h��#OL��0��a���a�Dv&<P}��������JY\9���/�|�H��M�.���N��/E�yJ���Cݬ�p�i��S{Cb� �:֎*�4�ԑ�3{y��V���v�r��&I.�t(䍆9��C�����m�5B�k99��o�7������W�)�Ѱ�V��������_ND�X0>8gV�,��7d��n�D-�-J���נ�A͡l�.oQ�����mYC��+F$��] ��;x�C�֌��
��=��~4���"��%Q�=�F9�y\�8ݖ�>��ҡ���D��	����S# �4�}8Yؾc�z P�v�1��͑�2�O	y7\U�E��bR\�؈�������?	WR"̉I���N�籁�����-�E���H���},a���䮻����+yZT*���A��x����d<bjL_�k@�rc��M�U����5���UT��Y��^�w��
��6���gȅ��LR�Wd�8��cyGK����y�S_t���������(A�:����你�aFAF��Ȼ,�w���3����!(�����)Vm�m�v�셲fX���l��3ϊ�� ��I�M����ds�`}��`$�=c