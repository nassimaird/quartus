// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
W4FTCOOJnaBR9qHddAcPX58wcJFPYHVtyyLyzxQINy1kTtE+K/je2KuxKJg6xA9fTU3GrNLT7DcJ
j9IComigAuySDKD5w5nCNIEaBGzgK/Tg2BJsfcL5d6HWqlV9dfIPgBMV8sMm4DUCigjsyq4qInfu
ikWaoFdUGipNjE+8vY6P5oUoDDPp7PyuhkNFthHZRzokO8E55F7ztHkBY8FfLrQVQAEjlf4e3cf1
9m82nPFiMBVcSodK67q6b992QYiyMfO01/gZMaxx604mpZtri73lYP7hE8ilZCl729ACIshQ/1UA
me1v8Z8Rz8HfUFt/+3xC+KaPaDJf40Nqyf+HxA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 46672)
GL3jKdBiEXCwrhi6/uiYwDhqOtRh6m0JonauvU09J/hTFPYpAR9Lgppg0t455fK3WNdvPtrzsNBG
VUlEhrwlqGtyhg5jJzoNTdeKJ+6iqi/NWObf6HHsNvqeRQ2F/ZL/jioV8es6Duq76OFWurbAgxQJ
EenqO7VUkdLtLj6LizbINZkfMkF3QFTpXiZC2cZg74qw8mett3LPf9vOlk1KL7TBCR2NXWDY6wlU
c5CZZDoe8YwxOpF9yyf/1fH4MOuCaCFyTiOav2Gf1/Lli4S9TxwjMXAbDF3SSj4XTOiuRaLp+3D8
hITwXHJ7U6N44vVM/uDrRhu08GCLkL3ZCr0LahZQnDdWbv/90gVrBbdEwqnqul9UVqbBiTX8eCkX
5Xz2hXUObqOA475chHt2meJyGaueY/d7tuymr+6p4O/lXqMngWCcSKIi+oe/CV8ixQMvJepxnQzE
2HS0B/vwJWmJejS+xz6lnIryXth1iBAeSDKRb2Oeksag07/84wvac1jiNK/e+oUGcO3/qfztNJgb
2Ou6liydslGdpmg+FbuR7e41g5CzfgEjNcHlpX6r3DQCZ/uJcWxWJ0/n9BZZfrNdkEniMKCWOn2u
l1qzl1YPvejUqrFDzFNKkGymCEvUTxrc8vMJBSDnrL4CPKKvZGq3wJ1R5+6/ki/p7FJWEmhfh8bO
BfFqijudsBZHkJul/aDb8ZGlcJMPAlj6vviw4ZptUJLWkBlWUB6hAl0zmrA4Skl0+L1vGN54LG+x
Ve7ZC2ysriqEjPQxd7y2acQfyDjxkjTdpBX8j7JYyUN3gYNEZ9EvMI5h0vePifZAGnVq0xlx4mDp
la4zJYUDRbGWNGOYHnvYOm4q1N3xJiUf3mUBbpFhfucybF4ET+B/cANgTBB/d2tKYSxev5fPzVCb
embSGP+TR56L++adIgh0RSdegpaUnEx4ew7BjT8dykKMJhC/LbqAHr9M3whEjPpISb7oz1d19+Af
5eG01PMDq0DNCinF2hwJfbwKoGgcB6QU+6F7P7wvUI1v/Hk0aNeY8UgOLXCkZSyHxMKfPjpdhDIu
mY62NBUUSCR6gbFMCgB9gCOvjTBvPxapHI0yMbaB29FMCJafhh2QKqAzfUot9Y8UtsIsRdAA6nJq
XQdvrALKs6bVBGy5B25eNA7vkvVDPx3oqrUHEx/+2oMMnNlml8r/BbP+0cKUjvDOS+rODnopU4Sx
B4ncici+7zvQIT0zCpuwyGd7j+0nyNsPH0vQVm1s54pxWXh9hAlhxH2HjSVGS1OYbvLpVPLwOP8C
N4l8axADIo/rGe18iPwTr3eWVMAYGUptaiwee8pEZtiF0/gpledCSl22feRYsQ5pl83zBHuoaBsI
BHTMgOaZgp+gSNe/dHAQDCQvR9adM43M7hg9jHVcforSNE0kqsI6XmhhvsP7f0yZ7rnFoxtzBjbr
GFdHlgq9JsXmrb2QtVEOA6IwbWN3AevcM/DlWxTl40SfwFe3Ft7H5/fGFHH1Q6R5CAT7Uxe2T7I7
OgYAfO+etKLsbeh74gxFeNtuO4j4v2bLW3LCk5zriPoy1sf3BjfYATpxCzjvSPjq4t5hchtnphSX
3Yppbl1UzZxprYDwKxWCvldui7pgTrh4WRS+qJUf18anWMunhpqoT7LMkh7+Td3FFIGWhBjQGZ/A
xl46lHukC6ky/f16nKBha8ZYmdTblXQy7S439BA2jDgMS41xz4LEF0/5SuUyfsA2003kF8UJDVok
YXKLyRnLimjsiKjEjNxq/0kDmGPV/5j6NmwbTaaSuLre+NhBXFbUTv3AEBy/RfVgMMid0e+xl89I
8ffJlM3e9C+Z5NO6EGmq1QvBJr/ZhqMu56Ltl5c9N20EQA/SrU5r2y97RUGfLKeJ4NibRc+tbTSD
pvXyItfdUeePxY1zUh9+3b+oq5GpXhNvAjeM2TO691NSh8g7TlZ/23Q+6wedYeRzuGvPZvxnYSVt
MRdh0EkP0jKCdJRJ8J9Q50LtFVAG/5dKvUxAY1SZAwgs2BaSSAqf9Swt4IwxUzV4rRuHXdsuRyCf
Ay6+ThIBkPl5v18VJaYktHKbtogFq7NOrAm2baodsO5nokJmZ9P9tuM6XTAkPbNL7R8yfNxpu9SR
OPYJv2NygvEUnBBBtlJ6ei9il7FwlZg4qnRqrl/AZyES9X1lhMuL1zWX9ZHvECi0DpwCh7d0Ks6L
rhSSq6FrlDWOOcBl9h6Pe+HpKX6hlHd6SqQwgcxxmhohvX6QRbXhstpgRgkFH+FedNYbVQGDd5qq
AkVTCHWSARZAlHTsuTyh46dCrFkxqwdJt0fHlCTqbHe7xxMeOMYyGBPmo5Rp8oxpl7DrA8PLDbcq
gWf3dDeBn7jmiF8/ytGbIiS2IE+EHy7gXqHZuRr+ba7b91rpEiqGLDNtxWZIEslcyekpfk2Ba/FF
ow0nc3btBIV3ZPFfZIuSUrpBw5L1CESsXquw5dErZDjrCruZyeum54yJ577/2EYId3IJQl2HhZ+w
6mmdx9jmMPi7X8AdZxgcR3qRAGq9RRUTcDMTi4YsLgn8XIEUujltnmClHnpHvZfCoBOWYPqgTpGC
8W8BDazQIQIeQnhYNI5YbzpFukLufJejf1BmbgdKTSo5uFClEOeCffiSAYfnLkLxfwnK+2JU5lgc
NrlaDc7KC0wQNKIzQKYd47e4WgEJIysb05TVMkyg4s7O1PUJqs1NdNiw9KkCkWe+tPJnXBZ0wFSx
SnG5sXP6/R0gyigMZTrOuf5FTPwbadbyjpUN+4QR0b95iZaZ6YMGbeZubVUGgwCUsJ41zCKD3V6m
gi0vdNazwYvM24jDkSt8XcFMJ9FrAMqhcY9Uz7hd/zsxQNoyh1BPyJiGhc+AJAaiKE/yaL1KWo13
g6mLwa/rxiumY3wemiThvht54qXV2jLKZ0YNCdf3JoqLu3ZvUmeUbDz3SsPeUiRKiGT1M/RxEU90
pz/zjRbR3OCT0xL/5WhWmBtSYHMXoLmRs4gCMzSDCciVIV3jmdpmKUFlqvIFfznJ1Zq9OdjBAsbX
PEaxih0t9FRiwIQ8R35M+JuzO1NyQpu5iqTkuoM19Oqg4MIXOMFPcTQIl6SJSGqXZ+psmnwIR8ZP
ABHrK0i7uRhCQBqgJX9q/YS4tRtHy2P9vcAQ8FamJYbnL6yebpH4ZxxY6qPWksR79ePJeOx1QM2R
q55jiI2Fl26iRDtDWwbWY+1/PMGvnKGfIgHUm9MR8LBlwZ+KqIsg3DCLLaNzJxUOAN018ZTMRTWk
A1skE08i2+AmLC82EsFqIil+oDf8cAR0u4UBWcr4DQcwTgnJm97Rvxyf7M5iRqgMtcUvIGva2pw7
MaZ5IBoZkSKZAz4vkNGwgl+XxG8/m0+3ulzDvSQs4Zb32KJJHEF8wngUSkCuK01JkciViEEmknHH
N64pilDVSji+pWQjmS/DnBqfrj7NfG1Kux9DITy53oUGi+bjliLAEicMt1TLVwqglevwQHF7BaH2
dljjkfIIXzxH5NqxW9+hIbihXoP8Z5b8bK6MEcYGEvIUQf7YAzr++iioQm49wzIX9m4YKabk7yxG
JZHowi5nojMIxKH83ojDXg6vgYSi1j7lVEWNIS3kN4IKfp90QtgGUsoeb/2OW2rCf7Tz4uqfX3vb
eLmQ4Q/uNdqHUNZow4BVARuQg2ts01NSEVSybuRk7i+0N/vhylPsEkheFLDL11WjdaOY22NRUME9
OfOBYRFM2zY2l87txZLOPvW/gDFAmgVx2U3hJSHlOnQwiPIKoXAcyFniEu1WCckVh9Mz08lc4UTU
BQX1nCyFjPkhlwE/BNIV7XfmuYNb2rAVX3Q/H9dxgalnSJe3YczS4q1egTxqmhkoU4Jjs37oa7/5
Ad6GzKSAx7Y3YdZAt2plg11vsLwpIBWrxF7eDjsRi5zAEHInNJLWLmVpVqxudwdGCOEBf8fCzva7
DYLmIJkveEYo5HljcsJbCGf1r6PAa0GuI7KxtnP2KLngfvw4JNSdPOyuF9KiYWtVgK5VzNEK/nKS
VKqs+S9WknxVWIuxKMSjXR3VNy1Kr4p63yBxRBY/BQUUcKVKgmvdninva5/uqC43tb0XmhIsVofb
9Ve3AdE/YK6yeQd6xHTDTAumH3+X8/rhR6AeJajqu/uEZ+AwWHrdcfxIS3N6IkF8+d5Fja25wvnx
/E9CvBy8DO3PXGcQHAgI906eJX3M42+/Oao4dLhYpNJc/OBgA791C0G9V7NmykNXOKjvOh4anfZY
0yINABojYtPEfTTZAxzpGzIqsuNlU1hOfx/Eubqvrb7Hz5fKjcmQzg7KCtKIKySbBexNQSKS756T
s5oFCca2NltTq2KpojX3kwZSIuqYiNdMG0JkkSs5QxrhwVuHrrq9Zve2aEc/mVZ8PlDTTTCOos6V
xcGYtP3ddRzcD92Bjhk4/5O6TjcFrXXhTbKIJ+6FJq0iqXxFH27B6CV7gFAA2m3o0Xbzy0seoYfi
eaGv1RPMTctRumtFkv6FiG5SoiNZFQS4haFbL3XWxnjQsy04hbkyWNVSAiMM+jtXsUMYdvtIUWGr
3SYgsyfzYfFmWqKrHumsPkTB5VXjqPQVFeoOrYe/LQEqlJV6hfa4c94nN0QR1cHIOHQHRfr8/cL/
WvBzCWBdWH4HqUJck1ErySWdccgm0r9QRDMp5QLYXaUgOYHYVUj904odxm4RdeD1sDHUbvwN97Hw
FNq4At+BiNfIJRTmu8EoOXW2A+OxA9/PQkjtN1WJWFdh0F/4LRxY4wmiJrji/n3JHLEZJRQFKdfw
8+86kEl9uNzXb3MwTfSAd8OLVtwqM2Kth3PPOTNU1q9e9ha+SHZQ+cmgGt9NPfX6jZPO5BJJp+Kr
gpgZYwe5KDRBn6Ej9JfWoZb5OUUk1eJZ95KFD6J+qkF7+wKgKbDplPBCY31hmOFaZEd5e4Pyf1uU
nkdFIhiEQdm7946Nu0X3omCWw87lYNeYNN9z6VjbMLC+VdSAoFN7gjCbnnqaBNR/T2VA9SkJ4aYt
snHDc1OYD9xRurMZ8u9vetgNNiTNFZ0rCv7WeHLuL0URRkJJwvsHP4RhCGoxtofxwEk0m/mC8onM
iGrp+1wpLokncL6kD4P/KS2z38k67lOEXDQKLmjETweU+AkXsTQEER6+1UPJcBbWItbrB+aNxxhw
o1mcHDY463MaWaqrMXCoiAGssYqWLFswbAjk1Iynim9TpyWuuT6hDBxkZSa08irwwcjetaEudFOL
ZhgpE+b5LXGG/1SykNPeiB2uTR0mGPiXoRWMpMs7FZdtK3AedPqxavhgO2IGakcOp8KKWopG2RE1
aUKFMq+fIKyQ/PugyTrhSlS8BklylFFZMdFSTKMt1JLec+qm3fpjr1IzcDHVNAeNOQYwSL9/DCc9
7eki0fn6r2C/hQXmcjjG3xgU5zmJ7M/nfKDsV9PmIyEHGk5r+HFBN/VfuZp5GtekMP8fpdGB8Z3d
yMMm9eUPRbBF7vp51JhXd7+fEmmxQgFWmw/EEUQ/MZ80f1XSEq+9D2Wbwtr/985uWzFQvgPzOEcS
hVH+X2frX8wX/acsI4zDHOhCADeWt/HmNyyGyWBQImsISYZrqXjpmivrOV4I2ObL8EtQkugs/C4y
ZLr2CcjRxcc3QhtudsvhGSbBEXKrgVjv8b6/LqPLBIRE6fpTvCS22pWOCnw4Amhhc3a80GC0KCfL
1rwaLNyNKwuOP1smWiU+71JjxPI/uwZMpWCOSbhs4j/zegjev956AmSiUX10zpfAxZ+UT/s2FRCt
EhkpSpG6Ezi57UbUun/LBLteQd6wVjTEpckjTOHPDgASE9IArFbhGZWPJVRAWQmJZWGcTGMI1+V3
KdzwQDYNqGDqCZq8sKRc3+p76iAzGKjjX27JSjr+0s0xP2Hh1N5XXxkTn+gyRZzNOX1cJDzQHwG5
LfyUnLnSL5kGAR06ty94at7ASfGtmTeQVjfp9YMtH1Om7k3h2QrP1veNf6hVbsgOG/vig9QpE56Z
vR4j3M1EYn7GXRG6+K9UMi6qemmLxnl/enC4AMzz2Enqa/fJYntkuGIziWEvyFgXiypDOPpj7FFq
bjvaxqFqPCp600DKdR+fCT5zEwNqdLvCMVONsbgkBdbbeFLt/Z88mmGihMTpiEfuZqZ24HIXTz/8
kqn5WZA8GpN6Lut28L7lAQqo34UusieymMo2XSfVSjrvpq6p96ZKPSZzH0/awZ+5nQqD3zEgQSd/
DsenDjSiM1BKRBFaYzXyYaUz4UH1xdaY/AHk62pizHyyrvjzTbfHac11jViCmDzPQJwoOYinXo/S
Sr5DfxgPKZD6OomTg6Mk1yZFtPsyseYolknooT4IRxhGGQPy87yCDhHcmNkDTb73OuQ6Asm4Idue
kAe9FJC2dTbolqoLgNTBl+RzMn+5hIiqTyW5CS+rPzIE8V+d8E0Nufptin+BdN2LdqQl10ZePmvl
MXh1fwIftn2UkfS2c4Grwt7rPjgW1lVOJbdez02QTfK6v/n6fRinSvmi9EdngMoY4IiwCDM7bATu
sbQDzAqP1FkvbsisP7RQX7RJGUDdrdIgTdB3fGHt/JyQ7ZZQ/KmEDZ+UQseELdUA9sthrWRqAkt0
EavNN0KYfLyDd/EIMnnOO/ylYDJsyrXLcoFYGTEnUX8GFsd73mtwV5h4lh3ijr5Y7EdNTCcfDoob
RW2uj9P7G0w/ryWohyplNnqvhwaXjhDc1qP0odrCRZ4IKylusRy2buaShva4Hc3XEqoJCfBdLw4x
LuFYNNts+Ba1GfUo/OlKHLCC1vRxwAg5+Xmm88zDmujQNQaduy95b80TCkMqws80kUaOuQRzcfCC
2dBYIT5fpKXBK4g5LiqLEsPjC/vBVfEzCDq+kb8fSX4flsBAMA7Wx3kZNAJYrBPIwqFz0kG8iIbJ
aShS76hNNmTUt1rDZctLfhvZ8XOIX1zNjUOkY9IWtobThokccu+WV9B8f/jsiJxiuqXWRI/VeMMu
mi6lJuZNshFTwbQBZgCsaHzoNOiwgGZDDzm2O6m3UUZ/yWe3+Nb8o7EPAfEsiNOaIOI+Na3A5ZSa
pI5+JFQa92OfbBGLsEbKt7IkIfG45JWmxpmUW+ZOG59LdLjXlk1jGrTL6VMRBt3RTmX54z+HZFae
CmFqoC+7cF7sX9cIzdYy8PMCgJzgpUDEZVIe/Y/gFdY8qu5g4dLwajC6uzSzU/N+cAfm3YJckbg1
LzIMw/crjCu2seNyEzo1nWw4GfTO1IeC8uw6ddIILpWdtYck5q+OGyzUy9My4kBMlqscPxKEaNJV
bBFUoAHPwl7F31d3buyUQ0ryP+ZTX0ZV2SZxyv/QsoeusV0W9fedyGsDQE43xMY7vwiOJT+5/w9A
LEQO0+02IGt0FMr+Gv0ADhgksZyrNw1YqJ4hI5ag9GMnQ2IvZiN5xDdfZqcwzrKICc8wtnY5UuF0
oN/CN9/f7Et1fK2mWWES9Joii2M1h3kY/u0Ki2+h9TWiamwf/RmC5INdlRlMQCqKbN6nCxSujC8O
HoHwWvV8QwKbjbWfHL2ppLnK/Uup5BCZJ2LPWiuEyzCL+gb4dynEZ/wISY++1+GeQmUBTfh61mce
jtkD1PnixUUSND8yyX3EAWU1NpEkzk0inFDZTAAgG5ihG60R2qbZGwwkflod8calynnZp0F2WLti
+9YW/2uFVMvkRwve7+Pb99fsI4OIS4gC3WQDJPshtMWLUOmSj6bMxnyXhggbWPwxY3beoIui4hRO
PvjYavMN5ufNe+17toWZ3zA6WMf24CKnYvjjQnz270P3PJNESNC8wbiqZok1AsRPNv7djqjXgM5J
3s9PwX+5exnCTDWjn9/RPGnJfhEqQZzwziwgvD+cQVPGcoRs3IuzDn2nD1eHTwRq/v4lzhujbT0i
tTdEmxlWL47ylwAEF2MF9ei1YacVHLaXrMOt1NbxjgZrz/NY+iSVd7yaH5D55g0rBGWvEiYk2t0C
NV9noqvXsUZbODttimY/xYdgjfxoaLYejduMVpSI6v3oFt74uTY1uRu3IrlkG2Ewr0x82ug8sAmo
HsJmUb5AXiW39gXHZ05mCEKO1B9KA8uEci9FXYTyLHslyvkpzlzwCie5mhVI9cvMmysKa6wFRNxR
MlWPicFh3m8toQlWeGUpt/+yT31LvAqyRTRUEq1lmtsFn52erSUYiEX+FQtDn60/Irie5vS1v3/j
px+vhCiZchsuIlxLLzWpQVuzh6WYKz3lyj67tTZPykAaQ1gsNL5fUh4DhQ1dEqAcRf5ryHcu9Nfl
yomvP2xSoX9LT1975IkKy9HtIiMa3xap6DaEThtzHdkDbvr0g/qNTaaiNzkI8WUuK2YBIDST8Pj0
0GuNc7PSi6KgfKnKXa6w846e8vQRc00xWuKYSCkSqtdZJDZAqiZa7Wwc8h61vyGGGlzbdgwxqIfF
q+j8hnh/dn18cT5xkGCwguy2gqakdBLCEPi2XSAm0t2gRbZA+3jcO30or0sxSHBAYlj0N4P44SZf
KDHvorBOJN0/st1UP5Pe+kCXv4wMnoZyOZVkVVLo4qGSg0irHnL4O/nFOszv5BIP9cg1ErNaQu/r
LB3S2mXtyW57ctfcCHZVfIvo6ATDD5wGAByhq5q/kgeH1M7t+eFS+gdDZHJ/ML8x3VHJl8gYDX97
chzxjl60ubFpkAVE1hd9fClKepEdX9NbzaePnhha5V1vwLqevT5WyTXDVQU1TQDUYDg0HWfjS3KU
bnO0RP05IoJx6adgg2BL9ovGfLByJBwcKsJdpFxEGEd3imYwQOBI8uqI0SKFM0opeLKwQd+0wnxk
RBmh6/j6Am9iuTXBsOalni/DEqvMeHOnncFfcs56Hl9tIRm6wzRIjWUfwPP4XhityR5JBdNrcbOT
fz+SjLWWnX+/XVjZ/Pxi/eRf4UkYnNrcTbXgnJV0WooJjTxyd6GYXhlHwGrZY6B6NOe7KqITPWLd
+kZGsqJIfWPkTXhzjAOP9hMaIv/iy3eQCJEP47y0y3xmPgJiyC+fgJVZpg9Y2sVtIl2T1TsB77nQ
Csh/b3aGP5kQs/HYcbQPHHMtbrbDFoXJXXtcKC9NQrEcB9WFGygD9VyUDPIA//b4XaWvVsxgJGli
ePeOHuMhsjCHoU/7uQgyupRGH508sCBs2SXLyNNURx+oFqk9n0wW0ZdCnREz6ORCDcA2vb1eYoYR
1AFmFyq7PETZ46KjJob3McGO0fWkaQSG5BMf6kQVpPXGDlJ9zibKkWEigncOteFmqucIUmJMy/S1
w2UfoWTFFzoXHCGhgHr0TuyLFH15IAMdJzPGgC+7q5FYJqJXuV0hCKfN35Sjsn8kxQ5DvqvvQ4hI
i5YbXTTuqCkhtlaxrQ9GqGySAukBTpJQ15z6M+070fEU/sO7qqkpOKAWs84+SjnbLeqpbHfcq3YH
iNonyWyd6sTJq5pjyHAk/OB3sbulxS4rCIyYs4v+1mGDHEj/ozRHgTh8SXjDVKvkpHQ/1XHOZGzY
00GpZPT9dC4GQLre8pH8hGH6g2o3l1gf+uZfaLbC/ljL57xm+jum2cL4tTig3wu0P+jNNTQNj3BI
1OFimcClK7CwcgFeP02TcpADSfxv31Mt5NYvmx5gRaoLk1fZ3HO42tU+sgR0KCj3CTlqV1KuyKX0
/OHHGiRdbqF0QCljdIuWOQn9KdCw9q284QCFVeDBpia2OeKF+3hGZF3kKphayW6b/CdwYC3DqgWp
3rBUZN8L1z1GLXxTg0Xx6X02gYH0zrXUp5/A43O2XxVQ0ydJwFROjTLewjTmvUrBDaiImGfyjKGO
N8s17S3/PdsaVzbbUXzXEeOFEsXwkGvlgqTNBgGOJobGwU5s7PfYdxTkNZP0BToUdtma1Ph0vOLV
ugmjRiWYnopgONr19yRP19s7e5WnIvBGCIJ6Ghjj0XPsnbjJiJZvVE7cRulX81W6ALXmigqvbBM9
Q/xFkex7ldsPnl9Sx8nnO/O1tmHyaBMgvtOYWKCOZ4N99iNbaWlP+y5nk56A1NGL+lsVAO7W6DkJ
92LQNUAPQHVGYZPaK8CnE/97Ix2rHe23iTPF44WnLxXgZCnANVr6WYljlH8XYvG8hKTiBzYujPbV
2tG1KzH6MkdCM7seG1U5kKW+WBxyQWYPWumTlS38Rcme0q+3RSSPZFiuw7Wr68yS6z/CTnGr9OZR
R9PUhtJ0V90pndi+nNOTZ45q1ecRizKsYBSpx2jRqi89nddJMf5D3Jn598h3zG4COrJnR9h+QC9P
napVJxpoDTRkFKffuaR/NAtpIhR61OdOrDqQ4AMyXg6v/kmSAoCSKxhUu3wfVMo8jMr1c4Mq6cy5
QsqIYL+/BXNGEF+mzxGFZnyupb/Z3/qi1nD/Atjcs94wINpo/+Xr1Asu6b3Fwy/Av565xSXp4Dx1
NI/lAviWsb+m049PoAh5VmmzInvY7bEneiGevUqiXsJCjEamQ03vP44JZKxfMiGPhpgWA1GvXBao
+NYoCM7ANlxNT/sc+JgV4y43yWSL0UubQvJ7ZFevF1SW8MVKY4F/3YN8l+xr3VaQsAv0OeDKZe3g
xd76uNEB2HVWx46Tb0UHcFzEk98xK8w+kZvJqVVtcX4kX32ZP4Lq2c5xtNJkRWyPETpRycdsVfrv
GZtXK5bIOBmZKf68XoKZX4ToM7O3IWTt2jqNA6R9aM73gZESIKMqE7nKpp3gjalZOvM1bO+vGMwN
QhuSen4KBV3wabDH9va4WZau9sRhiHdcONmQBFD4DPtUBR0aRsr6lz+N9WRH+5lfxa3M/1X/wPa8
MnoA+FVpQwik2L3NNlPt3/7fH/ymTA92DmXQi0LHL9TKZztHGoXVnq/b6RUyMkgi5bVXd7IGzqVR
N2TxHlBeG48vNWFqQ+Feyt+3NcpSJkWmXEtR20dc92q5M0aj1rEVDzZwln7syRfvAmEq5PrHUC9g
DsPgB3VygyXgRljss+7dZs9wEkt8Bu4OlGRPu2ZsqWd4+NgYsvHbTDfHBbf5A+rmNvxwzBoHg2tn
fauyey60snyXYgNSsorZwtvCD5yM7lF0JNtES8CTmN4sravmi38KRvZGyig1HfaZpcUrkgWasUSB
N5QMAW+JfF/djMk1UvpYpS+P5yKLHvflKEyBh45385bZGkRKBmA/WKunwR0ICqkwNHz3REXfOLDG
uyCLAoMHGVKEklWFbAl9hSanmhZlc9UFKxmwKNVmnkObhHmgJCFYojzbPZ7yUKWKCYeBAsLDN7wh
W9Wri1ClIER/k1WMOTUDi0VgyY1GtC4+dw1560SrO+LyfGRSyOsQCQoLvZ8sM7ih+tpzaOb2ao+v
rCmsBWAIKBxjN2T884DethW3MdLJEGERdiSwXC53d4jjiExTcfHFkfTpdcM7DZS43zRzLqfOfvKR
8oNNPbInIGm2+p8sMrFzcDqKo2IuXk96g0y1DWf3sBgD+dsDIjoOds/GCkfLEc3s9T6WIsZmRFKX
oubU0061m4g3NxbQQe5q+7+1xoWGMzWfXp4FNvNVF9NhBTOx8hFLFMabvPfpaqRbC6nkEn8Tg/HR
uEphJ7L0u7GmsK9q5RPrmoGoMxBoAXHOo2lMo3n2G9teCfQ7cSwHZusjbMAhkCm/INlWWg1czd5u
JZ27+9I1e+NfYV/wtNpzkHWzr5xgT1L7fes8hrI1DLFu9WbRxWEXQN4nzOJ010nBRh4LG1TYtIf6
awRJppv6ZuX3ZAE4WRikFA8QudDbKOB+WCZPQm0NwIObFIAMv6DCoRRWcRy2EegrQElq6+7zobXy
7iRkRPjpBqvqMc910H5seTtKIxpUOL3Jz3YrnE3W8sHtb6SRtS5OL36JmpE337lxo1kkCwaYg6pH
sPy5ckm5BSmNGFEDt7tsvQzONNMyELT1NdNSYWasQO9+7aLno4qtrMryVcKntAu1X51kZuzOlXWJ
677rfFyVAVslICR06qj0gkLfQBy0su/Dn+DsusXG9F8iudsnP5szaLZn0pxdGjUGzXwOYvSUcUYe
HgVmztJ/VSEEebFDrwj1oVGTmXxt2DyFH3p2FMMlhSRl28sP6wM2hhhfzjRRYdUhI8yqm2lKyTq1
UkH1cC2eCQTvptuCCo3WEolVqfyBHHdTUUXDxHubyD9mKQMmplsk7ayz/kIXyhdB9Hktve8rr39m
NJ6O08JKlMaCGSlzWFx8uRZ/3une4+JNKfN42D0Bn9E5maHJIFj2fmYinuGAy8/OGC0DqxRevkgn
Cj3GSDhBIS5WSy9v30aD7NXiCBqcHJdGx254oj5yXM7JCvNcTdco3X1mQC6yGOzCgnek3x8rxe9B
Wlym5x8PZ5PkQFxCsOBsYxbFgm3u/SiAR7DAdZ/hYYRPa7Qpc/E0qIyDzxNQUAc2V8YL9Hufv0jV
B7ypOIFKsZ7IwkeafFwiRe4Gz6dYrn/Ezx4PjNVWIzLp9biT7Iai0Ke8Mcfb3rbIgwKMhj5FZE1t
ej59TlslnPVj8o0taLBkKwZz2nkBtQMTDYsRRp5J37zQ8XRS0bS/+RXh/9DxYAvB2u/MSNQ7VX6g
STziUEHRkDgX+RJgVMEox/04W2UA/+v6F/BqST6XMxtZs0iFASN2Om/Y+C3aO7hV0iOt50M/aP9g
U1DDcVrnqRV1S3DWEuNHsY1ZGyUKhpVLAxFVpoFU9Q8w2AmE/6QCi1LgB/LTYonDYlfHDLDe9ydS
npQaLlP9sK04q7wf8uJXKYj8eNSSAT3Gn3CpoJYRCOq3EMQtQnqPqBo5aV6JoBiOTjp8sQ8qrQRN
yJJx2kaSRlBgJEi11gDkTQpTynB8vT6KYBgXckxuZot0QLh5fSTA+rHVQE5uT++2aUBITATcEH54
ywbMyKaQ5AhQ027LzdlKNSdTe8P+wgH/TeUwKz3rBBmKW+WwHRrtnE4VpiYXWtpyjlqJphoN/nJp
B6aAbWwVV3huW9cYmfWecQMO3pZIuH7GP0uXFTeBPULWI/M4gXTGZ8S1c7O21pTWH8Ec0kOcZy/b
mjpjUCD76kuHHRqldfCw1GH2rRSyLZQgR9NFPR0iZMxCjT/YKXZUvRPu0t7ZLLhndBj5jA8WqxRa
xNjDS6/D094lPPg3IpOTUs5dreP+H/gpny8FpzeNghjhcEO6o5wlPu3FKkHHg6c5541fD9yGbIAE
nULzzWTi6GWf9soWDdLcZrRcTiPq1I0XJZxHfqOOZbet+7SfFPNsxduOf7USMumqfJL9XVFIz8sJ
a4qgZip2KqDcfG5TezrPpCug/noZVqZeQiYdW7+c8iu8p6nAvGPHT7E+HvSAOQ6n3kwgjFBm8R1R
wsq4dUhCnZNHQ6rbKMA+qUIObShn6KwPUUCRkIXxF5d+twEZHhyhyDLciEbvCCdeQFcwKT5tLd2Y
SYPG57M4UqGXsAuaz3tdsDI87w1Fw84z6QEXVMgTKN5mIPKPm+NkmYFvoKboZfEjbkLNpl9SkRWE
tDBDBSS9c2MGuDGH2DDOts1Pjhtiai7eouQefyZci2Pi+aq4ZOCSOy6l9a9Cai+o34LI2aT6yO6A
tFSMLuUTOGrrDTopzVR1TLnCv0FuEPhrrH9Klw6VvctkIi10mu2Zeh+i3+74WfIR4PJOVAKvjzLB
+hjCjjjJaZjmhhKxxTDpcGv3niK4yCc1LNynyuzOKu0ZQvXleMTlP8Tx0sa6ne3x9Rs7Hq4sLNo3
HYuihB29KwyozKEE+KRr8i4REwr+XE4irVkP2I4VrxulcPUGyt26RnZgtfMDy7yN9cYEyFC0E9uZ
ubo0G4SsdD+k8Pfdn7gmr1nWtppKmtz80ZC72CGztoG+JDycD9kkTfnMg33Oezlijgr1tEMfnTmN
h9p0fuehaIDYAKwMDHKdNsO69neazeNO7T8/7G/KKlWHTdWUrzmoqeIlKQBYnsfBcIEU2DHj+8vX
rw3vXqw1RfAR1swv8g9fjqjl7KJtj3PWd0Lu9nv0DDCSmEOX1qZMgPkapAJx1RYTV3wzD8xx3Fkq
OPhw7s9w7LM8AKk3UKnDEVaSNmCoMaxHQIJdvhk2saJ3IAk5AfKt+wZtEIhrqv1Klk4aIjQgnFNM
kNIKBZdZEaBscOmcUCLPOdRj1/qK3uWU03Lk0VZOx1Dp+H/V6eOeZk1YUM6b3V9hwFyt108IdVcD
ehD6SBCX4Ze6Z5pqgwogefOkWU5KkPPm6fN5BTvRtXl5JKi6RSE469zvtH8+fxUpZmLQlxjfoAms
M6PNvsAoo5lpLx0T6LyESJnaXBjWoPDmq40+OMSaJUKyIaTL1kg3qiE8W+filyPHlyQ5mNLjZhFU
V4K/5G/BwbqGHJsioA9fUfZq3YeuO4Sk250GeWSqb9ehKZUp4/45bPIDabzQV+75V1n4z+Jwpa8X
0pnnXHwZGibWNzdmebbNHywfm7MVavakYwNxEfoaPBpjITGJf5ykF0DHyi48Orj44pKeHCAByDc0
79eNsNJ8DWk94XdA5f4dbv2lOdlm/orLv2RIQ8y0xbbNycV6klkdEFwfXY6B0mJRNmP5pK2NNUzA
eN10FCAvLhzzAy8m7lBmc4WhuOVytkG2lPld6XzGTuAs5FicCTw7Tjvbc5jKH4cC8ehhi05NRDNs
D9b/0P4Xv1XBBwhzpts8avBh//Eic+0ov1QChFjcEpEwynWR3YL9oKKVbqAsYHqhr6ENHuouUIdj
GdBFY3Bkf7+wLvCTZX4hcNlQzjASYvxtnVUCDgkTMiNntuJRdrkd2bH+OhG9F4f77Ug7QxDJjzzH
PWb5ztDslb6bQN8hVPccSUNmPHQu7NhL1Mgy77QRRpYLCeRAWKKUbI6vxBgwXVSBjGGdGxAy5ynP
vQYEwHoBNIKrO6lZXkTRVIhEpUMA7zgqrA7oPxr+yRGMyKkQ0lQn4MJPXjl1la7JiLMpUNKNAp98
2k8RZbcWPg99GcJsbRNRFeXtOql/2qtg3MHUcF+9FS7nSUgKJCBCYYFuBLdB3wMAp89ierhfG1I/
Jw05aeAWeaki1emKnk4gEhH5NgeSuttUYuGszO5+4oCbP96F4ySVf4h76YdUEib0DlY2tMI1h5hI
/8qmgx8I885Rj5PLxg2nGV7MphGoiEUBzMHFEGqfJ7Yngd9wJSjvvwVabX+2OCrBPTSK0xGRq7Sy
pIdc5i4wc+TicHo6vUzDkaQ2DCBNwRRj8zUc1ZzPHZR6SDm7RXtUsk1uPdN3n7AeMpps76EkT1gj
tbkdjy1+RFcQ/idm+WP3MM8jSWIJ4WJVxzV79Uuji1nOrxlTzcOfWFkxmm9wxAm2cyCRQbsJM9Tr
+2ovk/brK9uviCWZ/TQyY/0h9WiMpqQyrVycfphw/qnxqDYUfv3jErven5COpvWGhZoeJoX2BkxO
HCxSYTQbffUEKvexg8U30vvSM4hpr/Ts5FsIEbsGlsD2yDnYKZAtaGF5j3Ayo3WOWT03IKtBmsZ3
EXSQUiPC1q+P87gkbXj7vzNQyDwO+oGxvlmweOtERlMpTZ1nNQXCc4g9OfoJ3mEKrpS4s6iJ+45l
DC5vS7D1IjoxQohhjj85LpkswU3Wt6R1zJP/qPwpPVEffnM1zldkFava5hlV4J52vxEJVZg6E0EP
QfzqWGlI9keSdw57i92eqKDF+5n5jI/jcptVh8V+gE4w3n04jxM4+BzCQ3c9X+4MaYSq5Wzo4hOq
DxBX+jJ8l0aswYQWd7RCRgmKhlehnazLTVBRGFRaL0iN5GKEfsVkuGuXv6FjuuK6fO9i5c2BgYyO
u/K19BtEHimcBUu7zAU8WO9BcAS61USYe6QvfaKnUX+PSskolBE2BLz7oBCXOZWabrWSuNq8IYa1
R0EEzBAYW/7tWHMtnUM/HSnKAiq7xclUO+vc8gxtGOA0AozClFn7T+n6wpjYicOCOFh3q49ror0D
LRcIOlON3UwXLjKOjtf/06QitT59PK+u2fHboQBDImMWOzf/f1bpwXbUh2Q6UEkn5WtVALY1zb1t
o/6f9cvoPufl1jDwJUQ3QFJzgZynYFZuCxqnrbpwmrxQqVqYV3vfIxFy7FGVPbu4eXAo2wKeQeTW
5KRqO79KoYEdk3O9TB0K5MA3RzgkEe7dHaoqM5nirJau7e8pswZRbLCcnTazbRxuWHRXIc+x29D4
KmbwGS2Zw8OswwxU0RdJhWRuXCHk3ElcbQLbpk1cQfsp1wvE9z70tfiIJUM2c3YH+SoEE2+lxFIL
GR01Tg+7NfTRCdrVuhBPL3PxuILcKTVXoLOSSWUWt3DbOALkBtVjEHobDHqMYcg6iTHd6xe68MeL
zA6OgCkdFJV2cxMQbzQ6FyI427MoB9XtcPE8f+hZZPEgrtVzNxTUpcT6737sj6bF6EgORu72x69A
ZD82llDYwiaG3AMNL7KZW0OzSP9SkRBhaLXN2YJxCy/QA+6gOMbkxZS6HDQs0s/ysmPYpz2mC2Vo
KqqMw04Exg6If0alau8KmLBqpf03oqU5Nh/YF8i7sgZZw3v/ku8XSBcvXkkLqyS1oCBmRh1kIDWv
9Dqxla2vlQVYljN/UcD2vhm3GRiJ0hPCvT/3Ct1TEAu1iAe6WFAOzxW6O/QVDZTKjWXAzpHjVEYV
AJ3hW9NvFlzulS0XVKDcEyPG4/t1N+9i3+ABokK+u4QUYqX6FRQpF9TkC5KSUW41TFNvs/Vcs5sy
YnmtRUBQcvkbX3miZtHH8iN9R5WA7NMsV2IPxHzptbMa0Zn4I1m7DHp3HPs147Kttpwb6DpmDD3V
FeEUPu9HqIKlRzhXAyo0WIGLOBqP7/k5bBn1ZUJ44hgACyzY2ERpFvtxbY39EspsN7Wzds+WTYuy
kuGAD3xohSFikZBuHucQSnsM7hbQQYQqPOwYZ5tKsBVdm1/zSHelWySfyU8yKMfeBEClzo8LncF+
FCjrsQcgC1n+RcXbJJLSo+/9/s9wZH5XgF9q/weFEYmDb4uemZ3T4yafemCuY8qCnzWYudiyUPQ3
4Xag6rT0Su4YKqYgcQq7/1nYM0ufNAjYjKDw3vFyGeyegBY9UknmbxB/pX+2a0Kz8wafG8QFPg6L
+T4CfoCvi97/OsmGxLiQuOi+xsgyD4BowwfebvQ+gEtSSIG75FtGYh0lXT1Xpysq8q/bOsTYWN6r
GBaYp9yef8zF2XfWBGOT6JX4QWq/mpnFFdH3i95Y1DNOFZTY5NAlcJOzNhvnzrG2iEZVMtl/ElPW
Ngz7FZXe4JG0Ls6Yi7llFsmNB4qAXWj3Fe8cmJqXh0u/f/Si70vuU2y2ax7Hzl+Q3Gt0QDRBDsPB
KIpCpaEtrGc6KBrVHHIB15Z8FkKFc/G4ARhndA9nGrhmfo/sB9UrGHHvGDTBhVbRF5QLbG8qEzZ9
2Or/czI4ZdxGZA0BKMJVoBGcqPuqSgxlYOgMIVM/tzb6EFV4YEgq6CHgXggVOuaDLuc3Zs8LD7jF
7pMDoWkhqFTvnZLO6YWRBuXqgKQcofjmfRZliJYHDwa25erLjdhO65seVZpMLzyfMbAYUjUbfEdh
0tpq7HatSCREb9jnJNazZf9+r+vwi1BaaWIuh53Y5DJCa17DKXsXT2nY3PcpdqZ9uadW0emGDvOQ
gdMBQBg2OC8rr+WXBbeHdgwH/BnpMd5wgnQ+7Hk8V+lJzo+zHtV7cUtqc7ivLpaO2Lv+J1ZMOvXi
lt82BHShnXlLD0/ObpV4sIp9YV2Yu0YpL7uq4nt/GevhrtGVNgXW62f+U/6ic1mALUluWPjMrsjx
hFs5QBO3rLqNBi23cna7SnNIo+FTPwQra2AThK88D0ncn/s0Ccywc+W6PamaWpEAlAWFcL8qYjgB
swjxycGATVC0xe3k105mDOF0vrhX8EKUdlF+j/2i3Kwi24eUxzqoHr7EhbuCMHt0wiemw+mZEd8c
ofe9xHFKxFrDixs2ctg2uJP3mIbdshdT60534lnJx/aaZxXQDr7LHOE8M+DGrPDsXCLDQ6zjL8mP
jtUti2M0qWVC+vOpwOSe0yX6Knv5vkLOLJzKNoojKbT441cUQDa0FPN1ZkqnxUI6AJa+Cqj49c4/
IwkgY16b/RCrQt73WhANNEsv6pxGRv4MgpVYiOCE91f7CUoKo6yb7cA6e8m+08KTmxZQIQHE0Jr6
w1/AuJ+KuZr9B2LHJE4eL3Nrvs4pBbiz83cx39/wqciXMLnn0rBvKzC8fi5EgKAEwgznig9pY50T
ZLwgPOjzD5coIiRpNEMBl7hvjgF9tSL8Ra4cYV4w2Ieh9hAMrMSWvzgGEX7C+LsFBSeKSOw3wgAm
odppK2k2yubcpeUDnbNsLMFmJsfYKnL74UsNkNJiW0w0LeqemSQzYHoaCdyiotYuwy7ZYkvPako9
sx8tvn+gAoCUi778CGJ7rXaj98Y2vruNG3br+ZUHNW6NNFUNPfjEhPP7jyCbVUwg6c+Qwb3PuYat
QAtYDGMsYyNX03cbLZj5uZlEm4syRLgU/0/+5H2CCa5vQy+yKchYc9ES4qt7g9HYBcXiqZvMfTvy
CeSq8wOs/SvIw9jo5LqgtCGkEdkPVpt1qICHzSWeBoOON2PaiXvIxvIw6yu5S+Tykbu2ykNZz3Xn
P2/Cdl9R8JurGSFrrsX2mw7muOVvWUyvlXZo9rwax0BPMW2+07xl9CUTBQ15+TCX99SlV3pnpivx
8jSPDXTYfHKzmef4NMEzAL2K29fxLqpidqlQvMhuzIxQeHrC9q6MrW220kmCkpbUfpjeYCX8nn2A
VKrEHjeIGBKf2FsjOFu6AtZUQvhTd0e8qezgqMs4jRfuOlAv8EyNZeJc4t58XZj6++UkHy+jyFkm
oRCofmguO+Uawn9tmFleGuThe1Y/GlEthNY9Z9rzH0j35IOICt4b2AuJNbsDFPGtnrZ+rh5npjGH
OB1rEV0Ve4YaXRHWcy6GW1M+/BV9/i6ff1hATua4NuO2vH8AKcLEfLPgmSbPnn+Ko07sNc/juwrK
k+CxCjkHt1lEqj7xA2Tb8/CFvYkqjLVZfQIwWLl++d2velzYPRbRxpYPeDst8Lzbo1Rmy3aX8JJX
O/GsaHh/V/bfUE5YsAGhm9JY3mjM0ZVHFyzLaEDGyRucv2RHTp/OwvXYIKvXFl/oMh1UhW1KVDpG
uYqKCsOqLhXpgknrjD1gif1FAp+zqpxuguMROFpZrZWYMKAOSBjG208nZziy5hwHEWqXeQECJbkS
RFyM7T5sgH43mBEyYzs2R7R2A2oTp7makrpGjepPPTdqP6HWKLewTkMZCCqAqXDfFYDYgDLaqkgx
MxeTp4BQTf3dQ8kRwKATsCpDCYLUczRgtGUfL3wn+nyCF08afO4KsPi4vq2fn8jZ2Aw6t/luqkKm
GRwzWsgqWdB+45nuBZPxc3luqP2WzTnOBJd/WtBKc2u/I1UQLgzS4KUuNNhDvaJKQWc1p/ak0Fda
gNeQ3Oz7IOp7ew5F+VzYFwVt2UavAIwZ8jIpHT9uJ9YBAKNJ6X5sOX5dvpiiCmq73HkcCN/xnAMS
MTxf2yTCd0/LR3CcE3sgEpGbJ46NfFBgNhbTOKYnEfxu9bkyP0IezXMFAaMTzrvkPblAZDkQJpQG
g26vw26AJ8kJwdPvja4J7Grj9MBeeUlDlbrcZ9o/CA/timPEU+Ogic6rqYRg1it3fkK1GSD0ednc
/ArncPjHVSvzCVcJHhQ2/ntzBD+pDOZFvg7JuqrymOSs+80XA2SDizomum3xF2m5ZTUKfrsfe72E
cTHZz5dOKR0BILs7X+34jiLSu/jFbvqnaLjGzHVr6QYMkNMwawoIcaVQSilKmFtlnAOpCLEio8lY
RQTdkjyX/h4jzy9ZBSxhcmF6dhumz087uFba68L9LqQfowLWv00FW5zY6FkK3U28x5ZdWuOkqxdt
ZrBH3WDJwzujrBorjZvSkaHYd5q9gf0NtVCl0u/yamHiCx7xw4jAnJYgiFfYP7wSbCOyYYfgVfUV
14EJCgyOBPe8hEMGPk72pKjVOlBtYISVuBeANMkDX1pzqdkUXqkS0LD2Rvl4HyP2+/bnKsOg8xr+
GGPoAUK0jt5JHgAijxfeHTiRcIVlu6kViOLk5fmsFs2xcbX9ZyBEG/wHZoY6qkxhCrZgOoVE5giM
70r0ePMzqV99CQ2BvzBD8gHyzHjVMdZgCug/2d2zYlSZyJLnGPwCOKFJ4dKSE2Y1AVExr1mFkhJt
e7Qn4cuabOWSAwh1ikq3b9Le6nq9bAq0l2+1v7PjXnAXfsykdCNfXthCvCInwUpjJLcnCwfq9RAw
Z4OsxynuVt31mDEExYS0MZonMiIMk0NGE/Fhy9R1iMPHd/+HVVlh7H2n2liYInlcErV1jQ+uIzBe
FPNBDZSPu0fbT8PpHGgYERvjyPabJhXLYO0kYRUQWp5vgr4JKtnt1dwvzXcVVVPdt83MrKWflFCV
Tr3gwp9Vd8qfBDi8QEoUiZPElrnGhOEUhhq8foEu/+pIz4x0kEoMLyIrdBDoIIAXmm6nBAcJSseh
d0cKewoz0beexCWeBxoB7so1j5OIzWU7hSgr7eNWzvsq0rgcIscFiA+FLCni7M8jtaT/y5cbE8ht
Nxzgl7mYP9Qb64Lnl/L+Y+4KWuPengbgxMYwx7jiUTZ5gTOacD52qsqcIETvbOSXFgoP+82eVNe1
r+/u6wCnb6wBClL5WGiwrLbuX4bORlgDNjdZWy6X07J0ih3j4I7c1LwqZm/0otHVZdAZsZMdcF4O
BoS7MkcN2KlxdWt/jMRseRQ51rxsyZxqmJoSsCt31VakJ1QdlffclXt5CapRVBkn8r8fpuHAf+X/
C8F+nxQcBGV/JRNvoIWcfdqlsLLNmfEgiXUYk3M/JFVs447FwqfDYaKDpulID1+2L/369FP+ymAV
hdSsi8N1L4wgbySgdV5lgzr7jXuV2Jex0pDgOtrqwpk/0KFURTvju6qRlpsMOYAuEeQExJPstI+b
a2W12YzkPC/ExpWBj7lmTesuMvIFfh7GwTFoZXIDyCgG+ZdReph3f/Iry0+zI83yV9vknbS4iemg
7a6zQ+MNtzqF5dEdlNeh1j0xl6qxoLk+UIJSnC0wvJnZzcG9jMHJDc+Gz8rtHpDuwQ8HhqHIJJOp
KHqZkAks0W5DtQ9iKsSaQ/WAeg4FdJSYpwY4OoOurOuKTEocPOnSk6VYwW6NfqEtBAaM9aNJZ72y
p9hBvwEGCR74Nc427mXwtZTT4aoTxlv8GU+dj2G76VLUdYYGKp7D+Z4a28su51a0d39FRLpnif5A
0kIYdv6nEJzH9OUHsANzt8xnElchEAsUs5sxoh0tHc5v3NKK4pNnoCCixeeQM9pM4vc7rAeeSiiI
V/R8TZWzOzofuux3RvRtoUfNjZxD8n8UN2qJLib41+vKCnXqqMtb6a4J+2JsCDqfafoFTN/WVHnH
V2MjWROpfJJL79g1U67YfSU58nZEn0gfDE9ZgdRuQrYhTBiGWxjc9/bCf/eUnnso8qImr6H63Hc1
JOOdz5MS6E6wo6yMHIhNX5R9lcYhDAdaJUAvebqlF0KfcAvhUix2vaLgtq63hTDjVBEbdPiaFr4i
4QcxgdeRYicoOL47VEfvoT9Z4ci31ZZ1kwP2VcUwoekmA6j6F3j9bjseokaU7L4A8m43nGuD1XcD
1pTjFW+9s+JaCKdHXL0QA2L8ZOEUMlGU3hmlv12N+uO/Lwze3jNcHt9BmRu5yNz9ZNJ3zVpb+Q6R
0FLYQssGmcoKb8Fbg9FzM/v1ZJR0n85N4wLzVOoaVvWGXi6MYqkBQCqAhIVEyadD+GHEIAGLUu/K
x+RsMhhElyM65Sla5I1zpCEVOtMKO8Dcs3me8Sn94gPnhmYKZE6RWlSiLjdUoTyKLDwdgKgkQ6kb
g/FsL//TwLZzjsNm7G5tf442UX8O7XhbWNrQQyPyXRU9EbOcLqk1sLtrwx+LTJKXlCkLzDYo18tZ
ZQNo9oL3FnQu3giX9ziAVp0g6fnEzUW/YnRIKJHcLXTFxwC7H/WI7DunS51sAHNt62pEbabERUzR
Lukw3D9ktMyXVVOsJbMtVC7en/fNzHZpoUcdOp7PjcR9VNwA28eG4xMOeeebE3RNgt50p0Y//+L5
IgKGVxHcHycxEzG6rlpz7k42TuwLwqQqKwhdZb+Mdh9lJZ0kfEwJWmsXCciPowhkV7ifWtuk7Qeg
l/9Ychx3/gqF07wK8pPFBnIQkxzp5wd/OgqTEoRlghBiPUa8kmr/YBusrIkS4BnILMVKf4pHc2ip
4Uz3GafDNYF2s+svBh/+XUao4a1hhFdGVk9tASkuPaHhXBoyi8yVR7rEZy4HsxJv9IAbx0n1QDFZ
q+2GUF9ydLVPf3TnU54PLTrFIii5XEU/d7Ljp1/WloR06xECsdYWfRVK0o4HKmHw+D37fP3CZbCw
SObcGFU6awjBPnqaxUyLMgS45WKk7FBdABmT8GofOQWp5ork6teFSC5U7y6Gj4XuVz7a2lItK6EJ
rWfHmquxN/2cyNP+RyWKLzLRyEypFqj/xzqSyJ4THouSepRdy6aM5nVLXTgQX1eOdwwX0ivsX0Se
SvGr0hi268jZgkq30oJ8Z95DvL7EDc+ckNx1JSSeUxwqdbMweL5Wh/mdLaUJZQ7Yi/I5J8FdNwDR
mLcGlBLRFtE6O67CNg2/2bzjRG+S2nximfOjilI/Wrgx8UxoTj55WWGdBewHgmpLTpfljYQV3b8T
IHHEkodOkAjgVnmX2uUL4uSi64k9opsmeWIplc9U+upSzYh+polZyUA/NEQXXKQC8NEyepp3SiVP
vjk5mIEPU0Wl8SIeE9O02WI6fpEjKiBjehSriqcxw9FhslgFoQhpZB00BCwEq/wDt8gP4oZ2YKxz
LyPJSNXss6VYQuM4NJN4hUXItuhvvsPB/bQwIkvWxu30uWpq+9fXjhRBRoL88emwrbbF4mkvwmch
ZoQw+tKVS+ALvXoxi1zNsrZzSiyL5DtIbpTYYVSaVyHGoGYOyXr6VBkZYLLw1WwthHu9adKNTy+N
cLRVlhZwXY8s64KkIiXg0XMqMJv4OMjTvAHE2FjQZeBsrQEzxmWH+NrjwZyYTXp1mLP/0Xz0NaZd
fOk4JJDG3ymxWTifxoaLgI79ERT+8df9Hq/brytgwR/U6B5eBE1CO6yco9ebAQXigXBqqeI7CbOs
3LcmZgWQ5neQ+y9x+qjeF3MbVXoAqdcM0FkelgpByuLWcmZNU12NsX4rVLXX4IboyJcQMryutiRx
o6TUCj9AeMpHvOG6woOG6CS2wdDZkkNDJ1s/eO7Fpt0TMDPzJDML+6YgKCiJROXw2+jDjRkZYE/h
SIBF3eU/6GkYDjHm26Wmmx+gpZfCLRbqI+Smcv0wcMAlV2JsFmnVHtOLa4X84/JDtuWVDjlPvEfR
6aKK4JsAkmFYBCjjJLvPYqu31nRLSm9VuZmBMljZoIrWPgzbjKMEsWd32WJDBuYiHv+sg2i5OdGd
BSroxreiR2aHSVJXD8Pp93R5moB2QPnxRRGPum595gDmW4IEMPsM40P7HaDFMO4Hrklyl5y8KCwN
c7kpDs+8PZRxhDZ1M0UvL9iV5Z9iMbXnHjvtsIWrExaba329DI0SHNOnYU2ri6Y5Te8fRQKn44MC
aFi1f+Ka2HcP/61UtlBk2y1Ih/u1Qs4ooMpOUCh3mcNEMZhDKyloe5cEJ2Ym8VxwLA0vfral87A6
s3bJqyS0x/ve8qjONBU+g7dTHvzcUGDbGlvUTUilzjJYy0Hnh7iF9j1rGTvBmx1TsEQymWe31s3+
8xqlKuFAFBeDjM6TRuVeaclBzH//8B6Q9Vr9yf9NLB3Fp6JgRpuIe1EZ5mdV6QzPH2TmnyWuUG7I
p3a6go+XNQGzxPS56SaBTqYwfMMX6xoDAOglqOQ3ExXT1rZXrASPthqyIIVpx9+aINTzBUHl4D2k
82pROh1jAgQWhYlVDCkX87yMupdi465BFYbMLZDvrD6M7GQH0rZsVdRsQ+MUDi7Du3EJaOMfvvbQ
VSMF2dLyjylsQyOVdpE1Qwi/HF/6KBT/kLX8RBnVKlpWyEwyCE2LtmU/bgSXN02HRRTlf4j93dpr
RCRfiVhakMZS9Hzham1QXdxKiMvNSAHzRERfLnV6zClS2jBFIwkyeTZS+Fq1kBqDQMK6I974ocu2
gBCWv2C39u7Zv0tC16tCJL0mXIeamI4rxQHJ9rT0vNWISnTgaG+dbV3N1PeTa9GKLNw3qI9jaBkx
tZKMFLmJ7QmiOeORhO3EWisyczunz/hJctO0kiLr66ymqbJBNw1sxBOduHzR7aCOsY2y/Qr1+Gzv
1pNKXj5Z6+982O5BtpZ98oUdThTVboZ9LrdXH56TuY/s0gxfbhEiSpb1FCy0VyA/KSCs9gVux6QX
uEqXwmbzSslmQcXICDySGBtVPP04kjKUaFcepdM3x51VS65a/J8NIfuSv9NpyLv5g5WgUevnLlXo
nr1Ol5Pi1RG2s2K7SX2PjEXg8jHNRlU5jWklmHfTjOq6jAfKy+eGIGpJ/90HZh9u63eqAU110fC7
LJOvr/dt8EwzO/dBsvoO36p68tH4SruqDcM053gJ4RZgfTTUzTlpTeltv6itUZzUZTnRSZ+9j9M+
5oJ4YIyZw/emtlu+2lWA2eWu03GZYOn1zn4CRBTCBhU+iyw4SM3Fk7WzIiA5UMy4qZakMJxSqi2N
kz1GUptmOIQcc635YAv+UWahgBssMevkjKrETNJVaX/HemGz+2bOGX6z21Q4T2DQtNZE+HuDoKdO
chZkxChrQOha0yJx1L6mXH7hAstXMa5kH8qU9d0Cu4pKsuerJttKLXR9sQWihTYbDd5tNs3AUVqb
QQIYfi7fv27655cOWS6n02hjK08HiM5iIvIoJvIBWKexx5o+QUKvJP69SuGCW0UVv4lPFthL5ije
TV54d7mxP7hMhuN3LIS1UQtV91tpJVd1DCQXG/g3CW0zYIlAAvMr9M+Lw1uAG/5fZrlvqzzRU4A3
Ta8kS2byZTANMY6xNVXTRcRsG/HgvvpYBjz5O9URDnKLOxN/jTTDwnVitI6rYL34f5hKaycY5S2A
uOGNlCpVrqSxvZBX+bnKW28zCBH96vJI/fVGshXSYHIV/lr3e6ECiSXA0iZ8n263GWyThqAP8FjC
Ly3euxXzo+79d6CIfwhAwdHrEr20wkLTwNJsp+8UtRXw0TjOx6syQp9UrnK2TD1GDXKENXqAEn13
HoWn/WiKs0QIzQ/6WlmMcRURiSIvzXjCDIFiO/2fQmQDHykezvBpTd6KU/GGOmNdHng4abbJbN9F
WDe5CrjUxoxb0GRS2Es3SLJqKkDvAxn9ccaLb13bt5/2UdiQ0wm6OmuiZCwIv63U+FXmBaFPnahz
GF8z1nzH6U+S7awOo5YVo5bwWEruNUvMu2kPlXUUru/qmo8RYySyN2Nsdb2XcQjXid6px5Q1LxTk
1UUzpAU9jkGmIo3UsXqXAUHXZr7mkb8NHavQPbDwVcHHKWR43RxNKRdTlccGSlw1Et4vMzYflLHX
Pnm+eFPmh79kdwH+q4tLb/EJTMEVxKArvgXlqMl9jRQAxsJVf/8GZa+zlUjYF6vVyZ0j4YpgM22X
EDjiDt76nAXPXPmEZwaCe3u8f/zY5GjcA9OXavVHxIkdBXKrI3YYq5WB/TCu6DCuD9TD0QDEBSJE
NxceXGTwXRtBl+juRAmGPjUMT0vFm99Y4rjzzSXf3Wek2yVo4q7xzAhkmLsyUZk+yduZ3Pvo3YN9
sMoJl6KoH9QgcGRC3HucFf7g3j1YY+p7Ld9TtU7HvSSP8PvwRKiu567BapZVokNpCr/Y4KisqsFT
C4h6uL3Q/bsDsv8tCn5BkJvXtPJ2KLY72OD6DjmaDvya+yYDPdQW8CgAPcu3tcjsJN17I65VBmMA
JikjDDTc0UI2X5JBcX9Gwu8P1wbVhxr8+9XyOw7cqDwyBCG1qeGMs1aQAJTvIO0snErNfEPkUVjL
FupSVu4FcEK1hKZviVqJdj0D/v8LEqqs4F2IaRAvBdWluWoBiXjjXLvR4swe+56T3Ipk2AalH9TB
ViG+ut4aNbT4ZMdTOxxxt+JA/zod7TXi4Vi1U3uRKPHvFNH+kCRNyFJL3UAMQA9XNYdWpi2INHaz
SRdSsCxPnMHck38dzrwt9GaGFELr+sSqCYruGNRK557Ey31H6vZV0cqpqLtOq/3Ydy6hka41lYQS
2YT3g6ZI5WOhDJr1WnJFF/3JUHL6SOX6PPwaJ0u/kn0NfXDPNQjUnnAxfvUXaY6D3hS7cm2Mdx6e
OMa9mB0Tm7063uiEx2YUXq3vyHBvU65VKC9rGf3Gm6XVB8vphytxI1v+vs0N8v7xtF5vmHaTEFfN
jrOldqwmW3EwosLtWS1Nl54Qn9bMpmQIcw3iHEAETfzaiCcnhp5h+oa7IRN8SuTkM/lg9XFqEBfN
+oQ6FdTDCik43hJS8RsOV4VIb1dipDYkUdZJ/dReqNXhRsLI4VGEi1uitgeS4tfyOxD6v/34G6Q5
VQt8cuCaV9WMxfHgr8ckS1u77AJWfi5o3Sv7yInE2NP1F90lTT8P+9P3edwTRddOgFwW2qAe5SZk
Mgt3qST7X0c2xtftNaP8NGndrT+KC+F4rlYauDuDEQKTEWhHeGfvc7c7APw1PoOWLRrrsDVwJq/O
20O7Mek0LaUypQjlA7kC4V7/tM6XchRZJ+OhoEGEEtEqFHLIdA1FvAln4QkAT8Q2zyvTHvwSgQtu
GqsF4Dl2BuOY7g/bLti/Cig7G+KBdQJS0hg6XHcX7yWBRy/8u875Y1wXE7Rvfo0j8zQbONV16BJC
Ebh/4sWGnt8r37ofS1bxDZYYWIC+UVUDPkz3j3qCymZtKlWJM6ZrxNAK1y0Pr6yk+YD8SZ7PMgIc
+ifsvWee9EF1t1JvbaSHz6DDEO+/yN3ehmnpG8FOqxwpRy9KB+6f7oDz0fRniG6/QKY5vOSQjvoM
B21jADmwrK7g0jCGMIhOuty8xdco8qXJln58a1lb0I/f8Hj2GyuvwCFweLwjupfBYqtAwqyMvar6
ZiWNXlzhQmuJJ3ZPmzxCVtQ8G7gGlKfHok41B+wgUlF00snFe9KOMDqcWXvO//TFGtku/UKxLVGg
G9KdENAMVQ7cHaKwSiJ05BGqtxjvJ4jvH1UhC6nY89nqWDR9WzojTUIgerQNJhV6gOOFCb05vfDF
g3n1mFozN7s8dcIXW9e78Wn3LBnTRmumdst9D6jivc3JKscvIb7jHb4ro/q9yRQfnktkGBrdrvdy
rHmVIgxipJz9GMSBxEymtye5Vf668YAkkRkrr5N9k3mJDytrQvY2w+hONz6jCNPEXkAsSGRcXtbR
b6/ZpDsPFA1dWCcnHDIIz9TD21474a5anJqgTDsvNvA92KK8mEGssx9FeIymeDB0JhgBV1k2A5WO
WxP+4vNqx3L8eO4cMpj3BP5beZ+7Pr+ZBOPifvN8mJf8EWrGmRsp781PxDH2OWn6b68/I2HlMT0N
SURWWrrXaYFBD5gP0mdsqnQJ8Yzfksn8kbYrlmnJynstMz27oZZOaTz1sW21dypFF966MT2TgAYZ
ya4IhOkFqeZXipf4OHW5YVzo0aY9NbMpKPsFGwMMgGusVGVT0rYycM9S9EZsDMo1HGXPQuNT3t6X
58UW8axItXKVhfI8hlIQx4G5Fb87YRKoQahifxRmg1YCKOqa5Tt5WY4j8Vxv2CIaakWE/yegJd48
ti4C99uBBpiJwBdiiorfsExMUzroeeAMFvDCGEkgklMRuI8wLtDuYTOgt/zqJVnV8sNfsiAhbpAX
ezHamHNWSb/ZskGhqx/dAyEB7ktNloOlrYDCs/pBe3adfn6P2uOyrd+0Lz6LAxb982yEhsoEVwHP
vI7xhIIhHVvbi7kR0RpBnGL5PVREu9J3gROGgSsM9gyqOdQVTU5Tg7Uh3ZyFrZ1PJv3n5esFBZeD
MVDsx/ka2MLhwIKeHppGkyWDNiPQfN69r2eJNk6+jf8Bddv2rCxHzYIfNVHIc7e6/XHOWpuzlRW5
3TORTp9aQvH70KERcyTNMh53TQMyr2xHYSxW6+sOh7K2wwyOe4r8Iy3ahypki0WTnVHwhkO8tu3O
ZUsVB+WNUksGLY0yCMbcCGxZpdpbRlFmLRVvi6NqlWfxK3TOmJbDSrGn2k253Y81CwHZPseblPMN
UVHJgugYlDYgzUNTa+9dZJTE44AQPqmjntAzLrBc4iaQVNgjcDBETqE2PwoZiowp0q3J9NhVXpRs
Sp6/X8M4hRydVL7Pm5LfpX8BG7G4lVeiM8qQuzY9BsVguT1HAq8YiG7T+K1p5zFzBL2lmiuRyBgd
3mDfM8M7nvoVloLpW0xoSeGySglR7OU4wqq5xBDceRcqUJnT3bGgAlN7atPYrRfi5sCGCAGZG5Jv
SyaiFsLOEMR5orJFKiyJcEP0ZsfRtwyUbs/RrbLop3Pw1+RMB/KDGlF72Ln7RXJIEAYbTNcq9UZQ
TaoQP8CFEAQE+W6iUTVDz8s11Dh7UpPQRb20ybeu+0S/cNRuqP5r+9zGF2jih/21OLUI2M4NLKXG
MxaBsgBrgsXhfP88OPrsbBlWEGM4scrLrqVkspjcN9fl7yFkjnTgLWVAhQFpjhdAWgwZXhHHS9mn
miW9cUTJRJkWaVoTwoze2hJPk9M3g9BF5LqDxyebM7C4TQcJo1nhqzjgw76Nz+zrgyefren5Z2sb
pLb9qvb5sxS74jvgbt4f3Ojoe9IKQdyrU7eHtWtOo/h+2iYtZvWzh1FpSQ1J56J+3RymRTVY1zgB
g/tR88WipnFm+u2izYq2H/KzT0nAXw50bUihlXRM8kjPsSJ+wD+85bzzVdN9wwN2us67pGX58U2w
RwLZJxz4/EL1zoTUmJKFqZJhFF0CkvmMl57ALh3ddt8AAMM0+OmM8k5veIJfC7yvTS7tGHisf8dv
tKJjJy2fwKepfUkDgFEpOOcYDY2oqpAUOa3/LVFNYYXpFsZXB8ZaeC3dZeBwd7JkWPqleu7vos3l
b2JtyR8LReXv+3JUWwh6SeiNJ5TXPBxuO/pV7WtjmHnbHVkcy3t1VpyY+UcBIhy1pyLXkFu+A1Mz
7k8SMc1eOIsjkSq078tHmirqoyWEO/6y9xRV4lfHzLu06oTiES3/w7AsO9SqVzCEL2AurG7T3LJl
1gLULodB26EYRSgflDDGhbIZakeJeSBSY433qN+fvzQ7GWu9KTxuL3lXeaNw2jzVkriquaW8NODb
LpZgpumEeJKGhL4Mdxmww3osVdUCXm3R27EMPXh+xp2rGX5TB3qfN9dYIQRGfchAn39HdOxCBytt
2mwdHQChbjwOR3QjwJ+yNYc1kC3vzwv1i+NCwBigouaVzvZLn5fprEN1ztEzKwu37qu61vR/sL5e
EGMwQeUmZ0T4Loe34PvddH+srs6kW1Xcta25J9lBAovdfBVRB244AwUPQFpdJjExnG0F62Q/oUMN
RV8iXnW8/qbqCcRv4wWVbdMQapcM2OK48Mm/Kv/oVAAPXVzZ+FvgSm13vVEHP6ITpD7OGFf+zSmY
3h32QF6uL7kRcuGdzFLZ/73OHXbRoMQslkdO4OKUYOP8Dm0Iw9sJoAPznmmAn8cjfCwX/OAIogCn
YB/y6eBkJr9T0UNY3K/vUop8DsCn6Gf1r1W83UuXnFNPuO/dP3h6p6oiYc6r1AFPWP5JJPIDM8oy
J3eizUZyHyabmxmRM96rKNZFYuB4ie5vXEzs2/eVO7qsFHPVCKGV940/Pzibwqeag1eJ9Tgdz5uF
L4sv2pQgAoEx3HxETLCBinpmYppfkNd8DyH2WvsV+O2PLX5B7sPidLkuiFv8TCcCCk8t5FSVFdVQ
UzFGk3Vup2KK8aobkAE50m+pAgecShgpH7fkEP6kXuwwoExzr6FtY3TVH/1Fy9G7wAIoumZaNOxi
5GTrhIefuijGiwN0cZ+BhUfvaspeaGfP4bzfFR705JUhPViOpbQcQ4Q4AcfWFDlIH5StrxRTzpUQ
GZcS4Xir7biFHC8PwVqSmCP78jseyq5e428TCohfSJusyRx1K0Q/iBT9SkXl5W9bwIoT4x6jgDOW
NJeRBygy9mtFz50D/MA2hAtow1FH6VtTh/zX3Q4wd15n+CrskUHEppNCn64XLf8U9fxeRZSEGBXJ
Rj0lXHy4HyrWAGfJ9wDozh1KwtTn9PIOmpelxsRCr547UtvD7vp5IylHimUV4PfEV8szkuA+7CZf
tfsMoPT3rmO4kSAkAVs1JT8TDUGr3Dy7GFf2xiQ5YVApIFEGNNDP2MjhZWqIQ8eJxGKWEJtDN9PT
KW2CDWmeYBQUZC1mmPqiQNPayna0BKjnbJIip9k+e8c6tiUVrikpW5Ju6+qxKxDiDRhrcu1m5SjQ
A2xboAowgdqZ1uO1J4zXtMq7DuPJAebEHFIG2m4Srjd6tVWzA1hmtEY6PPTPiAoGzVeGg5ZF9DG8
Y85zsM2HN9zLdU86Ao6Fo3SJpQrOAjvVEcY1grTl+CeWH+x2i80UZ5D0jyJppi9j0vxS02z6IDJf
cWqkKugzxO+BZpVO7OE5wzTWZ1AKtL71UhSdWT4M2EeD5LILPYnsO+VuTj/cul/dS0KDu9/RwWgG
p4DxspH5rkPlllfnemu4xb79gXodnXvheAse7UCG84EAKMVZmjd9XbPyhx3JEn3F+SsxcXDIU5g1
b9cQ1CdRBJp1A6AyYc/+egGu74oZfCtLLkRF1c1l9WCd19/yHMDhetrJ63uO37f/E4ZEtm5N4+Ku
vzN1UQbqTbU+0xQVl/Uean3lhfKsxlYc3gVAY5AEjzJr50VRmry4bK5+0QuwhxdvGwPgNLxFka8T
/ryjE78NkxWRrPWQii6tFoghaN65P6Rc32hq83hjri4+OX+PFTxR76tQHuOc7NKi/H6yGzZnnTd4
io8iIUG8uAp3PIBUyGV9UTPRQXzJPt7Rg1jxp7d9qM38gtt31wsw+gbEWoQ/wnsBs2kscheoV9IY
TUmij3Fjub9qrKXuxroLky1UNtmD8KdDkLjyi4pfhoaBtN1xganccyq6mmIlLQ5ZtBPqHer+T6eF
oVpVwaf084Ywrek6eVp5bdGW7PxxMtsD/JHpFfAJKCSbIlSaiXfHeJIB6MXKw5i3rq+fazK5KBqj
dgF7h8jo81ULP+Sk8HJY7PMGlB++f+LYbPOF6oOo8P522G3jqU1xuy1tNzcvQtQXiSfCW+enwxbB
cTDog+0DM1Fd1Mo9xP0BPjnEMkJaJJP7Pwk60xhZBrMNC+P9El+8qVYh7tEsLfLr0NlwMylxtn5j
vLitkFesanFJ4r/7nUx0n4gZvbV/+LgAEdg+BnhfPo6E8oht3DuwxZPBNYIunEwpHdGe/tpkKBeo
1VNgcf7l742S6CIUTCHNMknQkzrJ27E+8Kirsv+MD+8QY+tPqXpCdqVT7WigYcmUK4a8UqaU1FZ6
/KTjBjyJrQR84iLThGSPgN203LLHG87paxitmfuP9g0V3+NSt66W+6wqm3Qf5T38nDoJE8TJCREH
7/FGwYVsM89PYmeZyAF1ZCv0uljOu6EFFA8Gfp9/TNSvPQSBmI9vWaYHruE8MHMgn5d7/osNQi/8
zpCULEJX+HcDuRGJo+Sz+In2KsKUbcPO/kdg5dyUZFarVCs7P1eBqFNzhO2HnaKIwFpjBUxgrMT6
5cTWr0Z9CrYaWKLZqlqwAca5P+VBirCbbHqnPmrbTHwIJZgHjY0+MlJMPwNsYk9zPKdhBXdDsck+
LInObdShaYRDN4N0OQBs8j8/5shzeA4QVAJ6VpE0N1JX+6urvf3/Tsln8Fc9y/GrzwnLWCxof6BS
leqU81Zl7jP32N+SIlxUEdg0MVNBugR9OHsgkoktxqWPwFvMyTSk+9iAORR8NU6WSBriV/e2gIVc
AKARNhaX01wZqOc7E68XpBX1qoDkLoka1Npp3KiLQZdDEJ25sqIY1tYDvFb8uKvWNYZy7ChJaEKk
HzRetp54xAl4NPd0bNN1JGIQKGSXLA6P6PBSp1mC4Wy8ABX6h+JrvOWvAAT6bHMkNitx2GsuVgfz
/i3QmrPidN2eKQVxdTUnsHaINbPz6l1anSjEOHFB1ikgFYJ5mp6Lst0zja434S2RSN9ST1tjtThW
RAqemCz4Ed6wmrZC3itxYd+Eb61Y36r1m9jqFZ/Cwnd5+BB2aIf/uukEkJ2sxvGV04IqzZee0cit
ETHhJr4AxCfQmVeoXy+4A7T3R5oQ7jzXLJ/KEMNjQLMoIWwNMklpYvf0apUj9tRLJeS+YzD528J3
0zbqrpHnWPYpRkoG2pGlirPwY1RRyfIyneJdY7/Y6KpMG4IMqjR8U5ppVGjwwKpC/8LOiRfCY+u1
3BJKHq4t9kI9B3TaHO80aDfWuia3WLcoXqPYmLa71cDfgygnIw9lZN+7jKeoQj9whwN5JKhKghXy
fzzrHJuzoH94R0tYQbBj1Mm4PevhygEhBzvhCETWvFSGkahJWth7WY/T9bo2PVZMo1ca7ME0XV+z
3i0mQT6ICIAcsOUOAPdC1vBwQRwJ5cAOoOjH8R77TwB5xwe5kJSaSvH/cEAtD1h+PqiOChZJgRs/
mnhKd173qwvcW/CCHgHzbTIqk+cv68wYhsSdf33eL6TjSg7p49zEV3++HxRCwIWpDySJSlaxGwbU
1shgfbyFb/Mg8sgSlNFh85OWyAccDY3pHXpp1jDUVoSCXeB0iIY3NqdVvKqXp6BfxMeDzeAnv9VP
AGG+tX/EwlZ+DtN0g8RYugh/EM//UCvCw5DPzK59aEsxEgNAXGJgSOF0ZTwKT3hdnqs0iCb3kGUM
cry7dYwYasw7QHe4hBR1UaIlN1Gxs2aAHM3JGAAwn1dKV9yYHw0CcqKJWGFqb3Ray9MoYYtISVl2
VzKOb4tMqj4KZG1VRupaeFfYE4jBdJKaSytYwDICGJPrkZMRyRItwbzDE54zqrHVYd0TFbqJku8o
T73weWDW66tAvE4bAfT0/RMOwJ6GnhHaS2w85h3PDOzMsotsrwVtPyo7cBs5/abrhfBvW/oLbN6u
kksBKxIPDweXA2itt14oA9XLJUXzElKdWsNI+M1bs6rq7rCT5x+z5Vh7oZW5lJM6bNPZ52hy6GU7
ywShyEEXDPaQJijhQtYr97KY5y/vh1g4IvTZ3SoCDeW0af7gqDKWJ3TXj20KbkmOuwnyzfO0M8S1
v6Bkklp6g6M1kkiOVsEkCT2vapkyD47VokPsI7XeIle8kSy1nmEfEWTbj6m6GOZmWaQ0VLzCems5
fmvmmiIuvYQAD41zuBd16kit8Dmfhn6ESXeqb6DvFSHVJ8Nwg2QOdRGjxhbCQDNou1lqqfO6Ayt3
R951/0NfVhKWokaI6fVbFgXdHsJc/n1du8+KfRYa5DdnQ7w3f2t7P1HwEnU/tyxQbQbDO6WXALgG
3jxmD937EC+D+wd9RjXdZQjscuCdigtVo/MpnRxvTVwCx/6F+cIl0StbvaU9Za+XHFVsT9gBnvkv
v/xoFdKN4jdXEBYnpkRD9WAgXAZw2ASDIIU+UHLP51MsUG3jVPpuNQoVhRMV8LXhE/iT9N7zw486
WOFJcmm2AeFqAaUg48yEuUjWb2z7QMdksGdqmV1IzIkAffYovHTbp9NEK7rG+iABJGh3G9wN/Exu
nkBqM4ElASnLfCsL2glwRmP0FkLPStPREUkG1BvZxVU6PGG9ZgNeiMSzvx1HI/o3OYN/U1i/CsHT
PbNiLtwaCmbp/xew5D/ToNtBcbA7L21tCXywDpbDM7zB+6cqHzPbt97svdY4AC9bBBsqh0eDvDyD
FgXRBGGbiTAa3AW1F6DnqbAeHu7wcnmlFeeoOVXnoUn+tAiCdz1uJoBy8PcFeSsYF2VXGjGnjX10
9kIzHLJEk9qNd6OIAD7DQhUrJvaowJlXAb4D1bOsM3KRDytpt3oCRdHq/MuaEwzrsCbPY11/mR29
hY45sFDRqWtuIIgS6qZeHrd5AjoJ0SCWd0+V5HQYTaLaGSTepcO35I08Dkf8ntKQ6u5hpRecoAV9
7l7y2qoifBoda3J7KQDtbH7vk7diY4QClVV+HcqLOAhG+PC2i/b8cu/yKI9tL/d7s6X/83QxNO2w
H/um6sTf7lZuVCGuFZWZRIQnEwvCn09VqGW9wFMOXG60hylQVzA5ImI7TspZTVUYCFfy2sRHqFZk
xs4xHBBZZh/cHptX+rS4JQ0dpDp3z+Zi9OoCpz9vv4qp10bAdHAuc0kqz7lHLgtQUbHW6922beyv
oeXnHCWP2D8paeUK9KZf9Iq0yJWBI6xLablWwX2MT6wSNzhmkWlBDtNFScm6zhPukxxYxRX1dcmF
R3okX88DWFlSKkoL/4V+eY8tWn/jyn7avJv7eIGOFM3+YuC7LpVnz5E7uQvjKuf/RxV9JGuRhl+D
O/ju8J/E9BY1ZZxYo67z4W9YFCvl4SkVThg/VSTg7N1DKgDGjSJchXUaVWbKQtqwXkOL+tUByBDh
S63dvxFy58dwYgS1k6TZN9Fyn7dw6zEvg9RFGaM5YYQUJJ7P6VP7OcadjeMQ1cgsiYluw8C0/Hdk
6d7e9Fio9UHcIr1MppT29xYAN+qGGMxsPrx9VxRXfFU9PqDMT9E0eOKegnEP2uJRmT86O/r6YBWy
hxZvgKjWydjvzhEssUHUSMR7cGMWiJTWcAY2rcd7BVyllTWu0/bwrrB2/dKCMT3XsWUpqAph4lWh
Dj4TVoRPJLobHHvfNPWJTVJgMnx+G0e5gvPNonMMinjhk0xICXxSJUvO2PsFyjZR3HOiBt7fqMeE
uiwhmDbIkDvHxA5ppSkZMoBotmWJalOASzOJN/S5kiG9yb+iTC5Y5ChQsDCAx9RU7zgx+/0PHaax
+uNrGYSymXt8WVP79Qxf9eMAARIe5G82Hp9JU1hI61g5HClnXSDHcXEi+Cv6Sjns6p35adQEDliV
2TJEwmx/PNlOA1tH3OrmDsCIafcLdnxsfyb1IlDwsuEcFHIdTVci4JtUSSdCz69TdCOfJpS5tkGr
H2hhM0pVgwDbKEs+dtnfKPdkgkstkPk4a2I2+3k/KvUmPQrUmCrBU07MlwomjC6aIFXJkkROmHOo
Jl0GE9wI4ODkmGGQVJ+rnUn0vHTZ6x11rH78H2KS0Zf4jDphe3XmxIaYxc9nShv2FT82wxBDhfiy
3bLzOH6OoZ59a2NKp5EdpZG3gnb8QNAKzVLZJfdRMBeg3wo+XFcFJeY/bLByVMdtSiwX/gYfD/cp
s0Mp8pus8QPHV0UKXhftyzG7eIpTtHBD87kocQrnyd5Fln2yqDzfiOF1VuthOfmg9L2d55NQlfo0
pAQieamOTjNnpCshRjLWQmsDQOTpKobIPt1p2IHHHY2LffdO1J7aXjGWVwOGwvtiaSPYA8hExbC2
QPfAJZFTip1B+rGdS81F7mLyDXmG3P/49nmq5hwTuLrm5Rpw1tqDEYx6oqDdUk7+IjwagOjYQ/Ld
6SaRmTAJ9Fm2cSGF/w2RsnSihw5FM0qyJTOAxAuNG9nUOeX98f3mfMKsRr8YgSxma1vgvjTekgnu
0YONWkukvkTf1M9zoeEYkOYNyYPB4HUzO0+NdK55GxwIOtTUp4jP8jCf/afeuuC+D2A/o4lAeFE9
vWDErhKToTLcQ51c8gO9Rx8tKcsfpwkBeifw1Bn2noEu+joM+7ftYKyeCVSLRJCrVi8w2uwfMqHI
YYJ3Zbi4nc4mk/8nkQseqcukc2+9sBygKzBt8Vc6QKRFJStrhKQHBMMYKn6tPG12b4QM50mLZ1Xf
n/c3vy3yf/fzs2O/UP14crIimyzQ4w044PM8R3OVBXWgjxgFZVKcovFWouPhP+h+3/seY98JHdAt
sIwgC/ciZbTFhnMHrHq6bslp+kZ8R68ykzFyQXS9PyziUkp86HY51BaNVE4F6A7j43nT8Y2IHhVZ
+RBH6ytPQsORfn6ceNrJtGfX1+5D+Rr7daYlFeoxX7DyhGrxfhvJJsWKopTjixF2Igw7LvS1JL5V
Q1vAgZZxpRK0cZnRfkYOLsMH5q3Plxh2T9JQB2RFWYAWHXq3SSfMBgNcEKi881SfXZuu4q8rUev4
Lv09nM+zxOCAMaABfct8Jkpm6JCehegkZQgrrbb7i7p2Gh2mvuaEybKN+zLbV+cqvHSd99AzrxUp
GCqvnR7o2TB6QwTP2CofCSlNpWU5whsmkL3JQC4UFcqqViKKMjzByoM+3Uwdgst21xjJRdG0ZBDf
ZARDwFc67ZvMszuY1fcDz3QnMNi77GZ0x0h2XKvV8fQ0w+Tt7DoelZ2lcwmEjcq9hqx2T5Z2V86P
YJ/emGunVZ1/jg38gJuBoJEbf7rUqtX9D/K+ZV4yXWcKFPmV5W0MM6foA6hlAoxEKdi7+kA4514u
ZHnmwtvpP5ORb0z2airL4EjnLxLZHy9YrwCS85qA0hsq5S811Hvk2eiyLBT+0fOomsFPN5nXBXzB
ylheE7dgesJFVBO8WA9Hmp8rdgBZ5SsZPAeRblmBYmDffkHFyPg+IBzjy6BYui1rV2vXokgT4rTd
w4eb7j2eu96Y2i12rJynemSPuvPfv0sarnnXCQqsqrtEqGstH6X29KNXn7d7mtg/cn2ikpS1/K++
cmBwOJWcwt7SAXKkr9otEDQmNaNp2/2ucSjD0NCqsZVDDsjgp5u9J2YVeJKCIukAgYHKD5TofwZt
3+IJAll5WpERG5ywKpEYjWg6b93S0bogAuHGzeLnz4KMWf4FeC7V84F4wyWpmUHMzHyXg4uPn4NC
2wHzl63cl6ChFC0y8PXm6AaU2I8KmMPwsSrQ6UjrpodsEu0HmpSt/1YLHHvYk8A+SBsbm2jhNotc
1MKXE69KMV5yd7hl96xbzyfd6hIOAkZ/CttK1b5PJksiGtepvMoNMlZymsAx5oN2DDrKDADk0ejb
o0ADUcTPBv++QBQeQYBm0o+z+S2sK+BxBxdyi/8eceNpd5YwmVuqEu5ILncp364vs1GWbrg5tZ7K
Oj6qZgkrpK15FtaW4j9blnoch0JZ3hBX6dFIXvI3evRuMM96m7j9Q6nlE1RZtub0Wl9M7Ce5nSu5
pYppeAoxPM9fioWfN+wmm6+gcVM3P4V2tlLorsI0GZewIUhtLBY+EZhremkrxsJ4SkylWP2snfL3
/wZIYXrJCeMe7tJ74cc75OzfdV7o4AOE/sHB7G4RVGCzhHqv+LCPzYOoLLy0qbVM4YVhQsWZ/TC2
fdXE8fll9H6kbjm/PWzRqRVIgzTL3blWdCDaFnczdSIjptr2gUeQWllPggm6/B8Hac9zbTbtcRik
RooWWbCZfXxECttYL6+aiklUNqxpULCVAJAVOTFCH6iZGSMT90U4Uxor0a+2xLUr11AcmR32Nfuo
woNAAILMD05d5wsbLtmx3BJy6S6wd8CkcZh7cWvGT9ybl2YP66eum9Wb4zzQVp9rNHvdQkH0Mejg
1FbC4kRqMTCsWKlOhkpgwcpcLjmev14Y/QaNirm8QZBNJ8VTxyip9b2DpP4S5GISlwuLrQoY8NYi
yIBep0A16a4Bl284Dkl8O3Ywwy5/TyoqCIhO7Uc5IlBthpQ/+19PbnVFRWuvdA98+mbeESLqGkeE
BAIa3pv1IeGgT1FRMDVe3RrtV1zNpUGsjbIHocDEyxTF2HTFgjYi/ZlIXJstEVyZXp43Ipx3r6bU
h8v20TBJ5WLMM0urTRE6BM621H3eJb4ISqLHIPlKi2x+Cgv0J5v6TL08WsY3C9yDdhwk6NiM4jK5
2t+dgA/hCdBHOEWLQsIe62/E6VkF3SugGnPVMe2wi4St1QOFmYMvXkpRi36t0IlpfnNd0AZzMs42
P3S4lDYJKWhxMjTvhGCCvRYr6zghTmrFp5gtYBAIqGynnKVpTj4X+lLnu+RzwOIKWPbd5UtGoBVr
qruAq7ygy3LxHoeZR7xW2uqLo1PEKo4GPwlBx3LhZMpTwPwXpDvKpKu0U/cLGvLaI0LOnclN1N8j
+aYXIkSKBQy4sbFQPNJM+k7J6EbZsT0UfXHiMEMzo7ujvv9xoUYaTvS6WxVlUtCwRAtfbDqXh7t1
GR2sotMcN+VRUgRnVNxFxwRcCTxJSSgX/KuRrpqeWU4DpC0jWFkJCbTL4cG3FWbHi5ESjF17LcSO
FV9vviEojFF8dvORr0H67N/C5DZqo6VpvjLHz+MuaJIuSasvN9z+/3HdZrGbwKqu2FNLDbtM9Ssh
267p6Jao3AiQmG5Pl10MOOKlqG0Q8BWkEiPSEuV8lnEY/ECHlyvjHTsKV+rgdxCBaQiVH1YIdnm3
ttRst2/PT1xbJJR+hOWuEJnUiUxqMa4Z7gLL5m0X/tQldQfe86IHsqBZftBl/ZGK0IYRlznHGMIn
zkL2rFDSNtpjZcwFW+AbV67/rEfut5/Lqzml7KGY0cWfV1U2rQHEons+z0KYzk9JLuSMMXHDY0l+
3oBkKXx3L/S8uZs1qubHfm9wTCIQH2GOSm7i2dh5v05lmLNY9+GEimYEZBZ8nBsBrFghH8ktn0s8
uV2XroO+H0UsuoMlKebhNSLJjDA9voVDGHN6mPq52hfHaBvlEofRqSAQksVlFX8TtAl/yTnFTJzp
DFSPH4Ywba+FE03mCCzrj/xVD88DfXYe4/m555nr9xnzlFmCDL3w/PtvhRKjvfzjjzLYR6Z6Acg/
PrtXm39yxYZQPtfuZt8Gy5KzPSAOdEJHf1P5e0Fu9Pkg2ES5YwewjoEKG3CdmhP6gAyf8Hz+QfNV
FQ64RyY5556gSoyXYSKYzSBDJeHmAIF3QxhghKxDT0TxaWiWr16pKiJpGr0k+yYQ2Nh/frT9z7fY
4nBTn2HJzOe/J1WjLFHVmcX3KnzIvNzdj8IJ5m3NYlhAawtw207WaYfLU85vcz3AxN5JxUkZDioI
ynwO0C9v+8fANwnQxtcAeybQhn/hzBL1Vw9hn1p9DnfcgAlwsZDL0dg6rPy7R90B55X2kJE/X5Uq
ZEMInwNaEaHyJL65tXm+nPB7GeEc8XdRyyzlfhi0Vvyn5BlHHPQh2+9HjNQkswMRJKKUDMbJnIOW
TyETjv0n2H/8mBFCaZPddC4Kxwc4egh6S6Ufn+yuBmNQZHgKshJrqeAqj9spfhR0USaGDioLa+rz
EJ1TgVtyrWPfuLXL/lQB5YEqMjtQ6EVx83hpIc+HsjHdMjgRuOkhSFHRetwHfasWrCmWFDayNAds
6eXFaMnrSZXOXyVRQ5w2asrXAwDczEiuA5sncHlK3WngbqnBoqZIADV405Ttt5mWb3E91FAeTo2a
J82RBZY5BXRK4HDEKscUHdM5tvFFDuggXLTF34QD6ICE6fxCEJ+xDPDnpupasKoIwWDp0OPJ1Jwl
XDNsbqmCstY2e28AF7k2PwfVwRxjNjCOCXQ2rBUVqKmy20GuCgsj1p9Sqy3Q8S4t4AW+7hWrixga
WweAsneYmaU6e78zspP7cgYWU1zluPJu8o3W1uhWJN/NqdplNqVmggAvefIj7jPGCKUwCObBF5Oh
PhFYiZHda17j2nQQSucfgZQCWLv3LUFMJNb4n8il/PP5OjHD8ztXRp8arMukK95RdsEchHBiWq0X
10kkDCfWSm9go7Z0gO6GUioZw73LNW8BZBfMb02VuefR/7bJtsG8UKasO7NjjSKCx9EBpWB1IDNl
s9qHdV1RzvbOhELzCkLjd0pKRXt0oBtJcwSjzDzkhDQGfYJ+2bQOyu6qWOuZ6iFtIel0AopIJH0C
qBhHibapoCxQpHyYwHTsj1wgw2xH5lZxi30mFSGANGEiRGneLhBbX3JkO4s9CGaTCEG8gUV9Q4HQ
FeD0le9lqn/8DCwzrnWRYZYQKc+PWTBHvBlKJpOKVWkV3oDcyk/xp+tFloCjUH4/puZRB9L9cR+K
Mo3lp1vs6qzwebvuI3R5b5Ciksbn9ppx4HyOKQbOouXb/Wk7E7i+BDJmWLLzmIq8mlgdw7KxT78d
owYyToowYg2oi9ShIlyB9VJSTQmbBgJW6B498BpEn+IcNn5c9K4ARo59mJeRacR84ZnIaFMhnG9Z
lgtOwRYS+5at71cCNGw2bNp2iYCgCj12n8RwlQ06rDJx0jPKMqwmuZHP/iKkN5wCcsRSbVDz1sBk
JQPRwRRRL03xpi7QdXGBrFK3+h+sEYyFIfqw1gg9cqMxg0mUHpyul45M/UP0jWm+LMYPCTwcndBB
OoJbTqv6eWHZeD6Xmz9KrTb8sckOmg14OqQkKYmfy61T48QV9lvFqt7FC+6sV+r6YBVhQDhdCIOm
zMDftv12x8MIfe39KvVHoSJdqSUE3BXJP8CkujZAWkLOHZAqZ494Yl7TeaKgj++MZ8SBpMEwRajA
uWo+/r10ZxQPDlbzg6WnGukwYQHykbKnDPtI/FGxRA0GrwiqhgpwQJC8c49c+ML5eHgILjmXY/xl
Lm53IiiW/85PiKs9Ezpch1CruAS3t+EnJLmjqOhJglAQCl5LK79kMWDCZGIrSIs1uj+POvscx9mN
R10QV7eSJ++1h8YtemBEgP6mC9PKFumxQnaxlm3ybbRLsDvPlc6nmkvGLJ5/06De91RHCi40oAQN
FsnmRcnut2UiXBElr1DbS3W2N2Tew1zgq8JenAh3a4AblQUsf+jnsPqmKm+jqHr53e3qcP6dChQF
0HR6Ber8C6fNLrY6nf+azX5O8ZEtiMYO66OtJ8Gt/cLYTikQUfoMyos+XKVHo6HmQ9PPMyFuE+rj
95ahTt5uYy4/HBtWoplzugMlSp9ftu2rac6QvBpZF8qcgIYrmRTbA0revNGSOtg4oSaQiUBsW4vU
SZN/Vc2UB7mgu0PZbn8KBVq5VArzq98WYU/TaP+kyzi5yhfYWgA99Hydo+9mGzeqDSBZUUA8ocbP
RiG64FZM60krTV8oAVIP5ElCy5oZ+KdpoVEPTopmewR960xBmeSKzM9k704cFQHYbEOFKqfnXEmG
b5cgfB/vxN+PMAcmxxPt/4soFYUpWMt/BmJIynWTkerJdPHvCGosRKg5W23udQ/+FqICS4htNig4
J7x85Bqu/WhnTDY8pujAv1qKj88lMD1SVaVsAtiZTWSqhDhAnnNrbeg7n6ai0eAhRS2wvJdy+Ths
nvqm1woVIp0L5f0P9KRCw6pAdZ/EoDxOjy+DccmUGbvky7gsRBUuV4WpwJ2LTyFBHnHuz8iB5Ge0
N4Mcl4FHIoytMqw2OFAbeOb7xVQkgPhhxBJ/BnA3gaC8KxVqRxIYFGQPbSQXdbJMOwsKIu3lw1J9
1Bp6zZEyJ+83mbgly1meuXztqthU8c9EGd20WexMrIMgzTd2KxZf6//WAZWzET49Qiug7Wi2xBCm
yxfK7CBK0p2ExgqkxEMJJGXNda0zLjWiKGrvcFHrW4OtSi8OHY+KmuQD8lkqWWe+I9Q2uorwvNrt
RcehUKvy2/99RSQeUasTEMYTtdppMgzmNoAVBB6nXMmgTqgYxFLUelvpd2cxyEMn3G6y8RYBmxjQ
lUur3kf4hC49AQxSE7E/cf17z5BzsfVLtWepuoMhAbkQzN9HB+tsgLUC4PgldwSFir/oC5dfP4gs
NWyB+8qo4mwwtDF0eag9eoWHS9+z6KZIF5Bco7gjKlvgwyAnRuJoIk+LaXwzAEme3fwM+dJeThE7
BucBLyi94xL5aJHuVqXw+gX9ICNs7AInETwh6lrmLhPKMwDttCZ2BOjVnAqrew89YaQGS30ig+kH
njZ52W2m7HtuJJIYoIjmJnZxUL1htKbjHuTFflw2SrWp6+C76A7R7WvNIqkdcm8dbhsimKbMZOFP
xKhj+7TUz+IdXUonfFkFNyviYyBbafc0wqC+GJjA1bACE9spI37UZT5wcpIVhHZl9g3qchY8ByWj
tpyHCT8lWfd82DAggIsDsyIyaA2Fy232LEBniI+uDAqbSfqK9xZTU2QIoSmfWmXgC9wBe2dvbyGi
OQyVInGBC6uNK7R5t6TrrJ0QVy5fVzlYPWlqoQPw01iCMjj768QQkyV56FMkt4f88A6W8hZsw3It
y8P+mDy4MPPE8vAq63+fvk9AT/AqAV9+4bvhx87EBhIJmWiArs4/zXspiyBoXvROCEgs8N0Xbuct
r0Wo8bJto8NMOCpnxnTCPfi5aaiWrxbE9gi5VoNGl0jx97SoCAK7yW2eZW/ZvUsGjw99L1mEkrWl
kfY6pKUUVZyzhlQQXHs68uIYF+/D/VrVIfzdNLpJfeCi7C6+wm2jTS7SnN0AcLFjFLQPgR0/vNbu
zYa6Maj3p9eaSYmmUupnRhWWvNV8Tzc3+iVTTTo+jgSAbNbGxMpUed0Ko1rO1CAnOJeEsG7XAR/V
T7NCM/WiRqxyJvhDMVKjhkRsFxLik+Vu7uhW2N1qUtO8i58IiQKI5OSpjWPYgT+y7ftHPZuL8R5v
QTMrHHlBD5SIqOU+cAk/Ka+RXftdVZgbGR9JkiEPHchbLEWpbnPVWZvNW0RREn/9fmYK+L9jr5MP
emHBGqJ+wXicjBMb9q+sOMMXZLV0Xa7iXztWaWSj5g1YeqDPIz5D4ngSs5srNCISLMZ3iDqKgc74
0N3doGzAxxq6rVWelJpI2B5jmt/hdL0oIt8RIL+aWMpbEwkRyh2GCwp9A88lbEavayw7T22aCmHs
YNueV51dvYyXvuruYAO40vSgEM3kL3EM8VqMxtRWEn+3C6bZ/FRWRiH69LHk7VpnUlz5ECdDpn+x
RkXgWKDdniiS+ipQLQQDtzMyjn5UJ/Q9OimEyfeZbswKFJauE0GwlEYi0R6rqezCzy8UnBZjHhtK
jdN1RXGqg6GnWenqzveCyZjV4ax7XYkFfTbive95vi9JFYkp3+M9+/h6JYfPQxq1XDgaCVvzv6e1
/p8I9OUCz2vf8aqYgmPk6c/rWBSOF3tO4uRLDWSL2ahKUZ/zewQ7gviQue5ylRdpyg4NqxHPcRDL
ib4Qsdtudz84J3lChd3Q+m9PPryyFgg9BfPdeaT51Oxwg/wS1s2Q9Wdvh41Xzd2URQmCpAlggKtp
eUwF4wNNXSAT0jpgdr3Mo2ovVThUGV1EYFcGKftjI5ZfemDQALgFq7oMxLjAX4xOvD8wwBGvboTk
kbZ8UEaJo+PRlQWC92IA/gSnlBd29YGR7vgwO7r1QWBIi1L+GSDtgz/XOgPXgL5omRWkcSl4jom1
KLOI8wbr+k9L9SN950x2/RS51VKgKZj9+8GdocwldHmM45JwNwq2K/60Vrzunokjo06SU/VUxl2y
yOQ4hxwSug+5s2N28GoZzxVtF4SC06/Rp4wvvQ49V9FRHq5CeVjpty5GVEf7pBdMp/Gku5pKE0CU
3sCSGfs2sOj4eST3Nsyy8hf9wz32t886HZzalf6rBeGXlAKolAEYc2BrgGOSts3H8OyrWrWEd9or
lfjwCzAFzHwNMA2aCJbxF2MDBUGplPVh4tffUzKMg+82I/juEW4a9GqrIxkS+8KtVE/P7JhJFD6s
OK1oQfR5I9P9QIXzydZ8/486dUXICTr9D9mkzpvwKzdVDTqBPf8mvPvztNykCHs9Am78074SMiSI
RjCdmc2LEdRtvZFDrvGx950sYqP0PK5qKBblaujHU+gtksnhNIQp//4/4cyKTqatkC/rMGtpnGRC
+wiPx0SQpikATniim45GYmyvUnLN81uGk7soSb0820stAzLBI3CJD+FJtXeGOSN6JWNTNSEw7PMO
0oE6r/FNRcIlXNw/28eXJCe+0mBiUwhIx0CKamIC6t+RCtBvzP5wUwjQcsP+abVFMaM2llmYwZJG
fNbqge5sArXKXycXbgigrIMCCoqi4Z3Y32XrpdZlVpzDsv/vKPEX1kNIG3Hwsb4KYr4HHtkkHGQU
ZJBgq0/wE+UbjQl0JXCMqp4cZuwdry+SsueSaEQ9Mwo0K+MoENOWKrxhbRiWjIMnw6OW96nXUfMd
vVjadWBnv4HIf3MP++W96E2nRIQmf0b4/3Gg/B+pp2WnmAlIFP071FQs8iTu1dPBPkp/dFpJQJpl
b2tTSQUMPc/R/j6BAW+nozJnMkl6VYmXKGy1YK5y38nnZNw0Ln5dlK8VBoMEpK6yyTxMNUmjjOXp
CdVRfcvMZquXj/SeIh7qieAhz9FfNtka+x8Tddmw7iBOreDaI2bmyx4JzDD2dJxbyraU2kT26kJb
JR6oAxlLLfvhCvWDYwi2HMGfJvxIRUh8hfI9zOLzJca9lN7D+mcUCVra/+9/ydqONo8hTDe2xYFx
nX6fbRMYPgy8okNCGpOymfKE+gyDapXHKB9z3R+Smu8D6Qvlzm1bD7pmQQAaRK8XvKFagqAYPBh9
PZzPvYa+kagGJEZuH/HqRh0uoB2ZBXcJ3qLzELLmFSaVMUjhmbdZDt2vbqBpxOji/G+bFVXk9llO
xHV53B+zpAxVr5EE0qymQTYtJfhOpJRRInYxXV7GIOlLT2/IrCiSGmjrdncSEE4hpRVLgCxSBlK8
mCdaA1dRFKLjj0pYWQZ/CwmmC7cQw7Q7bHSE12pFRUx8VO4oKTGukNrtVwa744Lv4M/pMH7U43YS
/kajESl91hUhAfAX2LCntl7H5EUhzMYsEwXS4yv0JZH/T4c0Zj4ZEjjboCIo6zjLdG0F4vTPf4Gy
iyRDGNewisAhB6JHA/gFKIMwgeWQEDBWQKbW73+YwR0NyXsr827/k8sZjE53A7MJgQ6B8CQ0ZU6B
my453wdjgVpuPLXdkdZDX2k6XujC4cKF2PYqNj+Leoww6wqQhe3+WXzSg567Os7QFNVWSQHg5DhD
mXq2p0EnGpE8TLpNFURVYo7zx4TZuAbPVWWjLclFBL10nFy7R/nH93ZQm9Y1crsLk3QbXPaqfwwg
yyeFzgOYJViATEcN/mbspPrtHL2wRCyp9PLiUJXC16mGsdgKKCfDkBJLfUFJ4bbSBtMvAP+4kefG
CymYIYm3dIgB+TPFsDbRQCGpVoAXzFK1XMS6Mo9JAEgJ0f0ZJzkzKm8e3VpA7xdKErz9Flay5+KZ
57wmoM6i+BPk0DVaZKtOriC/BugtfqYK18iQKjV1SoLSz37MnZP88nSmbUQ6Kh1NYxVGIcopNN8y
VUrnPRxUDWmqHUtiq0DGviyh847hhtGZHWzCDy9NmjMqfJQg6OrQEhU1ilxtrFPZ3z2kQzjjASkj
i1fvkPdi1LxlWDW8iRm8fgbED3ZfkmasVBwaFb6Xxu45ZRkYPGw64ktwKpWLNSpjG+6BEtIS+e/2
6TyL0zcmksFNLGnrfmFsfAqYR7JhfzgXknjQ4dCRKeSaE094y8v8cOYWlgtrJf+Rjqg/H2tyswY3
1u8g0Se9NXbLdEVsuFHhlUBVdiMp2PxxZyLI4opNqJK+1AKXmSMP8C7FieB9ZuJkL49y6oTlzHwA
O3tnuZPoTBluHx5Wno/PRqhZ3xZOjj+FkKYV5PqgAxEL5Pwezqlt9R33IvRIcwnFBBiiP86ajxoX
oYrAgAvXJ1i83KlngWHh2TvMFI+UFYPRX76YkQJYWe7SRFyyyXpKSTPJfN1/NJLWesuZk2zjQlFf
fMUNI1ZOTGirveuqvsDbE6vfvR1BLJHg5mObLPNvrP9aUqZBNScI2XxwXd92QuZwZVCDyM3m4MjK
tAqfan8xhAqTc5JQ/l7XrmQBegrXPXdb8LN2AzzWnzKXzK5fKqzH4q5OJQaWUr5cCnYm4KM50fHj
OWHsQgTfACC3+sfrACO88cvskz1mdqCDCcfnTnhb8u8Sd7I852CGfBc0arUX9pyS5mFYCMaBqEKl
sVNiV86YEGs0fqkf9ErYCaSilKqGp26zoN4XYv9y/2r1S/qBOlGkS49ZhtkY0IQWKZNKYJ1dJlPk
QXbmwfk7p7y5xx0Z7oYw8oCdQ1WuFQ9ckvvf5F8GD6mm1GRVqEz9Mr7UeP6oH8g2Fq12Lja8cQf1
cvFJVIeh/VtPuK5uY8yYxIF9Kg1D86dI5ZgEazaubrn3EoUzOzeRMUsT5pGesjBRHUSQdhL7+EBI
h400YIyudqcHgMdffxXU4Yg5M1JpvSR7y34iIGumrXeJTAR8Nj4gEgT0CNVf4bPkVY9B81lR0jgN
svvGGPgQZe+R7Zp9HIQf9yDE3znOWkh69CnwlX4H22Cb46P6FvOpqE44QEPn80tsqiQC+r44wDLd
Aa4RqEeUb4RpMxkvMTbmKvFknXkiSZnsMSwl8vTiHpaOqK4N2BlgXBxWI954UyGLYG+Qh299Pwtt
Isr8VZmZUXYGXGn//ud7WXGO6PRxXk9td8ehDEhJZDkiM2fL6nrvnvCfmCRw/wZEAcRYo76MIVuM
VSYlMymxLvwJc75IuAgU3+QhqNFOdJBcVZCih5IamdRT1F8cRlDBjerOVpo0uyBWXDD/AIernCkT
hqA4+E+TPQBru7Akp/4ophCaWxskjQD/kU+W1aYCBbn4Yiuq24GfBw7Pe+MTaXPV12RpdO6y/Dgz
8YNImr1KADODQSZZXHVWyPpxuJNu47ZcD7tlGJ2vPHcFejFRKwh9CS0Wv7szuFCwmcy73Ka6my5W
hZkslSqsbT3ti4jJVCaRSZnVmRhVZiZ0NDEhpzfajH5yR8W4QdKhzEygK1FES6BLl8yQBHqBUh0D
at4eU0XajB/MRdg4zCiP5DttEhuFewlIB0YDFCjevisRZlvAlglTmfzor6ymRYRXSmfNC3xwlLae
slNCTsIkhj0nywrXiOV+yM1Fz4EssK0m+jR+lfPXsgh0EGPHvPVa1kTmg15gGMRqMQT6hqM7LY+I
V8Xr4hiEzYHY9H4vBuk733Fu+cNJUAoYTDmGj/9J3cMS8kyqAFUdoPeS0oA/Fnqbcmi76pe+o3B+
HpvTb/Qp7tFM3fMg3F19XUDnwKohxJM/5Nm+FNZ1efNH+t5uKPO4M/i/0FJ1Nr0gP2xspxdZN85B
oldwPd1KJEVGOm18csPUThgn88qWKLwEbIfM2+bdGf9i0XEiKQWmcb1LUoSv2+FpLLoLJBQOLXmO
psmlwRi2+PoxTq8ftbHSMw9EfX2Hkdib+Q/+ORKach45VTX2aBIpX+3AxETOzwQb1Xkr7KmfVh38
LlXj7uFkk71pDg21/GGpEsU+MIOpAsLfjYa4Xb8Hp7aq+JRH8cLElR871K34b1GRUldymafMUwvw
dSv3xGmCczh2eu9HGDQ9RH1zXJSlG72jDXvtogdaEKObEUGLCrCABz+SHUzw4mfH9v4hOr6BMuyB
z3QZR2ubtDRoh9VNnTph2yTbxmKuILVXM+lBlA/e87IkDEgX8LvZfxV3pavz4FKaoPASzDGk0BlH
B59LUIrHNYi1upLIvA5zLoR441988g0yFEoDkpMZLHXEH4v8g2dhkLFe5bqNAXr08aBYaDmTnZ2T
nl1CL4/Yk1KQYDyXPAkvxGtOOZSwtgdpi18LXwhm/rrI4yozdXkn7FsetAbhuKd6VvDwZE3rgeqk
+8fmkI6RSoVKOb2yIfF6dMnKPLXxFFYVaEUr+ZpJHGen3ZoAbItQzrt5/gdEN1pdO4hjkaMFqPyU
CzmOvDEaXCl/8mgYwMq7Gn0VeccWnDobd1ghvw+QxsPYOVwTG8jM2gB/2Lv9rBCUYDmcrdAAmDF2
39kv/3vA+8IZjpNTvqJr7Po3h8gZETO5Sr3MXJ4KrjoOjmVGKOrHS47n+vV2+8ObdMqaxXTQJy5W
cayeoF7m9DN8dbDhDj4JnGlwqmprQZDb2feHedUmFtamOEDQ+QRe9dmr55jPN46xIqj1r0xIhvJ5
LWRNHiaKYrV4rUQsOSrpl8T2LkzGyDG7PXUKU5iiGlly+waNcormJO+xH0bHRvhf0jmJwcnEMjaX
GKk/qbWQEmodfz7Hk1Yp/QDEjCvDnd4jWwXAeQ9xzRi8GR5B9VlKtRciLrI12hv4D8Se7bqqsJBd
BxnYATT9GmVuV74pcI03WtDfr5ZCkLxJ++qeaavNTItCnyva5RyzYKy91xZBrSdJLW4ySjFjr0Ik
YhI9zltJMKGm4lqbK1w5j1tpjFS4Tywt20n3+GAIisY6VXCVZ5hDYaRTLwr0uJOum7z4tmC8mXGg
KXdmMtI3tgWJmnQV708jYEFCWt51nK+ERl4QLAuS3gM99DYGMFGsRknBtsysw3ZNhuAuRO49qZjW
y8l8aCDmRRfits6TU2e9a1DizIA8O+PRpgrJXjz2+tap4NGSrXNDgRVRxanVwYKY5T2cjoB7xRr6
vT30OgrXPc5FSUoZEau+OI6Wkj277nBwX+mTJlXk1zOv7DT0BgvVDNAGM/rxJ4n2MQ09SpMb93Ju
EuLBVyGjOh5znWWE/Jl86HqQyqDrMVqu1XU5WJqOSrkXrUp/SF+uHt1Vozvku0NFb9PdGCJYiwWN
2kQOb4Mna821cJnhTw5kBDEeLuzPFSNNndTCkAXSgAdnUb8OEAIqOkjX2veuY1Xg87++d3575bSz
KT7xR4wIrh1RCsaIttLbmqXABpChploDGfqh6Efx9cGEaxusWGRci+Ubcgf6J+cKrzlMTv8B4SJ2
8MfQOiE0uhcXtaZQHf3B/ZPb801b88cBMFu+bJjXL4DMmdSQzajxtn9L1dyZZ3S4IpUJeKyKf4w5
+qoG+kRAkHpkXPUqr1lzGaQkmBOXK67BOOyJnVwPdp+G0n1czJrTL25JQosVe0vg3yLn6DIbZvFv
ueasHrYa18u+lxuNtB7Wd3rcPLLAFX7HsfSYvKIIkerKjOq9kC898z/hElymnxN5EothrL667oCD
74Pg1BEscMbJeqwAVRstkn/NHv433dAtB8kRkuLTwzMREyQYzRp2w/NJlNeFIjz7ZYSuHhKEi7h9
TMkXIoDCkBpcqXk2G3ZBGtm+CuJgzilzLkC8tgmfmpcot52maSa54PjFYc+S9m8wLQAEZP/0h/AQ
FwiGmLBEnB5j3wtNfepDFQOzQD2OmI/CqUBLsZsL5lzDqE2au6DhbGA3fswdNkgRMEbLQfKtYWkO
1i64dtrbFxFGf15UA8J932c5pdznO8uD3jnonmFWkDlZH+rLx+l56BjBXngN2oJL+mRhMSVGthBh
VxyItSCjpwXvBz1bx5Kbq/CAS6yPYkyvUNw9vE2kTZl3Mwjja30tUX62kkVh70hx5Dm9B0B9pfj+
GhP4HRXQeWGB1rRxdechI8OLokKf6I46oNPRRI2vGkd+Z3P244W+eXyh9d4Ae7/72O82QYmM+Iae
fi0qAbsAV8zumwLE/STLmGzxehTrfdmAgg6QUadJ2N0pUuBJ52hKKDi9Z9cOqcSFKdNjLMQnQMap
N3c3GsRK1FCru/i4hBOxngIdovvcdZNPGNTYgXIq9yHYomOSV8a1d2IPxHtENybU39s54kHkYE1b
zcbAd5O1/GRCIcrerNH0TNpblQfr9BgXK5+3pW6RaqCVLgyT70qkqthI3Xro3B+RToO6qeK/XjT0
fF6acNMQAY7fjnVHsPvgVuq4xielamkUKku8MNYtmInE8A0BJD8IQJHWY38+4VmzBr7M+G9qY32r
rQxNTfQm77NmNXIOD5o9ltfEOWKYy7kZtBWbyi5Ldo5hYUW4c8A1iJ3Sh70gNnB+3UmlMqpmR+HS
mkf5MqBG510KZF+mXOiU1aYZ+IZjKFN4NK0WzJe+GEi/d4Fb6pKbAv5mzUPZWa1v1di/Fk/oCbT0
rH3ViRC27Mzac8akIhLm4tylm+ck8SglnjPYPB15dLf6kkebluL1TO+66UTvuMCpvjAlJfx4uu1G
qN92yosSgx3ty6ltH0XRrKW2o3d7UEHWCOnLxVO75c0KsS6sKnpn8y+b7xtBpGuB1XPW5kV2ayEv
T2TWUKMs6WVS3DFjvuTic3a2vCL8onUtWa3lKlz73KiuyW3qYImldljMSEfGRkXagQOrp0SABBC7
BqAnd8GHsYFiqeTKp6r81k4dGkGVO6k/qZUjlBZJNZ2OVtctuuFC7Bgp1429+zj8AqwzzNiciXc6
fsRwCwV/MbL7cq8/4KqFc4S1waS9YwiIoNQM2OABA0WbL2gKQOsbEyaHQf61I37ojN88DxdM2j/+
DLOF99GWj1/aI0/byUyDjVIWC+f/6BLyFamBmU7Dc03vhVx6HSXbJSd/OhCz0bTOwKaKijyyQxht
PO1EFuzUOKv1V1DpsUmn0J25tD72caAU/rDzqEvifgSepzk1K7hJCj7TKEO6gh6McgLwZsOw6xIp
xslvJqRf6P9erBnTFbW7ma/a4jQLCXsy1wm/9lAN0KeAUxgp6oBZx23JkoG170Gm71Sr2f1nrPqt
JZsN9dk52+tQHlXt5pmBZOLeZiLJ7GuShvgtOB+5WDjN353rUwXLdrWKt2W3dRQFxMF7ZYdy6dpo
rQcNyGUSgMKWVu97hT5UXrhcBYp7Dz8bJzooSW0tI1NTwCMv3CmWIp55Yp36qIe1gARruOvH8E2R
oHCJYndErjcNJ8N1VcdxM5kw9YWPwL1mTMW4BDQLSV97GOC9NveVkzz9ZhntNNW47F2sj6eWFIT4
exeazELkAhL2JVuh4uVhDj/Id+90L4Kiv3jLN7atoQYXDrgIpljk932vUGEpa+0NgjNhiVzscj2n
92CxP0RfmHVSHwzk/oKqZUW3haeDpwcFP2NAMUiTUmGf9cNlDNnsGEuYDl3Hm23hj8qYuYNTx+0L
gFZV77YkqDFWxAMb63NutJht6lRE2RI18as+ELEk3dxSrVWflF4f36To3Fo+N/1DK+iVekkEXVMz
V2ahXie2MFgM2WuNEoqBdI6WUYAX4XtpULUmy0tDKo+udSewG6Gy1j8MNVCAnUJrwMbTXwNFZ4Ng
+yQ27c/MpWbLDsqPdArhoA73k3fhIO6hlICAVd/NGhSEti6cFpKavxUxgPaqUDNUQrJagowZrlcg
zvC8/VJIM2tYr7xzGIFIOa3fak27gVjG9ggA1XMGAiDYSeH3AuuK01PZmWySmByphPSs+qxHpZDu
EWaJgMXVky7nvKNrt6/3gj+7iTz2bmMnotFKkXv53rSchDIbtQv/lBSB5v0ak4DA4zFAyxec/wLu
w0WGxNrbYygnHm9GJEf4jEdPIE6jYNt7kV0J3vuGsnSOAygpHhVP9RLpUiKv1t8G4DzM9zn+ev1y
H9LUKbHW+t7COL+r1QhEGiE7c1qlk9oEutihwM8P0i2l6GKW4YINg8BsSjuuXxZiUrvS7K79jD4V
n3eXEDxleXeyEhFt7/I+l1zGrGhb2UJE5aN85VAVZ8akI+OxgVBH2ssdOvu8zDo6ePhgRqLSFqh6
ngY4i+beThBbzM4oIqera517VNC7pntH0/wDBTzkPdZ2z3bocgntNEcuzBoBBcRdaIr45VHx3Xij
CwRCoKJwPGvKsCmlYIYBkim6T0WZroks4BVTpDeXqTSD7VUK7uhZ39tMqg/pPJBXl/LIuOIDeI7e
GfJLvx8PZ7i1/V64HxSXMiE8LpqWExzoYSyq4Bp31YaZix7ZEj9cdxG7h6KzmgJtYT4M7iTLGx4G
6YzXwEL6qYLAeQdjg81sp1KPawgLomaCeWB+ZgBxFSevj7CVT/81NNdvWD2QIe3kLHYhAZKjTxZ5
v1o7Op9W0m49yD/B06InNfpaWQHv/S7zkx2DgbOSVk2DdCH27cqNuTE9Br0kxDCyp0uFjTSrQbxe
nK+6sCwj66InnnAfIfzg91jUeBOwO8nbsAYvFPCDretJXdZy9qtvHyFepcEXFflFH/eHsJvpCVw2
pgxZKHAGq0+YyG+hTP6YsCtlTH3JEg913uhFnO0JAOwnEc5Ytg7zlAZi5ewY8piaT8jnth/7R6RR
qtbmnHJPx4kFR5ZEN0+8KIFuoNBItx6tuj/8yk9s127FQ3Tg8SDpEsfyYfqkcFChFNKYW3Dt+pNR
5Ek9hAa0AQLMY6yEsXYYfc9o1IaBoFgCrNZDH4oqVf9ddqOjVsrZnYeilq4Hzi4+CvVecEAwSAJm
U+rA+MXecW0RtMKbu1IHus38RrLoFy7zMNzxonj9Mvfc3jyxsGQjejFvq2EC5KoOlTSKurml72Ma
6NXJh8NM5P84tyhGGsXA+Awa48KP/KRkjYAKDDML6ipHv/AobpEvas4q2yKx9SVbhqb/YMzJ2StB
p7it/SI6uoJTt0jRzqE3w+SUgBVE0i0RTWJE98+97onRqsZCFykeZbhNA1qNJhSCC2dLE96wX/K+
BRK+c2JICHrYl9w9vUGUFVFuk2fBw2sMv1WeFDxfp5JQHGO7b2ZK4TwjyrgQt7vDRPQwYhkLaRsd
CfiQES9P+nLxE9YwlcmWaqAvNp5f6IQsrOaH/eBoLEONO8h32zFm7oa9c/9e/e2rLZeL0DzSRe05
bTKJxvtvwxoqRgnj4ahv6+YUZaoSlmRQdCHJg54Woq1sZwxB/rJ2cU3yWkHDF0Q31YMvRq6pBLA7
VfIoJXtDtjMx7zrOCuUP980EUPx5FlOgHEijHDDloRL7lhyHyfTKZ5A2xEh0DWNYrCkXI1+Q7Kja
u9UX/MHMRA+jZ16UllCRFJtQaJ/nU1+gfYXyLsPVvv9wvbWqc5JlYhwjMD157zyXsY+YiiMbuNAJ
+eJC1knV9GlSk/FtnPwdFUeBq9aHWTk5t6hd/6ObL3x0gyDRLbaRum3pLr38TlwxYAXfYDb7rN6w
50EO5WZG4m916OMi/uHla2bRcgg0qrztV+diwy2YSBpak4lIaiiYOfBXPyzNZ3bi9Oa3qcN2+6Ob
Me0+MELdgtmiTfXiExz3mCOUfNfM/5ajxdVlngAJzKR5tVlXoe19oj/zD8dGxPWBxnT+I5m1eiXJ
Aq7fGmKHMCPabtM5iFcafJqW2wIR6tc4d7XiYsM5haEYpa0pEYab6112F2E537SWx8GJkMkS1NKp
L+TWx9Qxcvq4czmHZBupRs3uGBxiX7DLKsw19Wi3Lp6VvMIarkidW1axQ9zRk4wNltDvM6neCvfE
iYKrugZwdmcYVhx8h9IG/t6XGLvMJNgBHxsANGzcckpdJ4uRy7OJBJ+sTFAgKCLkgFKwpeH6BPaT
mvqcemzozsMTST25q3qnu1U5PMEapTv6VsGRz1By5YyvspudMaL/F5JUrkzdP7ublMcomkjCf8uj
1fxX0+ThMpD9P9Vyf61mG4Xt28pR5ksDBAfJftiHB1OO9bJmeSxihQmpt/lzHpe/otkrE4IVbwxw
In6SSaDVyPxdlmWXSlG4ewEjhx+deXJoyGSwZPe34KYrdNSRQnCPvwFFojfJhxPVcIwQ8XTpAvJC
Ti8bW+pe/7RvjB7axu1eScfQbrRKxrpZFlQ3M7+vCN6cnasUCn7xExCbS07v+eZyir1RJFCcIDdB
noo8ATKaly58oPkvH+WDj0dSo6qTevh/NW6S8P7aI9nlOtnXl5PrqZvoeaQNvfV6VmvGwiUTBfHO
SW2t0Sm1pALghjjLeGFvIT5NuRDx5BMpaETpAFrLT7BtilVxJYAMHR7G4iMFz+jKCMiljw04Qyjw
GhwQg3W+lrtazJm+Lj1fzNE+a56g96W3vctY5rrPgbhVtSrhCsC3xCEi7b9mF7C57gmzO78YE2py
bKsXNvSPuqzp57sywtfClosKp/N7cAluA+7tM4VWDCuNAMQ9TSyOWwOEPzLNdeqKwrZvFV4MnWrt
svUDmeyMO4fm5WMPFvXczBysQuQVczwsiECYUyl7GhvFRYUoRRLHpKd3r/kI54VlvAPUVqaWwko6
B23HBIP9YH13tRgOnaR2qZaWP5SqpeO4c1zLDybJmAX88qWkkfxZBBYiUUT2yb178tkPZqQTK4Ir
H+T605ip6aZBQw0nV08iGLXIup9hCWoIBEkxtRR9VBXrV0H9LcU+KxlInYb6qD5ZP92QyTLgwXAn
5zyEgXj7EJJc1P7k0qKgvtULGg4+uwR+UeeStGLwBib5eWRTjZfgoK+3ESsMOZ7SLom1AJGKTZBO
sAuvXAohdmn8XEoduYAmacRh492odw+Fz2RpaH68eITb6ZLxCF0Ub3jeuB72XUm9DWAUfuLo18fm
RdGy4uiQaDzMe2ENhMbAXHueFDiKJ/hFvoyMV9Sw+KDgrbkqL6JF/yAeBXVKBoVvjBbKtENlwYOk
ymc1qR65s6HeFDHYTnAcOJwKrX5fepAwgi0RmOPBuI/qFyfkDZL/4Qxu7GH8f6Cre0fTDTsttHJj
bLZ3GRWmI7N4ubqRWfflHkBTMbyjIuoLlqk522XZxaLYUk6KtQpqY0iHx2Tt+VF53iasX/dteIFv
8TTS/plD53L9EULBG1imuUq5zZ+ZywqRrmqHfk9FQSQv69BOS0+NJbtnCDXrx1UetjfL8VyPpXJn
4x79Nnwh9yUX71g2f9xIUjDmb9DIR1lbxEQuH43vkjySA6Kw2J8t/g+PqzjaX9LzLXosb2sjD7eQ
V222Fcko4RDZELrkARovZHZr5Pa11kR1fquJBB0CIx4A2Rj4gWNoujNx/MjJjNfk/YeqSs4jXvZj
mbZCBczJ67HVp+sNHJMty7Cq7xjxBG48r4zlv8i7nq3pHPVNKG8rFcIRZUIouyLinB4+IaFj1fq1
9gnlHMavRBLaAyVpqNHabKAvFbdxDMYQQr4+SXTtiUIlabl0sSmSrMKZPslJhmtxWpJbRfOt9Ymi
+tIynFhOqUJiqI/gQUATSCPG2cIvxAgLLPav2iJxyaWXx+Zm+s0IL3p7TmNPF3ElbJTs+9cEtnFf
LdlxRI35bWDoTmKY9I/yO/0i5A31HmLVrK9DwDVRuMK0XVwpSlLLYmYYucKeSNCON9ikRJtEbNZR
puotnMAdEFEtQCAg+3kBd4oS0u5FfCTNe7WQSu1W6iHp+m3vZjtzGfhXEnvMChTIQiNurepGebO4
sl4SD4zbIo6sdKe3pYF6YkXbW4SXQtjBwOZ9SqJGwUycLs0Zxpg2JI3/PcDqJZqYRaHvhxv0wM78
qmMSxGtWg3ny6KASVvpNrEaL1yTBWGCtgLjUa0lFqfEyeMbbyMd0DNOZ9BNWrPN0DYwjvpyNWQEy
/PdWhQdJz6OyEkbihAuH/D6qTp8w8PATQ1YeXegR2qNVBtrs+tmJsghfiJc+wCTQicrklvfgbzbq
e2ebzffAdxVp7YQybidiO4cjdvx6xGTmsAYwZne1VObAtKCa4zadwEKvpOoEKuqLxUrsDoBWCEuk
yx9JnPdHXb/Wcix5TBjsylJwZriBhABXpPyFvbjSYPBaqMfv+FT2uZGI1MxBPZvzZyDsrL19NK6g
Q6GwEcJY+ZXKKnLMP2Pf1zPpMgFwqKu4lHkXiNf0cvTiD9g5RAGpNi3U7ZqEMEUGvjhzAOy80pyl
x2eiKgbntW7Iu4J/oQw2xfQ0dRA6bdXxxAuP8XPXzgx282Tt/2E/7zSCfZUs4K2UE7JRtDM7C4in
s2qPKAPYP7PE9sBbdKl2dTT8txHRngma/2VOnrc/heTRzwFPwetcqpK6MS9KRUbBHHsjjKyfxPdb
UeUxkTAUEsXuDgmpWWCcfE5deQ/dHjsCFPA4lJsEu3XioMx7pLTJUnp4wDxrHSmWA6v0/xXYwqJy
Z0THiUB6265L9FjcGYKekkqQiUBwj++33DIWUwLmmO5QrdK2sCrIlUbTeAlJsGZF1SGhjajsmIq+
lgCnZ0hU8Xl3QHIi/xAynGL5iP5o9/NQbVsqvESVxmrh+3d2Joqjr52Qadi86mD2T1T8xZwWHWzA
nJsPZZHsPKfkKDKR4j4VZVSRYYZQXz7W97vDBbL2slgIJiyAVktOd89UPnT2pxxCSj3pTQflcGL+
FHL09mjXk7fmR3xvIifKQ+IPAKt1ePsVdqPw2jgl3Dw844i6wf3QIoCu1RjtLq7/R+5H4sOdBMfw
jkqOtKWEmcgz4TisWvsg0gPaLUmRl3tbIz4lWQgGGYBUzJKwC0BVNAF43oSqYZQgzDCjfdlVDUqd
JnY4jhDeU90aS1RYYTeU0oh/yuA5x3fqGV1dbBHTJSF+GtPVKuHXIrngKMp6YjtdgtSbVHspwoLB
b+kxmPx6iX8Sex5B0aMhOneebh1NAJgsT/h5aIKfV4AfRSfxsRrvZHPgdX1z5LBGg+9v4MIkoXS2
JEQYWEbXCsvN6+CGte7abWex1AfLRdOs7RRq6uEG0vBttdtSrqTlcDpK/s7cGNh6y1kEfrbTM0Vm
WhEyPaLQvGC4BdiNN/VI9AddSIVBTjYt0PrNi/Vxu1k/S0dfyYPCTxu+1SnZoWitncoZ9ipHZgKg
EO2RiM/lOLlh0sSCA0CHd8SmwwNKpk6VjatGmZYeUey6ugc74J5ASpJ+pyOkjX5m2OG9xNyBnmd0
EPyjX9So3zDwpaDQruQ2nsxnLINelpUIOPaXrLapm7BFcfQp7ktZyQ38kw5hbJYGf3xMjz9BrJOD
qQ9XvjkncUV2XEOa5HPxTR5n2gCBZpmujeJ9f47Cbe5oGQG8XEw0WUSXkqj98ueEzGK38j4TXNlf
BrgfDvfiyZd5h7ZhcYg9E3rX8pZg4hQpCiDu5IKEOCCGfi2FZ0SSPZ0FjHJBkYP2+aW50532AhBJ
BWfyBx1A3ksqTx1rnay1nYLH2o/7M+C5L18xD0wnk+zHkVughbSwV4VQPSnGSLzNz0QURIRzuCGd
OkcDB58lvoLon/4YWvN7CfLjh+blGxjq9O11Cfc+1I8mWsg/qft6XcsfOpuAzS+RTkoK08NeUFY4
R2WGkzOiMzcoQGBsfrLlqYQ9ADctknxbbghaYZvnwKz3GvqninWH86PbO05QVkoTNhbbeR5uO4aY
KEsF3la//bdWUf9C8jwFUCeLWgBur2veN+nSL6KcO4RZkxlEIQIN4F8BbYxn9n+e0B36rMy4oVC2
jZMkC/2u0fMMq7CFsEKqj5NqRGJEB0A3rwJbEXnKpLQQPAsxRgqGYmFlDaC2OlXeMDqogAGqrPX+
0z01b4ZqD1QNisv5Gc3IIfBYMR2+Bx1z/l2Bcv4Ijz3BLfXiZBs/A9b2vU7NmZtolvGIy2cjepO+
hTW1/UGp6hxkk1Jk58+VkhZauTBVHXH1ymO1KgULqhTQ73igTAeSSgkT0sCTXF6USZx7QSwa1bK+
9KCfNBsOEy4lbAaIkmEFhsuVZB8RT/r5kUYXGx8cKeBPA5Z3fBTo8VAyevoG9NdhNOX2cLCYBV0i
6U+IhIR0FTLJxqsn0xacbBYm7r2m7sJ+WdUffF+nh8jOpBRfVWN+hsnFxrj8p5/ae0KcYMZ3ZYhH
0FJYWgYxPwOl/j0B+PFdJntpcUsiDEgGnjSCujKoKEyrXGg63jUHIcmteXPRmeP3EMHZpZjj4L6y
0pmJilT/SQaqdlSu/S7MLnTsLS4ifMQR1De53TkH800rfD3T/O8QfT8DYTME+opLg8zzJPxAF0//
MKiHGzoa3VrKYRRjwsSarFQTU9CpYxb2AtZU2hQVgd4Ow58NGxyeQFbEPLXSschJtDaeaioNheRh
vlCRcbDrRcApYuG4hq14YXwrH6HgPtM7eXJSo8WKu9Bq/v7TlVfijg4voZl5kBmYzcpLqARkRD8q
w5JeY4LVyxXBgjQEmLB4FC7RCh25dGEr8MnIJn+yQlyPos+WxjopJeNHOcmSrDHRh320lQeX7An2
I/5YMMOXT4eRf0Jr8gmE5yRWUKR3x4lUAtuHEPN1GwTr/oVhy8nfjxzsGZLPxqc87xtc4kuMIIxR
UbKzsOiY06CLLU1HAZ70tLI2LUS+vc4sORhrhUp3xXGUrH5KcxeHoWN5CJZBlQQokcUUBnlQUdYk
GeeF+tNIDUqzq/888EwRenrz3m1lX0PbcKvlr/iDXMn1WQrIApovXVx21LyFOvRzgAhAiq4k6iL/
nSTDDNxT7mKrmlRshk5rq7yOjsYwxYkdntJHxCwg16Yricc8MLwAUPhDL0buDzIbyYhOwTeNKGz/
+wXJOqg3DHWGQ4wCLEQI/ZnfjcOSUQRIMkU1ItAgJvRRkEt4hFjPz0fz9+lsyTH/CQFs2TxZ9DtO
atmxI9zzP/P2as63u+TA/ag0zeOVqGbQZla6xH1Vae/gJXnoLukh5XM8W6nD6oeWwhrelOeoKW0n
7FeR9ejBGSG7e9Q4l4+PgBjxB0FAQKyZHms3UPv1gYxf9L4BO5YmAAoTUI4dPkj3BBtZLCWbAs7Q
n/rXueDPfaL7+Cqep3gPfILOrQSZAxg6rWROklc4Ahy5nC+qfDHnZqDjkEi4CzHARIcCzeNf19xw
KZd/msM0JhEPvoI67Utk7uIFlZAp9CGRsPtzr/sPWBxHcPbYu2T7OQgsHiUgnmO8TuKpNO8Fj5DB
cDpFDS6WIdNKDW8luI2LZA3GXR/lPjdlpNDK3aRM1t10LmatMKZXd4pj6msCz19mpckMak+TsWD8
5+n6dqf4XsH0CvG3xsnbN4sQR8iphcg0kWp06NbPoDjG7DE5qqs9mAsxkxabyXmvg5to45cTvWxp
/WuHf67G4uDyigk8dijcdL7xGWCLcRGWyoDzbx419qPPWlFOFlA3clP/0Ch69RsYN4cRSB5gdX9q
kax1eD7guDL9y4HvjEGPVnPwgXHlMR+kMEFiv79UJKUMMoGSCGuBZFrVffQAqm5gsaA1TlGTZrrm
LhOvUwQtGFBSCuFylixMSiRPtTCRTSxXSi1FBcdtIhdCVqZ1JJ8ugfvCET/mxo3hRuAeTm3B4n2N
lox9yJaypbHxRRltozcMqwAfW86QG/WrX/BYfxvv1bISDEewp83Dfsnxb90qVGojwmkqKU4EECbQ
Fr1UxaDDmDcUO0mq8hVGLiJECuAfXsvGAYfShIX5LRPM0KqQmVJb8mA+CnVIQ7UpWBQ4PAn+6l1E
QKse5tBv47gupVuBJdv9QlXKju4+scNyoXEujonQFP7FI5HjehA8ReAGzKhuuMb366SGLINyuNJy
fKw14o2uewwSiV4g2cvkG3TNmFyGx4Bt5izWPXDjHrxN+/WXhK8znaXUv/F0aVcFNLgRwDG5MBzI
tGNwUIHUeuCiyD9i1lOJ7BYP/eFf8LCsVIHfPxmG6Fo2/l98q4GyMLP5E0K24jCju/HtUu4+SWIu
3UafonFL6FfWJm4k4lYJ8NYksRK60wc9i6TqW2P0Q7h6l2d+Z/23WOs8PWVlSX6DSzeHw2Qma2k6
+KSLQOOtPxjMRA/YtW7/byC/mC8bpD+FjW4XK2yebXWNDWVmrR8HEOoYsGYoWoiixcxTcwMfgXtD
4FhOQnNgtGL76D1SB9E1XVjpODscLdw5oNLwt/rCLeyd+06XOSupUkfDaAW+C+m9DgHb7+75xDHk
Vul3w3qKeGutUXOrhJXiFI+3/VqDQUS+KqYABuuNoY4WoSqTsbT4SF9V9j/CffwXqRq7NX5AlQhi
2tYTinai1vcPrccMJEjT4x15I+fG0tB0Dehiz7tbN4s0sejGGWM2PBoxTSaaoDRswi1ErTV7gFA7
J46oOA5UhkDD73Q73VB/vHMAp5WKKpocjKcLxXLeZ814OxUD3kANZ3ABOK0jpuxxKCQLkR1lWbv9
cVgIiRPG3TT+90XOaYFGzmzup8fGeir61arEQJyk9/zfpu3uWyT+B5XC9j8HF/EtOM0w0gcTWC/O
7ox+0+aeR/n7dbUx2w006JTpwl/ta2mgrCK6wsfMOFC8c1VzQT184G2BHn2mCSrJpS+fQg4eJHxr
KPp6nl6ZJHI2q2BwLuD1fxIdprShoG2P/9CSjaRSNw+RjPJ12T/DlaEcG5zjOpNz9zatTwynHDfC
Z4XAU+00RAIwKJUQXHIkqL8kkwZ1vljDaAdoLohQLzq7wIpIXn1KBRaqPTLyfltuIcCTb1X2/UJX
/Rk1Y09MpWGpD4V399Ra1tw6SnlTX4fRZPf/o+p87LjqQQ49xe1Srjq6N4Wyq20OkfgYYjS8tZ6e
N7Sc7hpnR3rpQRyEUMnNqhn7wivRsasB9nj2AemwO3r9NK3xMUvorF/sPGNhlSZT5qyMS/NXKGSL
hC3iYuvh3QVXxZ2+FcELAVN4x4zjXOiB86LhqXJ+Wx6e/4yOCjoTFN0mA2wCaT1762wqy5HpnaK9
CPnm0Vi7nFZsScVGy3AcRjjT7OrBv0COEjopX7oXYfIq2pLDT2Zvj3pTU6ihyCp3wKVV2noKrKdt
G+5Mqav88uFgAENTrY6rfmQ0G0y+5tWsDCdrJG3isaT3ql3o6JKXtkeYOZ5Sw9gu5TWyU9N7B/8K
Bx73FvAA6s8ypLrh+/0e8GRltYtqcC51byzigJb8MHCFv4ackWJgKVZ6PTKaERBVO2sL2H8GH9GK
OgaDHGdhoR2mUOIWwwF/RZ4RikzrmS+JzkGSI3RqhtTzE4H5MQVEYLFe7A4wMS7H0yc3lGy/FjhZ
SfW3MHzPY3ImhZs3UeNHQPzNrRXfH/DPc26tBgajR3hGU/WCkeCgO8Zhusw6t0vVqKV5N+c6aCP2
jkKFROUtuZomxrkGBlTWw2vmfhou9BTXKuKe8B2/TTCn3yFhX6QhVoouc0ElsbKY1ioY0OQBCBo7
g5IO80n4f2mGw4Rd6Cz/V3fMI6ghB0+M7ZoyDPAJQx+PK+kHhKUeVG9U6jU+uKuaAokZR5Wq4xPU
/3tOgfC8VRSN6EVAx1EEyK7sJvELQJKqJZ2CwqjtSVgl8oAo2Rx1N6jsuIcvVDqQIJrWefXToapW
WAZCqweDtjq4XGEmDXS0lkdVYSNWDA+m2R7fsKWWRCERZ/E5D8g98nvho1dXSTyr8D3Q3cYVLqoK
OV2ljEmUANoJwHmzoiRr8vBRPTzmI1uCfwaKHzDh92DTPeyzZkIdYucJEbqZmqXFEsQRb/Z2INZo
+H8cxg0Kuu8Avt1+rqGma6GljBtmv4C9+o9ejT4HVIa2jWRwbslZYqZ0p73nvCF6GWMEwOaUWArZ
FPWjv021UGWQYPCfYayeWhq1RBHvxCFMw5yS2wUWAmaxrph+en4Lo4DUvG4B/vK4loY4T5JZLFYK
BgQ26/cr0f2JSyZs92Q6klJNg7fzNIVd4sAAjMQXdhrGyV6+BcEwE7u/y7ZY9hcQnTQlDatXSNyU
bdze0hqnVgOOngTKGM0hkgsVUyGf9Hut6tiONkoIWIs7X1TuAm0e1Y8c/xe5oBhvvAtm5xl5/578
tnJE/bU3eIo7SdYXYKXLYiE1N38kmzgo3q8EIuGalCpM/6oYiZjwEdHtr+nZhTzi0RJtLQeMSLre
mOoJO2mbOXv8/nEtIkOwZbj6Nbv6XcBA9f5gJooGM3Ygba4PSWpfYxKFPqC6UDH5DDMkAnYOplpS
NBaGXpLyKKexLTTMJQ/r64hKIg+pHIcY9F6H/r5GrU6p+He0nCDghJKph879Ihqy5C8QhlzzlfbK
XgpHjDMV/55EExYGSAH7R4lkd0JOtx8bYjLv7XbZrSo+siSSLMynV/lynlY7wxkvS/F8N5nHR3a9
NzQ1n16aYwyEybtmeuqqvRfoN84ADASNbtpBIFd+xQW16lmjkrkoSXmTxtYH65zRhK1/KkJSlAnD
JFvDYmxUNGR2RiGg5kK7xpJoZlT4ku4aVa8HkBMsuPZlP2yZtpDiecwc1sNPW08unQWV2RWyLqAg
82TnHPfrhGcg+L9W8Cc1vImG8FMSDrXMjTSr3KEfjXVjCqpqgFGCP/gtt9a4B6UGtFytL3zsEMO0
2tquDLeAj+bB5jooHKi6h/CTcoVo6OEWqF2O+TxF7B3X1a84rvoXtddSTLIOAZUoP1BUMXNGabcf
gD8XteVAO+15hN23CEAvGhOtywXqxexZirl37KecZyLNouqcHtpOC1LQzZlFHLnppsSpTrox2f4E
+39g20vfHpip0cUVROmAMIoKuzdEkyW/mFkzeK9AIUc8eY2n2T4SOskYWrukKP0E8ldOdO0eN/9p
2hoIWUY/TsbTq39UxjKufGNBPZ76XlvHOKvn3pFyh637EEK1oBR4Tl1snET33y4iTYiKEFhr7AZ0
3xEiSlw2rXL0lDATrSmJxtJybYYpywEnnJc11ZPBwDH+SfYbe/CSemRU75O96nEhwknVwRcPlvA+
zoagOwu9geI+QrKnwJeP6lNoKQa8tzCK3Oit3XHPv8O3ZTsLexUSTS23hVeIdzm4U12U1sFtW6F7
fQ5RvwIP9VoB0Qk3gDZH5Hv/7uUpsVrKyWKCYwoIxnS6kLO1FY/2+tpz5TgWARxcnRbs9laXjGhr
0djFS4lq14R3yx4OyP2WBXvojl65sUevs5epak9juKXFo9EGI9zB9+n9dIXCbKID0qDF9eGr/YIT
aksF4yyoeGKStXSS01BmVbq8JlYTyx3EGgbCNAU/rAJt4+XrQJzsAhLS31p00El+gjPenswloytZ
XVoY6mBcbArOLy31QNFjgFI4qX7A4OJOOWDLa0ybkgPpQ+mf6SoaBaqEOUyQXw==
`pragma protect end_protected
