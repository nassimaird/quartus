��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_��~�og��B-��e�g[���$�Ԃ���#֩�&l��=�̅;bZm�;����O)G�q:w�|�w�����H�)�k`��(l�jF��?�(ݸ2ў�_��]�'gD���x���w�l��m��-C2�kB���dR�׽
I�?-ز�ZY��Pl��js���Ԣ)Ju�؍�%;�������۞�s(�d���*(��bR�I'��ht���D����X�8��=6B���gXk[�Ŏ:�M�N�d�Mc9��k��s��/XqC�A�=��Wh�t�'�x\Ds���^|G�v>W�3�=5���\x/������R��+�j��[�^tqb��S?��8�ݐ`e�%v��*8��j�W��;S��`ۓt(4���^�Zn��0�z�>��F%�:�.ބ��w�j�������0f�p]�u������h�e�����oE�ð���Iq���aL���Ӵ
K��O�sbO��0sr����q+���Hf��n��9�˶��s܅
2v�g�9xF߬DEt�5(��&�R	��nD�Kp�o����&x��6�c�춍.����dGg��/�y�h�Vv���)�a�k�[0�A�����F���b|��Ɔ�d�m�.��"��O�YE�h��x�5y�n�w�)޽���0����gt]��_h
�g�k��Z�C�� �O�%�����)O��jߒ����S��n��n��OF2���ѩ
����7�,a_�}4KXA���$�{���VZ������y�=�us�q>W�R�/}p��CR�-?zT�Jo�C_�V��6�)`�������	�=`�^�d�����9�|7����Cb>!�!!��n��x���e��h��\:����	�����.V�M/��U��B�T�
���ɳR����^���/�3��6�)�#��$4�K��A�n��#
�''!�M�}��� S0��uS�aU���LX��^�3B�?:�*�U�d��$�	�J$����҂ek7�L�:h�{A3d�*�����g!�)���B��HKpu�ĊU��'�0r'�PgB��]�94�@�0�<s��}B�"�R��@ڧ@�d�N�E)�Lޚ�����Y:yq��д�E���iO҂@�z����>�}�0���I)����J`�8��������`#Cc��h�_����E�KԹ�D*�ƽT-�jnM����Z��W�Q-0C(�:}�o9�s�7mCE����sv9�c�f�D�4��魺��"