��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_A?N��Y�jo���e�YI��#~B�t��@E����2u�@��G^��8�=�Q�Ps�t�N����ꈱX^�1��Fȑt��X���ސ�t\J���6����9*���$�L[P��#L�pfR������N�Gm�IGlr�FUx��盆(0�ܥ�!٨Im]�>��r�J������<{��	,�Y x{��a���T���9P7	����p��(p>��7YN����aD��Z�<�ѭu�W�B#�X�fn�ٿ��f����x�ڦ9B��B߳&B�24��f�����˹'qF�R��nE'��r=	���Tf0��6,p���g&O>Z���^y0�S.��RF����v�����CG<����G}J����y�'b���Q�;�K����ɘ>��سP�̫�Tہ����`J�� ]u�"��Mҧ��Mx�(�Hw�g��qV��8E!/=Н�-�9�E"M�3�n�o�b���� �P�Lc�! n���v�c�>��n�a}���D���(��G���'D�i����}�U��3��;K������Q�&�3����aLxmEQT義46��W������N`�hl���\ �ew!�L1���a���g�]��)<�cG��Ħaý��)�t2��a��_��t�D.���Q6�����̕&H#F�^�(��:��i*F�Y�n�����?������c�E�	Կ\�cb��z:��W,L8����o~��@�F��r�iAds�U	��̺���<�ʹ�m3V3=TH��n��@W	��#���B-�8C�S��nU�H���|����=�,t7s�c�f�4#U�^ :�)�C�+�2�(��a,��:Q�� ����_2�����c�2�U��zMjhHGd@f"jV��:��� �l�Rb���K�#�ƽ���"�}q�D	� ��=D���K�ߊ��3�j�����Z���:�I/s���e@i 5�0��}���Or�Z*���u待%��ia|?E�9?7���v����ƺ�A=uC�����`� 7�n��	��U$!	<D��:�vG�,..����K�.�2[o+����x�͞][�SNb?6��b��R'���w[7*����oh$���V�{��\o�'�A����em�J�ݰ�t���x��,�ͬp��D8�����Y�AP�ߋңi�e=���[�:��*gJ�
Gz�<MT_D�¬hb�qvf�q�n� ���B�ڨ�z��Gij������ޜ���t���9m1I<�Q�$@}����4+re|>��\������?�^9�b�)��Q�i�حo��y�%���UQ�H�����$��᝵B[m��Ds|�a�m�E������D/���9#�&p��4�}�&q�2�pD�b" -~�gԊ@En��H��_�52zZ���ݥ.r�	R�*���%�b����	�YKh�&���[�\(�D��s"^G[r�
l�h_�C�BXz�ɰ�f�M^���4h�\|�%J�m!�|��A�
�b�ԉ��wa{̥M/�-�J>���M�%�������!hq�йqp��_�K�h E-eg��:��h$A��俦W��9�v��M��>	?Kو��
�n�3!���0����+�����+��k�E$t��~	�3�}�衱�6��?Qrz�)Vz�ZP�|������X��*���=�9
��l�tm���=Hd�v�J�-���wѮ�#?�qyo�!�T������3��	�\B�Q�X��C ����i���^�g�"��qA�;��6� X���v�1չ����A��婺XP��
Lx����灰��#����[�'D�_���4 �wt����l�����FP���r7Ԏ�zgU�pl#�@�s�L���iǐ ��[l�Q�9�=d�1�t�xsK�TC�}��D�6�Sy�4����"��䝫�@�$ߦ��UmZlR�Y)BUEC"!�8x/�y�D��}08�Va�����=�:/���pm�c�F��KLfR�T-��J��SJ�UEl����ܠ�e�[$)�+Z*nqH���ѥ�v��X�l��q7a��"��D�0�hit��N�͎��Tx�U�F�6D�W���y1�	�S�	C5*�*T�J#/�35,&і��[̒�2��}}�L/(P����m2��d���>e�ݴ)�Dr���۳-��K��q�$L���3������\��5;�4��C?�D2�8V�N�ڂ��Y3֛��#M5H� �d�/��]�F�-��E֍׎s`�8��E\(�o0�u���l�M�b�[���f�>ڶT��PA�!���]n�;�MyԴ����Y���8�L`�/ߦ����̨6�
�K�u�V\�:�nH��);d���u�}�����U\JU�#��@#r>�`v�Ek6�[c8��w�spp>D,=o ��M�YO�2`�_��΁�0��8�T~�F��7�9̈́����o}��l�GD��Fsdx}��Q��A��We`ƈ�����=!8p�>,^��E�I*��w ��
b��o⫓�$X�	��TS�*�ݓ�t=�1|x��	K�k�Ύ��5�G�:ayfђq��rGg�
��g�W��lcC�]w������k�p��b������-o?��ã�tq�2G�ީ�i����S�[z��'�A����i��gEŃ�����$ Y8.���N�,�(�ڐ,5B^���`ͤvd�ر0q�A`�O�Rm��ω�uZU�i�"�TOD<�����C�I�}�ԩ����� "�|�k��i/�:A�LQ� mw�2���S6�r,�X���P���M�#�d���>��vSW(VK��������?8�aPx���aɟ��fiK]�"��sm�`Ј�H�O{�88#zh���r��41���S�	|Nb%����Âhճ���RH��A#vgC������^�d����J��ܝ�D1o�ϗ1��ؕ7�LAe6���\��]�ϣ�v�t�)M�_zJ�HV�oy1���Z���ީ/.sU/�����������_�ѐ,� xϏܿ��Q�Cҭll�[�&-�6#N�(���u&s�w��"��;ԾV�k2