`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VthMJssoSE/miwKCPh2AH+4hT2LIO8TOLsB0A957FpbwTRzUq0Nfeu6L297SKBUC
Qk3ZfwDJJWavV8w1IfjoZ/CpX/fsz459WKgz6WWaiG1643tcW/ft2zAF1znm4ma9
m2IO5LlyPsB6/sXXlN2UROhV13EIc0ItyU4yeVXayhM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21152)
5A3f/cvdfTafKz4g969qXQdcDCaKJ0niO+lm/uavu+Eklj9GZ9biQ9kvGE7iQIXP
luq0b8OwyrjkJvVO2nZIg0u57oVahzZoCj+vfm+99nSRyETyoTLeWsxV6icPD7Le
7AwXC62c9/qQkWwLaPH4OeMrTYFNWdY0ZBUrPXqran0cfuLfEmV6mLuITP530SPu
tLAJ6iuCVZUMv9MbxaV27mw9cfOr2jmXS7JZqLT6+oWTl5vj8MoPhG5i9JkCQPMM
njSNa6dJ7HR6xNTO+W+wxhxInxqZAIsu2gLzjRGdAcY57fwb2/8XbnCawcYuENbO
TRUxWibJOLA781RorM9GvhJxcE8pzkRd3PRhOZWUG86rB84sJsriV/DPMkeOU/nL
rz+pHkv2AJhgO0AvEA9RjfNDTry1hJgdjPKB0/VU8nOtCWrKBOrV7B/ebN2iF/PO
Z+UMkd5XMAWbk9SVDB4v+X+xLOCd8ahw+J2a6eCVSoTjzm46v5TxiK6p3ZiNoROi
RSFdb5EniCsWY9grNXi/AMwz5244EkiwiIxXGFwESI+ogITTuKJMU/UP6771C8Cv
f0ie8QX/8D/4AXtXkHWTOObETsm0vgz3Lue+p0tHR6oiaqeavYK+/0DkAn5P5JOz
gJoBjbDuhinFuaaBmHW7zujVn2JN5lvbpBTAXRyYp3EwysR5QJ3ZRTFA93RIK95j
C+/kETStlbmHQDBq40N52XiWJBCTEaoqP+amtTVyPZ40XjySrHBsY2iG/T/BoTfJ
q/38HX86WOyQRjcfUvJyRCWarDabMCjfNGyWXH7Un/mL8ciFQX3U8YXDxAnWTCUP
4b0TXHvc79AMkojjWkYO3XH9OWdkh37Wp8AD5qZSVjl3U3SNEwERIK+EQft9xf2n
M1yLnCxCw9qERkIaUAdjoet1l8NTjZ4FKzaRB0CDx3Q5k9A6MASP1T7BgITNO6r9
tJ2nEfjtmeON1QYJP7rHJCEm9LdixJmi1aaiMe5hPihXzDMhBt3oZfMybNVlJN7d
qHJNb8of68BAz/SDdV14on9DNdBIULLIPFxIJ0RxF8GqMc9FszG7o+YrznEbdNOh
1mSJZnBNXHdNTgS5j4FxlVBJjX2E21Or+2MWDXhPFs+DItDDHszvCAghv1DEaWIQ
UCcV7aTf5LwaAh+SKwi2gI60XoW7/3Ek8xVso1gK5HqVgJLUMaOwL1627pCkIMpd
xSauFsvQEalMafxYl2D+INZg7n4UotuNTNDB6OWc+oRsva9oOwBFUAwPZ91ZFWMS
AYoV222/vo1FDlk2co6ggUDo8Wowxs4juDeBu+BaWVB/qnjQq4o+fitcYqaAVxJK
JMl1lGAt6UzQxKyxNeMm655ILx3DZu0dmeBD7GJMQ1XTegNe1ERIBgQMmCvl3pZ4
mBHWqbNdZVpQNRTFMW2rkmE+SreGqa0T3cfEn4ke+PuXEBbBlPCg7uneGHhAh/QI
gt+bmyoNXHZ5x6KUmgTh19vpVGUFNZEM5rgVmv1iczkWVgDUBn3Rpc7B8HDCptO3
Z4OCJvQ+tljqJTVM+StGkXAmQj6YRdeQovNsY+5wepKCN65FN9b22eT56OdnwmpZ
B5+zk8BJOYU3oZf1tAFrJ7WtSFrmF/rHXZAqz9ctRK95N2wDJP0cq/TEaO301L+r
eksVWGMy6YtJnd51hSVAYWGk7GJf8uu/UZsRLk3+bg9hNUevquGacEdwrFmzc4hx
ttfcF4Ft3uKki4LYIsyJWLyUHg3jbgTJOlbYXISLruEd6Kd0Ntf0GAq4xx9ppqKn
KCyj635n77Bi11iZVPdxcGiurEL9D37SBCgeSdOHC2lfqR1zlQBfTgNzlqUjD8t6
i7W7shleUUHCPlljFPMjgxIM4CHlGxY+bArFcFjkdGS4Q436ECAlphPzMU4xmAVX
q4GF3Fgl8cfSjiwSwRc67KmfC/ecFNaQTPphO0kzd/4UEoj1Sye7n1+rjfhLH1SY
x/AY+TAZTQ1aPgRtii/td9IBESsZluMGn+OuX7rnYyDnzl4OafDtUHF8ir6AW1db
yQXJF8cnrE31eXohzczq/ODELcAgsdzwPGsJJ1n2AEincaUWISnpvu3tYLsnB3Gc
13rH1Y1TOdsTW7loOL0JJUlKC3qTB4Nm5+ykNSFFthlk7HrHBLK4XY68Bhz1kncZ
82w/5I2lex6Pyq+JPFvS0dHfQ8/c9XcyB8x7uZOwq5a86YXuM5hSaugNx7y25jKv
DSv8OpPoUB5d+7HnTPiqCppYYGr+FVUbGXa6w/4VsbZUJfNHPfxN5tAth+6PxDPD
Z/htzOl7baXNp9G6C9vZevEjlN5U+b7hlvy1NVW8Mr1hIBYdHKRFyJpw7f3Mzslu
sNLkyGdb3mlViBtxFDbHiWGJBeAS2acrZjvjCmjCe2uGWoJ7nJ7P2DMop0DLGDB/
l/2dGpr7koJ793N1Okap0Y/QdkfjI+DiGPWhhlq27XnHiOA06rD78yXKuEUApN2f
RPJq0C6v3699hEJu/mX/C7ER4bXhLW9y7F2Mgtulez0PPun0xH7dq4JYa+qbcvZ5
/Psxwu2rlua+xCPLz0rjpbQclGnCgpWvQaOGtRJHb8+m67OXLrlIBjA2vyFsMny7
Kv4QooalPP7gBssFBo5KfFPVuenEI1Ct0fZiPmxAv38+8ioaTQ8PibpiqHLI7Y5v
pjxoFZqdUnuRckCEbmDPQotrMBIfLyMfjb7MMFb+JMXEXHR4kKSlnYGZpcMeVboU
UljQ7mp9YMmSTQMeaH7lpzvl9juqiTCCfq1Hb1bgUVj/jjUX98WUPyDtcKWMd9Ee
dHQ9fSGFaqBPjqefhOU0ETidNxI50XT6yncDdupH6pEDKLgrPgjwy5IGk0hTlxkN
1aqsRCH4pK29ETd6K8XPAz7LVpoUV1zZx3nUsy/wJScjaziOjt2xRtXY8t98rcBX
1Yjw2eqRNoN2+hFcyn0G5cHTEgsILkSb1ZtqeIyD+yUQp59Rmf7xfIIXXh82n6o/
EYLecPZakJKHpN2aTGSurpL2cJgoot6YKOvmB0OGEbHMuINA22wKBV7pEmTjvNck
aBNck3q1Ddi5D9S+MjKmchhavReqFOCYtSPewL+NUKroyWvSZY2q9UnVLCHvmuCD
DDzGmvupCdLisbt+NBy/vfr2mH+bFKxjZgciyh7I+CSh4lPraep25oekNrGEjJmQ
NtByBYkshWPUJ4fa77M7HOcSdpYhuNHYVz1oRe1jf8/RtqxUVqrmGQ39UthAPSFQ
egvLGvw7sg/9AtHl5YjrfnCGakjfIkzKWmRUR71rkbaICa1gT5PIu4ScMkFgG+kQ
eNvgu3UVpvpf8C06H6L5jFYqehmil3Udxru83Sq5aGW1cKopdUM16/G6q57vjpuu
FoPO1zLLwUXRNGxSr9UcLBZ5yhhEoCFTas6CCZTiFBlrlliC1qBWQWorouU1idTC
wC3o/waEHQ+PSX/uJotKsBnYG88L/FSaQdGitgUZiBndJLM3fDVMXdi5Lnxwusbz
VmLWi9ipu0YfJ5H6FWL0hMIXaEQWgmOOaoqaEiRJmCkOPTN74loPLpTWc0b3LaxM
iyuBFQVq2WTFiMfZaigKndhfdg7Ota5m3LogRBJVSYKE52A+rFzMydnJIhXOIlXz
CAUOsrS6QqP0pOUSmymqPfzvUySgmgNXAdcU/s1MSHSFO7X9SGrc09dLY3U2Do6r
pfq5RgQUgi7k/62bnPKBf2JnmT09vXPvOLy1wqwk2MVoiSMSVvP3e92XF+6cQHQY
UKZ0f535diBt4C8WnZVZansx7d3vhoLF+nfD14T0D083+eIF3yz7pULSIDyfvKtE
QbF8g9eowupcAcqaTlauI1Cz2OyxtciZFbSLdfFpejgFNGJP54GhdLxDzfebvddj
4Dyw3760iSXKnCHOzUw7vJgVg2MIodqo1CGzR1yAfFYUYowjHD+tTC7PKZ/1UKnh
U4WJZCL/ibD8gHid3qsaF2TT/13l7wOCFjQJyKgPfaw7eAHdsiaAfAB1P7MjltXF
FD7OdxJ7QzKU2KXTi6E5MVFiCiOnsiFB0HsW2Bq4Jx3vYt5MaPEE1ZdoPCZzFh6m
3hpy7dxV105FGasHLYK0JuZttGMQd7eXhDY2XiMMv86YmlTLbJZB8OhT7jH+eL5v
XcvupQsMlzZhY5izxX2+Ug8uh9Ikm2EQGKkXmZzDe8PyDoB9mAJ2mKeCiT2lXShd
LPxhl1wqzw47WdUb1THLP2hKFB/QBhShYt/8NH0w/tfVrMyeM40f6jg77UJJJ3MZ
Wd5LLNmF7YCjlirK/livcXf1dTL1sZFY8dKDJoMsnNvagWUvVSMUKzpMWIDUHkAd
yh4hiYGC+C5DgyqBzIRrXLnyTkF2/ZFayNb01+MtBD20Wd/KqIY4TUU68sJWRf67
SjIMVUz9om2u/R3VthRD9/q0D0E6IgBDK8iVyd/k4RJCO6t6Y+v3lFgQyW3M8Oyz
Rk5YEcoesHL+tHExj2bOOI81h/1jRccS/95fQwbd2+dr/pt7dXhEAt1MG1bAZyWA
qUu0wA0J+fZyidw36nWgIugWb/wa0Apk1EZwxgfa9WtBlylF7A5ujEFJJwZ3e1ek
FplSR8wZPqwgC+5r6CY4HNaUrYRETfXoAy0t5Un1g7lRBWQClgeDdiF0Y3BowPtY
FAJ3kZCHQoUisdAJF0ONQNvruvfTuHKmBUA2b1T5LJ66sYgOKguhfjpZBVD9sKrY
hck/CpJxcbmIGDSB1+ILv1FTGZAKjMOlRxUFj0RxjsP3SMl1VvRj1jSJh81qxyU8
9dCqCuRS60bg1NXUdKaHlVQXPVavR2b77waWxNmmzKz9olLHfW7vL0gk92SWw74n
LcAGMfaFuuWqB8GSwofpgNxdb8Ca1uyBzh/KZBgmwl0fsb6T+HjAPbeAFAHMji1l
sY+Cu2STfwhbqwKteQfQgyZU6JjjZaXVk0m81uoORqIqfefPyaKvLxIiz3f2ynrm
UPSutTh5KrXkev1PfvVQOTZ8556EccunXRiqeacMBlg06n5wslzd+iwTUn2+C0qA
yzg8BgHBeqQRkNFDctYQfaQD1bJPjBlkj8Vpyq5IoL4oWph7bt1ss42hKAHszZK1
UL8t3JTDOh4j2085yX/HWQHNfQ5M5DKFDPOxZkJ4ycul1t6wR3koLLsu214qexGu
eJAxb5h26YW/z9Gv0EE3aZ/lBSfv1Hh+PSkjbjnyNGfirTI8b3PDaaB06C+n6jXC
0DKga53esOJknZ3nonbQoN3wGCRecqBL80Hg2X0ozXBqEK3I9+1dNVUofng4hFUC
f7+mZj2jEC5N8AfBOnXfGgv2vBNsJ091xeVaqpHW2Eq/NAai+V6dBWl94TJBEsWe
NloaPn2NzshaZORSdTTk+7ClRdPEe2SZbNlYzAT2HnqBLaWQy0VyX7eQ5vy6P+E7
3bolpiUtE43kIekLQynq0+KMUS1ZtNa87Dex8rkeT2lA+PuULv7pRg8HpHCegC+E
mTEPSqBs6h0gdH3UDggTD50wwTDTpnV7yBsMDDvRXqiG5Cb/dLXcugYqsiEfPXLO
C25cvL/Oy/ZGgefNA+rI8S0I2aOt4H9lWttx0GPUy26RQaqyAoCLOjzkCup0e95W
+UJYSq8lotKnRsHuiSjvFlLWPS97nw7IuCugL7kwtcvWWQ3IkzfmZ1t/jeB4qocv
FW3sckQiJ7zHDkojmwJJfsNCIzd2HcSaiHZRZzRUzMHZ2e9W3gFDF21Rqd0hyLkZ
Qa1dMhb6yV4qPe29kGeczyCTYvdOJm0WERXps/uvep0Un+VydJ9iUZVOK8pwMmub
EplmSV6nibHKj/7be1iKur0rvtaVA/WfCKKgy71Rqbf6Jdhp5HGpojiWz7Q31z0v
g+vbnlk0CnRE4UqX3cHg+c/Xvvh0wti5I/sLgHBbQPssNbmT+PhzDvzmB5Jt0/Zk
Tq87hC7gsRMgjceqCye8ZG62+ReHwMYt6UATtbWksAjJ+SNMY5G7RUNrW/mDPQHP
RYhcaUntC4TI1XS4jCcpTg+xmLZcpea6PKXUNCpFLs5Ly96q8WeStyUXFUuZZ4jW
Tk2p7knpYoCsilJKBq88T4bx3hXlsdyeDvyzS08lz5ZRSOKTzWWbYzbpRVmWeVMC
tqAiAUhMfThUdj+/PUu519IRdR5/+GaUkK+csJRLxkMe7ZlJqNmfGfcTwPHKinb+
dCY7R3DzsQeWG2u4Pj8xdOKZ36bJClHRbl5df004dAzuU7XkvYDrYjCz8WY1Smsw
sNDj/I4FchAvOZeAFrSm3VV1+EQxm9PGi3pZ2DhspObGFtbE6voGFWariZ6xuaJ4
7M9tqcPkR6T39BclHTRgq4YlsTeFptdS5+QGW5uJhgXVxtW+S2iq+mKIOXh2KtM5
2LcE9G+eLCAkz4xxrHnDepyv9Zc2OiRn1FZm0xJcigcBFxL8v1sl8d8AjZr1Zyzb
5rS3lznX4qaEi/ak0l8FH4X4+KbGiBDB/2/mQgIw49xnLR9EP/QkOAfzRY7hCQRU
LZijK+NWw9hA8826SUBzam980X7svxot9V1Mf6+UpDZj4UG/vk/Zdm+iX3hvTdQ/
aGnm3j5JSyAEuMGYfNil8RFddLRRT3DoCswSFW4zgSoUYRGoCmkplJhaJ2+5Xbre
rnIxKJlTabDI8j2e4JI/MvBHFyppNGBXq5TJjIpyaoP2Ne3eKiDNXD+Nq9LrSmpl
RNvZCHJQuFhSygJsn7zDqriAqPQrI+c7989Hkm7cmKvwvKgpWvmq7oHHA4Bmz7ym
HbECa4gEcKtKbd6OhsgwBFBEwsd14Mcl4K+cOI0WN+CbpGaLb9/jKF5hWnvDIO1J
OFnT+pVCfrXliyfll3UOIy2TmRuz8UXKjN1SGofomL8Y9WMD6ow4ny89EBQoudGB
Oqg04Igliv0brM8PUxilt4Ewo1mgSElK+J/KdS2cywhB++UsuQuQvnp94g4kVFPN
RwIfunezcuAEn2vWWPh2hmIYeZpw1O5+f+ZpOlP5VZgCiNLuQ1QLuwHZK62noWxI
nSVpiSeWXwb5GPx9TTMdyymf90EaPkvNBXk+oELP+297VMtHgwNEQXpk6pOcNPuJ
kngXMsidJKJKeZaAgfIC6fSdJhTq4qNek9gGrBiQvKlx8/O5pReluvprWfEsUeNZ
SrMIM3qyLKGjcFUyl5xS7DC+Nnm3POuYJ+a1tDKr5att8SdGZeVZlSpI28zU4tLe
CffsytEtaro7ej6hBamD/QmexPf5YZ2VPpfdf1rfd12gC7AX2lQX0TEgzLBTujb1
ohPZWX4hnLJccLlc11jzxbs4r/xyhgbPzdIIhwccSNCqqtGlBxQLHfw5D95EP2wF
xg13owIRFbSSXFVNkauiN/2Hl1l0mJwhnwJPeDYY7Ysm1zGxbgOzwbCtVCka86jB
C/4HeTohbti8o/CfOBWqO6KJCcN44Ny8S4WEqOIaR/FvTkzDaGY1gElzRnfFYDSz
V+mYWBehEAnOBAzcfY1eikViVR6l+SZVRP9JS5DGmDCB7snhT85b54kr8E8rN9PJ
W9r9er2o1gLuyjy2Aw8s6/mB4Ht5SBhmLEiiAs5R57qYcypNyr/5utb6t4Fci1dH
uazGacEM03+lu8xBLmoyBWl7qpXVg63uzUEwLBWgtHdYMHd94I81GIKJMXXZ8PFN
pD8dlj3s2BtCVGMEuotS82F6E9hFzSEQLqFAcMDpB8DkwxvvT7WKzrocBu4sc9Jg
Rp+zXLxSHlIHIi4nabui2dEVgArGzw4zabZgHHYAdpe/87DP59HHS2cAoQ2++q9v
TS6ncGnK5z0c7pk74ldbtaLA0PNuMM2qXwBRqiCTgrmfOwuyzl3U8lCRGmDRaERr
9Dw9/tnq3vAHfFmavhcjyWeyHVzSETO/cYPPtRIQUhSxicl8rAYMNy/K3Gs5wWMC
sw4cNY4PHS3e352hPeQUJPd7L4SBrN09DyJ/JiBehrLk0aecnBsPxoBa6hNwtXhp
6r7xXo1ByBX2aMb9XNWA5rJgsS5T1LtAoiUjLBlmzWG80UykHaCxfC+RIUdEqxhx
X2fb/bsuuuIkcfZDyH/kGd1Ai1MVuG8/4sJEEsCMoKePJbUtqplTcbYzfv3Sc9MH
3ptpp7CjHWPSxyuEgYtYJ/KMG2vBBVIhKIm8WE+ySWT1VAGuYz0qsbaG2kmH8DHy
8y2SkeHApC77r9SnSfGHd+JaP5C0hwXBc5Ho1/iWhbozrkVLZVXYAQW4Iz0CxdQv
/pJ1YKsQMAxWa7o2f54YK2Bo8PZO15D11dQUgJAnqfK93x3gPgs+XOJvZpKl/Uq+
dvurzJ63Jk2tnlC4rQwQpo6R5dSRLbRBHS8QuPGCgNSysytWJe0S4RmqFBah0zL3
PlKzltbqQRT1NZAfLktf3JNF2lN3j6mA2ZHxKzgM3znK9gzgrjsr9zxK/vqHuOX+
WvQXHw6q7MKbjR+V7lhmGPVfck42HoWKl6kw2DzB4duqGC9z11nytIhyryfXJNkr
iHLRE+T52kn84OjcwCUg1+t9s4lf22W48T5EhJ8mtks2+kYH+aXQMRsy6P6eSSsO
STO+ESHj6PvPgDzrhAdT8mXbBWyWacuCpHRzoUT5qlPWw8ZUj1L8N7Zk2Diu28Ys
T4PUJOsXvm2KPCtUlEKJ9Z9oGxOuvkKaB1BeY120wrNgDxEEhfm0yrZu3lBKL9uS
VEbK1tBz645ECF4HT8omoSQGHamHC127U4MQ3Xe7j2frI7Fnzu2nU7T4eLtFuALL
Pp9hSczefpbbhuhY+ZtoHVOyJP3b/AVr6+yrlumfTimgKGNjD2uQ47xzzCFBBME2
cGIShpMbhChu/y2HnrT20hONiDxmZflYDQDgBxg0ByZNYudFEA4Mu/KkIAyXCjX2
JpBIpllpjNqHl2iCcD06IpyFErFCIEFgv9+1pMyLM0ML/TSOG6wvnaT/9XwrQBJQ
CorgVSnUJc4ZEal6kY3POySqseAEySQDR145J3hrpoU0Gw8YOtC3/mrWN0Dqk4KD
j2ckBqu5clK6cq6bYr/qaWB8KIGwjd84uyKZyXw77qvhKp3gZY0tT+c2jfcI4p1V
838qmVFaW4xfZ5vws2+/Xdf0koTquOyRyt3rdSNTFZVEbIjxgk9F0g8ymYSfY0UN
BKmhdBQ35+Jrc+jVCVoPpHs/DHryFNE6SVuCXQ//CqXh5gkaSRIvrXtTBO+UONd4
4Wua7mPzp8Ylf3vVn/P4hMfwfL6EcECmI5YD1LsC5kIkrP5F7wL5qWcKwVNIs8L2
GWFl03vbidkdauXJB/B0jBhiSd9ah1L+9L40hVl9yFPdCb03gbBIfOwjDPe0qlbg
UPuNu6dR3Kpt6ShNqsbvHVkzeoyXcO2iHxOMLevXGcs6uPbTjeUDOm8vNIor/2ig
tyfoa4hnGi7ExHgY3LWPBy8pOemnoXsTQ40jSCciAnQbh4fUM8B798qSIFfPuiIl
iRuolDWnPR4rZyaIpB6zgnlHKNX0j3hSfRgE7CKo/2VciJkFckaeBUNqYnImvHp6
CGpq0nUujyFE7B/xNGKx93tlJMG2GMAw8bgmW14HCyWEGK98p/y+rVSlrcFIu1CC
3tyAICTlfjESyVU6sg8j6XRzqi2elCMnuHUraPRylKPKLLfSKIcg81oNhjuN23mM
VcmMA4NvfdBWlxVJbuVOsrMHXxD+gJej9jx6poogo4jFI5R4Y9uqDGNCIfXu2GmF
ikMPGYgnPQjtnpD2R0TRNndDaXS0IRzsS12xc6WSDsNV9qHR87FSeKlnZWRmvOSl
XVuqeFLmPZ4XBane5bRQL48TiK2BdezrX75QbMBgMeTjbHv4e0UaSXtu43LtoDDM
1e7VNKnHAJcmPvNimCK0rE7Za/BjZEOKYP5yexIf8ZLxb91RmemMb98gtoJorb6x
zAZl8fsyu6YEz/u++olySsrklOgepsFwQbrvT5C0r7SNxmxwuVJBaOW4m3IZ4PGa
DKVJuQ0xeKreMDxn+I+DLdLPi1k1qArNxrCkO09ceC7SsxRVL2bczx1RD0btDvRF
RUxZ29I5V8u8/9fx4JBxK7WJNYP92qaExxj3BvGMkStMH4nKNiCxt9xuqVky50G4
+LUmg4C9eba8pfzQCPubKBNLJYp03nAl7gQ4O5tdU7vVQxsWsxxWHRluk0m2P4O/
GqfCixY2aU2RrrTpuNgSVjolEsrEJsIgGzD7z7CEkO3uW/gZjqEg1JR7G/+EikvV
xRiLIs+Ia8xfZrLPeWF7D4VXHeesWkGAApA5k6DLRgz9n1mWGHS387wP8JAAxfsA
+qxz+99DhfhxGrwnKkaQpDEGKMXTmqOXXNkM1H+Sz+OpP8i9NfkV5Na/ftZrp3IT
GJMApdEOo3Ihn3YvDZk9FjaQp+eNlkOTXhYOMhjrDdFMzJIuobYU+IXVU9DXtMQc
KdrwH1/FnBy/RoQ9HXE9i7LcDQoGkkc1IPoG2bx+HVD/CAyVUtq4oolMvI5znuFh
NfD1pxWoEML1UJ+KyuaAmvVNmPz/bMOH/kzo7tRl9UkIjJEEy7FLdEp4FCjvrXBG
4haZZzxd9/gObSrmS+J5WYRoGZJ75QzzT27Eyyh5xPtCpAMafWrlExQZBNk1VnP6
L4InW9Po1oO6C+O5qinun7rdzDvHldHr9xUSVfOpDmHG076qoyIijBbcgcDvLmC+
qn/oSOQFfvVl+0R1YJlDuyLfNvxdFL0E1ZMHYJz+fvXN2t4GWacxoZMO195dKuqz
/L/qcAI2ewy64ieOr2e6c5xWS7jxWzahQYMReregV+ShUdywTkveK1g38QaPD2H4
JkWh1EhOkYIo31OPnZ4RgW496CbmvYhvHQn/SaDIyX6yLGkO/q79Dxqndp+E/spa
tL9GGoe8bzR67HBMwk/tKlHVBKHx8A+sKPczbIZbPaRAztiESVFCMsIOKEAOR5V0
prkf8qgOlyvD2xIjcGGxcuQQlbPW9yk0fVBo/nDNpl8M50Jne7VIFKYu2m6GNSRa
hcEwwiGtDhak0i99PG48Sdbcj6CGeIaj7EQMud7wE8pO72JE0l7kLTtE0u5BNG0N
ctyDeVsZtDEQxx9kgph1URU1jNoGzp0qs3206FwdfyhSQn9BOrsGQrroS8Oy7YQL
TehyZsQU+IzTz585mmSPff+D1Z4aa7ZeRAIp66FHK1Ud69gGcc7EcXXL0ino1l1j
I8+Ot/wAW7ilHDp7LezbfPKOmEC0LxOG+R7dlEY2xO3oTGxIDiJuG1N8JspocK9T
GsHmcdBB/d2V7YTVnPBDAHaPZm9E1OTeCkmcicSLCkArPKmvhzrwtQDj8pcQyIDy
qQb1dyug6bths4wcX57gPrmf9ossjbExuJYIRA28IvxnrwVFxDhZccP6V3v9qwz8
ienmOIHH3UJ8C/kob5Z0GOKi4G0UMgBWp0u/IUhvKm1aOUErjbObAyJrZ6dZ8ZWj
Ts88jOPTEvGSQEVPBQpHV/olMB6nklKSO4Y3zQMUwkODTurUWCF19E27Ag9ekVjl
uSc30k2r1JBdvBNfWY+2lY4pMHcsJ49U4vOjNTdId5EcXSUhBxwhHMkryZTT8SAD
R6xFPozV+xVhoX0dDcwmEjQkfS7S8eNFR8Xc5vszMELV59geBdrPAkbXMw69puzB
a++55nHJz1ZwiuuN0FgxTgxhBxJqZEC4IrYWcIpw/lbieRyFet9NnKHb2ovSadbX
eerVUzafy2/pC5XrGI/swymoFzSVQ/jVPcYObCx0vjPDasT13yIO4pM0m3jAR7d5
Ye3JQYS2BoA4V0Vl5RI9HfaKoX/hzeRsCak7W8rtIzu6wiEH0hr/oUGYfr4J/K+J
HOHXNEiqvnrPZUMp2lJrcRjewJL9pDmyjup1NDBqYb95tAHhtyZ6SpYpAy+jQgfW
5gl770mI3UsnkJ4rN0VHJNKaGjMjN7ufCpPUMeWG76baEabXe63XgNkIrMz+8jWd
4yeKLlpPtaz3dqnqcTmKvUKmvPHk5ayhy5cDjjKIXCnzf3cY6EjTPfvEOFe5qQxH
H8qUsgmh/ObcTpznkEgstV1mEgMb5eOAALSvokf+Ws0ErAOzAiRHooamSv/i31lE
rJ9zL/rEPGY1uHDvwzhgOvyDYWCu3Mous4ykXV+e9cUou5Nnmu6p43Cb5eYHnI89
3JM93M0nvd/m335W6z2xmWT27hlyY4nnRASY2Kenz2HAux/kf8Txrwrfdvb3xSMc
EqLp33VHmLkJ4TZTNEhtkxhoTgQA7BMVizuDXtULrZ5ZhvQTwS1cmjnUddXu6iYi
n3vrVLCw2wyAUYnJ4GhLWMBWLAt6bm59cBpjhpG0wEB0cs71R/XyHojvW0q7+WYe
8SyW7mW0+M1kII0rqsBcgv2ZuWUdJE0EJF0VBOxm16qp4WBRPxTRThjo2XCjawYq
YaesJ2VT9yPZN37nWa1z/hVca6xLivDpdLdxXsK8b9SIzpyitwRXuzKc0BeJMpbu
JTvBjrjedPGIgWDPQo0VZYdfwPrUzpejxM21rQxeuPXwPkf8cjLWZ7XsXeZhI0IY
YBoq70KE7IobhbtelpmPqLk5TVjGxad42TVcbd0kDvmdttxmcxiv944ljyJDTbjJ
mDAToXl/4hRx8kS0OF/BBcQc05oNoih/kVZoVtZ+btvjaXCDQm8aie47Lf5+GDHO
DXcTHAGUxQTc1yLa/MSG5dO37g4s2hyeqZe4y4Hd/EBcg22yI9EgVxwN3lM/IloW
5ULumPaDMAE0axHfvrBgN4LHVnlvPjOOV/DNJDrESdW7Muje2/DsJZ0R84CKrQ6+
rrMeq7mM3k1A1hz98aOdQFa0mgAoK50SCGutrfpHXbydOQ028ynkkJ4+4iw9eDJq
yhyY7K1D5lU3BZJTSrkQ1gq92jXaBA6PLblak3m4PpiiLw4kX5NW9l2gC4Lcd/Hk
pxJVDNQJhthpckrMVeGBRySbaPwp2GBMwZWHBoqfXjJdQ/13dKc1r5TW7b9RXQIh
9CEh9POeej488Qs+tvYAutCRUNYsdZ1/jABh0Z2rsbL7VYfqkH9qWASTbRXdd+bY
IyeXRRGxATt6m4JW+mwOOb5K7WoJsixA5DqkPoZME2S/KaKmXKel5/IiD8j1YzP+
+uCnwCjufbd7KpP2sIp+Ab0dfe1XQBFqzCViGsbDnfcd5JUB6wCHKDWlud3cc+de
iYqqJSBZXS5w25//UBfePqrKQqIub/RdKrekhkKe8VnSdwqg9ZJ5Stpcg5zJs0eC
4syhRRLpYYask4AITnzTq51SCK8WSqG/bCSH8Ui+hcqlf2L+pdzuhNv6zmN4ornF
E1eRziITs9W2XkSgGf/Ha+1ScRH7FDal7MeIguE3RHG6YuEjv3jmqGZIicEDpQ1B
WUNSJUmXK3aijHMxlCW34uZNzYSsSIvxfoe+eCm8xhRknwaikX5BbLnITCFVYTX5
nAg/DGzIYs8lB4ilZn4BzbifTyqZbFlMKFZJVqp/FJVLwSnulApDt4NHVE9uH5os
/qSqmba8I7a+v7Twg3p8/VS3eu6xKVCae7XNQlPqoI13eFoUaiP7KEckxPUfuLFT
PgAPIARUeFaygdpq0WLwtIFx5YEBSCzvy06cHaAEi/ZcEw2ljI9MjmtMgMEA9fIz
V2uttCuKFoZul3IcWhdTiu1DXBlHQClXZCO8O6Sbdo+ugzHJtUUnKMfC9mAv/5Pw
C5PahsTDrrd0AzBHP9tlJsw8+EqNXccuIx6rSe9CCcQ0m5MQ/Z2//m1LzmhndwTb
sSDhxFDp7q7Kgp4apmQR+5pWAKANIyejycvl6+4hgsrdNSMq8k1morARAKEjLRzU
qtRBFn3ZyUiaA6o56LDbq4WlFc2fFxKp73pZOYoToC5hC1a16serB4CSiOmMpt7t
TMISai0lEHSwJLk0gAD8yUo4u8+lMld8+uKIr1K/fiwzZgZM+IF/1HNzVBNY+nMI
FwhAx6aNe03QyYLXtMF9dfOB0jVmXX8RT6cAwXLvQEDvjxRKHdE9SAlKGLBLWFQ0
lI4ROiDhcxdaCsFQbNmQu8wTSKQnojHhOBK4vnAIccMK9ip19oi99QTgrG9pqJAM
t+W5S9RooX3lWsIIawgh5ulE5PwpVEb0/hH0VoA0f2KG9ZJERAQvJYgQ1ki50I5E
y2DO3QCskqwVy02gQi/DH3D96qrZfS6JXxMX29Hvb+L7l9Fx8wrOt85h7Obn6lto
AAnGRGtVMuEdqgbSGUxdYIgd5h0LDxvanA5TOWBk3b5NeplS7TsgeULKMKjOhYtT
2FEr1Bq0NDNvLXxdumC2qxyNlY70n7rRLPdteko60UALzq0L2+JDhlqIPvnMo64A
q30iZs/CtyMcyGO+4F+q8asKwdowoY7bLi3mCjD5JNf4sCYZTRO2Td9FnSWDRsbF
To1NyeuOVyEabB5aWoKWlMmTMXbq+NHnEn89SaTQzgmldJaEgbts7T654KE/QDrE
YOKZBNYUohwhtpGsIkBz5CO09VNiHNGsTFXHvpNg6rb7tzfiLg2UhCRWNWH8/l46
JyUMw0o6ZSMPVFttr3ldzPRzkz5Un25gedrJqmIYD9dQhFxfak6NM7qE6RauTPMP
VqQkO5vwjl2Cs+p+5UbuZ6AS7upZrufr0XwNMwZoh3kBXcHKyP+cbWTwpEKM4O8R
+/yapRQTitCztfOfh/u0hWedEFcoDrdQ37cV+6n0DBqToBBU3uRTMDXn076uUzRj
SwJPf1A11mx20V5d8nFOSEMJ4K16xr3pD5LUElue/tYImqiLPrbhm97q63guxRUb
CLlfuQo1cpsdqi/BvNc1YCLeShrPT2KkUqNlB8mgfxiEDZcq7qcXTNRkKcWw0jSX
2Go42Fpdx9M9GTe+0scsxkViBRpBx7NjpA2iHwyf3YKmv1wH3xQ/jUXR3QWE/nFT
mHM02Ed4ROvBJYiqWiJ1f59yhKLTK0HznMjm7khQUakyEDlx1LhAyGW1W34LohD4
ZkKMxmGKZu8s0WeTTuZXtUKjjbQXw5/JitkXNsm4D7x7Inyv47w32dCt+UnAQc7d
lUasimLwIU20Nai5JDRzBnH3SkXsRhJxjcPj1FC5jWVfubJkfM5DIHsJx9VDZ5IY
yAblaXw3M+62ztSGgb5By2a2SQOKt/ok3HLyHRpJX72hMcZ25FSb8Ykmj4RVyL+d
4vam1lIrVm0ze2V+xJwPdPXhvAuRVVCO1ySOIxchUCv8/Aw+8Agq/+DZxTD4nTIq
Dpy4ql3SU5XdbuArIlzntBPGo+Q6gCsbBurJPvuKwhCYwIHS9ZghZ1rgEm9KUGAH
Xe+fm7vXF+QEpvU/9GipU/fMh25dMT7G58LtdbZVY2LlFjorlzAbOrEhg2gkaIGQ
qa3HPmOWEA10Yn8DOvEV7j6o4lG4lAEXdATxKMh7qjFLQhLC7ZwrodGiVcbiF78l
f/ugpdQHMmVLyMT9BEpq49R8aReWlvA2FxDdxal2QWHwfbZ6UpglNzhSc2R8OZCF
xbSxpE9F+rRREfPQIsiaIccgLXcG8QACaR01M14R4NiQYkoUDXQXHzQ/5tRp2qTK
uDvhRPt02yfdld6jPN66uMLXlkgNiqdTeZPgyGMOEaR+7Njcyk1Q4cLeVkClzDdf
wFxiO44bb13hDeamBmnoy0Y65+ixOmAf10RehylIHloCFVJH+MjhFV4BhNel5k0V
yWbt0zGN3lefWzbicXCLJXDx2HgYoKN0ftYQAet0bFx7LbKmID8IoicTHyxStNt9
5T8vCgRyEBpFhXiWGGyy+01yCN/6k9Fd+kjIa36z1iRWEon4HrpnnD0rSSnsbM4G
cfMul74qUYmD+cPNGcgrqGzQqZ7DuLOqpXM5RQT+RVXYvPHAn6lmoYh7x/3V7sGj
vE2GgQLXYqgGool/62ki5BMcb9vz3mY+YfnHy1xbxdgn1HWGTSKLR2EQvCP2/V4S
TzMPPbB5IuNIZVBqDiEfC88oJ6/O82+Ni9XGRZhmtNx21WqjagCt7yNuQoZN/l0c
ooi4GoRt+ZeyxnB6hZcSq5JACYUmMq3DcLKDdo+D7K3G4Z0LXbEx+zTkyrPXtrMq
sm88fyfkum36HNsIgYu5dWyl5GsIkwZu5aYINMafdiTj9mMywyssKtB6B0Ke5Gkt
VLX2NyfbfuewS20xMYy3cOsUmhYoYsio8jKupOu0sKHhjxCYN8wXA1880qTUDY/Z
IXLkJTB/nHT6b+CoXPjst0UvKFbneHDRcWE3u9ypwcGwFiEqSAnWJ72RSkujFY7Z
hOLTisWW57KitUY48PYhVhFlVskCeZ/ni7zhEZr1Auz6+Wn5k/R8yFbwf5/3VKrU
TSefdC4eXcJSpje7gTgm9ARxUGJQSgVYx6kJz1/USx7NIx1s4kjDnKW43yEfiwgZ
KQnMAY3jJcpvYRkZIm2YIzNSssPf09woq7ecerXVWVwa0Ue5etNEaSKi+FnySl/2
Bwt+IcuX0zX7FbfFf9EoxZAQDCLKVfEpQD1DqrhdeyQ4O90KF2KNifJRpVaqyfQE
+Bw0F8FuAd8pEHwitxEOMvV0AWNb4MRwgDEeTeRHuDT5+ac8ytOcPzOMm1ZNLEp4
1MoSUAQsomSR7Wodf0OZt3KJnZKTXMSv1nu0UpqIA2vEQOZ84ZHHCbOn3XswVk0F
h6YC4hWJB8C/MtnugBzWRnwKg1wAJf0wgwMDCl1LRi+zzswqP1trLU3+kXCkoTtT
TuBZ2n3g5YkpROK5LzvGHrzrJtAXfQDlQSy5ER40Uwc2TWQ64DpH2lEceOQbOqAQ
r9AHHncxg9mEuKUIr9v3I1V35ojhjcQGefCNnP6bFx/9CJ7Ctp6M7CXrwXV6aCX/
7iumDIzEeOuU4QVVGi3XFp/WPKSoCQ9RaW4HxcTKryRAUY1vjaSfrGnKfR8nvGVD
vGCh9W3bIixSynKzTr+70kyp/6KhEfF3kWoZiE0YZiNlEXn33TF2GK/4WcFzxNTB
go8PgrOgtsm9xrossxXjPSA3LxxydaqhwdNrvVNXJE0baag8Nr27b4waPzdUcRgd
mxTMxGsrFxNNO+gATxm93Dui4VwgDWtRMJXkePQFVehlKTiorPJtqzHePQLBRav0
WFSxDWk9tHrV8Pwaw0X2aUePwkuvqlhAjHi1VbMAxnkAPlx+5hxissqYPrn6/8w2
C7DBGsMoGEF5ThMT21USeme/CX4/VwKvL/o+bSHjIQFJQIwRvapnKE+8R8rg7spo
ZLayyYIYx5JOUEDYWuNDeZU1jeT0+iXahtys7xwMHLBpBagVx72JYz9ZKVmGKzUu
Vzmlvb4kIdIxWYeBMIsFVVOKpII0f1E19/EnbJs3jWiza8XUQtqqzr+szWTyjM+L
p2iB+UsI9lR4WQ7v7/SkYX6LM4Smiqms3qFcmNwYvYeo7xrqKXh+GJcEVh57XYTS
1VUXKZPKB7/DIVqme3Vb9JuMIREbA3A6QQz0TAgtVQgiAGIQsf8E3HlcDp/hSD/9
uIrp6vk7Jjs5/ht186F8qhRyBEiNO9T7MIjUbwNBA3kKdf90SMartLdqL69/TM8r
KqRS8TSuoreffyFN3kIOLA/OU5/xTOVOx0DtKP03tJs3pADYIB1GBdR2Ll8ZemC9
LDw1sGMavFwMTTBHKT7mnBnfAIfOSMV8lTqur3tv38KhYQlNlf9ToL8CVzIcslb+
344TwwV11Av4L+Mi+5wjnXAUWpqxI6o3xsEfnb8y+KlkUzH8tJq/rKDeWIGeG/46
mx2qSq/Ty/UcFWH1eMmCpY2HE1MiQ+DuG6cpZsfmZkw7c3v/FnWtRmcjoptbjgOK
xShtJpsrAr0JKDWMiz/pVivn7uU2ceXzCKW4+H57TwLJniUsCiBs0jLrFg5rUjvU
ONB7iVkCtZX7MQdGtUYFbT8PpD0Ea9xgNMjKwchT+fTizv8Rrtuj5GMWjexd/NeQ
AG1eZcDtxLAaTdS3v2fgvhGBTofXld4egi+T4kpXq+WKvfgxl5Q9ln24zn5+R0xY
8f2n/N+VSVLhh1cyAQU1OckyOv36fyofYf6CHIIJpCx2y2ezxWpCSeEe/XeWwIKm
+mWaRYyxQBWNvAsW/TA799L7lxzt2k021jqsArFe0YjHxg9aHJ3xSLi9kAv3UFw5
/MoWk316VF/4Kl0AjO5mSq0vhQ0yqgNaCseWXwcPy1JK2WQE5Tdl7xlGzEk/dzP1
2+A35jPdjOdaCSb3zQl3VUvcQxx17I0NrA4fvPINz/hi8SdwJ3QHihIhOpv8VZYv
OepJDF4BXbudafkObFy69jfCtOlPvKBopKdr2LNCwC9aYQSyqzz4wZrB/VgeI+/D
CJ8KjqHV9iSIPUABSt3hCQ9RI8D/k60vVutxxgvnPyD2DPTMQtDGOcAvforPzMZ7
goymPTTbxyI5XqUDI+egdIIcMrCxglrXYnj/UMyTsqOXyxBtGeiJ0/8cLZ9Yzo2x
fMJaM8URD3KtwMj/g2vFqBl3ZThY6FwL4c1z8h69c5JI+HgPJtOFeoMmjUhva1Sx
Ar/Or5HengG5T58hWfe20emVg6feX4Yab9ZO4Rhi3/SOKy9gFJDW54Cr0juVz3oS
QM4hu23z9lda6e0mLf97i/CSgNAFd2zdycLf5DTINcki9nyES5AfDmD5Nc6WX9r7
4GvEiB/2iFvGRrsBGxaOdG+8ZsCMtJ2NR+hpiE9pi6qtpm8FJJkuPCfQqGs10FD1
Zmd9zrmteFrAPsynLu8clmNWW7fEcN6zXYARAmkYb4fqc4ogeyAgkq5ukoA2vFy7
fwdxJ0h0CihOQOg0EksZYSrLNCF1E+xQ+Gpj2n/oujRBxh2mT8Q8YbL7QBkkwvGm
G3x3F8DWgTiSAGqAzyXA3iXNPQCprIjEb28Thxj7cMHl48PygHAlpGZqC6gYahYk
hO98Lv36GaxBeyQOw8Vb8i6ZPTl9Pwk3SnngJ0kw3oBGEihiPt4KXNUcakxQ8I0F
hD4XQbqQ/nbaO/51g+tyCB5/eQk2CiJb3/y3+GTu0WWO/gpzwOWiWqomnnGJ5Lb6
XwytarrpW7OabT4AHNQRAzBu4HsRiB7aKuMaU6TKwPwOHx2GMuX4QPBJzExzAzBT
tQ+og/MIPqkYy7ggNUV9+iPBbepkohlozQpkIG2yvRac7ut+IgGS+1n55zZEVaZW
HqCP0JGo90SmBY/btrtGVGo0b/ScQ4s31S5g1huPY6NXJpnY6Q8DEFC5IFBqB9Jd
gVd3YraXr6VuyhbccZUxrR/cwUP3XS/GtIXLIlc7GL0SJ4mPprtINKK9PKV7Zprj
XTMlHk8TggNxtFWv0/kp10gZEZ0WezrkQ1h8t71WsBhmsaE2IJOLOGTFYxG3u5ZN
eP5fosz5RJak4FqREMH8Iezkfy9ttMYMz9bifcnohscES5nJqGu+gdHqaV/2OCDV
V7pwK1rroD24NDr72YNPIsJMdPd5lJZHQTbfCxm6Lktz9ZnoZ83oqQw+0/cfBuGJ
+9fiuGU1fS8tlQVeioEV+A/gM9C7IBI4irHYzmzqKh/gIns2QsPB9Yse2MXLgpu/
vzLEyxPSzSV3FDXqrNR4JdByKXDubn+8kH3kWa4TO7tZM0MObUVgsUS1o9yWEE+Y
4VL919MS4uYRauoUagW+Y+es62QCkV5voS5aRlZcfY99jVRnCGLJJrVtpHwjrpMI
7ZoYJJR1iExCIYfsAxNOCGU/BtcsRn/QC8Xw+ua10kfy1OzM36JL5Zj1DEE3fwMf
U/PGq+vn/vChAbpJ3BzAA3D815jRSOL9hiRr4n/h99u04Xq+FTUdwBKEYVA5qB4A
a8DJqCRuwGZ6/lvt1oSFnMFCD0WsmNsq3JrqLnPyCq00DhKzduDRTfV0tJfCWq43
jrtTSOIAuYSa5E2x72NeClmxJYSHeRTSp07kE5j26c51mz672qg0A0wvgF/aslgn
uZa09jFJFTQZrcFWAXSGBezhe4420wXGK8X+9viRY5SSoQsDq09EFz60Xjbn6PoD
o5VtZy37ZxrquPYwlTFfIwsb4mgcdXVS9bnQCZ/edLqtqGpTY4o5XOgUiJzMv4QI
DXCpWN2fEIE+wEULrHODmuMnnzy0QrDua4ASS0IjIylvspe1QXD2kH17yX8lXGwB
C9aQw54eU7yGWVYyGkfHqk3pUFpfXxhSd63b2yo+vtoUnalWAqdMfQic7s7J4Z9P
zI77DlBUYSBEvMai5Y/nmFyKrMnjK6C20whMEAKAiJ2bx8n6BQLcJKzHVGmYmbvz
C74Z9Ny7+eCk0BvAJDsexGRbyorGnVeAnwNOsojiACoMFdd64tJ2ZFswd0tpgX4u
EsNNm7JxP5YQY/y9tFRmcYBCzuI8X5a+sAdW+MsrUW1Y1SOg+iSthmlh7T3C/+GA
eAcMstB0iKerpmzXUJ7XhlbqYsmKzIp+eecXKOMPqtUrJL88vWuLchDkLqKPUKzm
g7E69c9QavQhLM16RsoWVFooenlhPQ73Sz6WM2QoypfwYVcDDaH+EGmxQAE+MxEi
wXAmFk1Es07bR6IrTAllLej2tW6Nx1Wwq05wBasnu+YQEyP3JBVe8yHfwMVUuILf
lC3mOYSyjDiuukc0IUhyfwkvg5yqyXAjLFHpBunuJCtKSdmIgbHEdyLek+TGvLcs
mwZ0x5Q4tioxJU0CipJMvI88Tjy7nXFbFpJg5CdB5m/g20ujLNLKTcKHhml+UF4x
FR7zR/7NrwmDUymWoxe5DId/N4bZeU67nMnl95OJTI0u1+EMmn96PwfiAT8H2OWq
+5U4PETMDGhzqo+d2mSttV4dsBgYCOaK2tOShHfDiISueEtRL4SXr1iY598SJE4t
FNM+xjWb8ao5HsneoLVLPcsVFpp01QDw9Ru7gEkNNnBj611u1gxI7Oyn5kuZbCZF
NWe9ByhecBn8M9iWwT2wghCEpwda5RcXRIAxURCLuEW0yLJsSggS2Yi//4si384p
6myo7GM54qKmEo4A8a7N/sEWX5ykHEMBNnNLfDQkpyZWA91VBB/n1hSLCjXNE707
WTEImi8K6wKtNzYpeHbEwq7hT893MwfAyUSODisp1ZoB8fV2lG9bNgxyt/z8Clhn
r19SDJrX2xgL+8JCsa3xjA3IA+EsCGOc5RJ6I+c7pqfBspHVk66//tBDVKwnLwu/
jXpJ+O/eOR1Syv6m9W9MPNXHpEPnY0bBLdp0nwzJzJO0nRNSrLBRLuXtZkN04SQ9
y/ZpxjwFLraugR+Sa+ISPHIruJdf7RmYkMfgnkRZK+Ux0fsxnO8IBkDPI/b3quHM
RsZ/X/9jvUdEbdV+60ArKTJgfVTwvWfSpbXtmSfqccD7ldot2X8aOCT1hoU5Hv9I
ZRuwFdfZF8/Jvp7Tu7jqJZjXdTdoBdmHhhKHTLXk/3DlTJX8iVfu4yNRZwM9mAbR
Tb6oSANIAjcFlp+km3hfn88f2vPvx76ASFEI+lAsSkg8AZ5mFW3gmzBqrQBZ8O/H
FONN3nFIdgh98sEUHFsL+VhK61YowTWc1UnVyc7Bl47grM4olqkiyOpDGiA9bxmu
MJDPbQxrf0msyvUunSNUVPb3mBAyif4zf1Xb1BchiGP5MhSs0488bDaOZtpNB/Eo
Rc+kRhbxNHLphwJ2PUCViNAuFhOA9SuklZFNUm5AbJ1xZl5H01e7VlCVqa1zsqoR
Jp6JPN5ZlEh3Y1L49Y6vIZOzxjYyt/4y/F23yGU+NKrA9d5YquI2Vk1w0e4pvz8p
qvxmz3hQ2PLtxqZZx/uPi1JGKEjlJGd8Rwh5Tyhmh3oRaKUXiN5/Scyd4llOAXnf
J5eu5hKitTNe8ehUr1ES4gCUjSZOdYr/FV98ot3rRuEr/tcYFQW8ehkHuAQ6QZhA
zUpooKSP+LnVdJWD9n5sNhfAZGQystaj7YEDhi++1HRxBgKqjuqsmrdhfzT9M34g
w5/G/ZAJPBQqCB++zTd0THDp/I6MinHY/CqeqaVfwsm3E5tMoT0f1hjGo5bC7oen
2nGk3X+x7RsJZk4gPZB9iAdAFogQeH7Er+tSO36Wm4Utt2Lvk23s6DETEG2/4nj6
qhu5SsNPOtfyaqqGJ9eE7x5zf1IjZufFdeyqdPx8ITf+uIchUyPgWAWl4AfLQua8
woCXyrTY1tRF6QT5wBqrFcBP7NatojPvPFpkHLc80eM9dKgqO9eoPUOZIrBdgJ0B
q2cYzqXzvTTnacFSYqU70Y6qeSngDP72IMY7SW6VQtsTbOmSnQWWySPDyfpksC6Q
wBBkHfU1wNnQWek0mI3dI8EsvFpUC2OVudFkjFR+kEFxItJ+f/49VjdX3nnIYk0X
OPYR1LJ0B8rtTY1wpIZkKCk7cCpH8BiVJCjGsbnH6M/+xtYlclrX/WkJA4xQGqDl
ePpc5cX8mFsJ4g7hiZcbJUtT0SOW0ZZlGzx584tnFLDdDq0MiUKz8WEy679xkuV1
ZlX2SrM7mVW6wVTbPgu31c/evo7H+YHNt4ELhzg3VW74p5/T5FRpDMIvwuQRXd8K
gBaXm3iI2ki8lKMOd72bTxsDkKCJRP+m5Psbs/Z0vgMu/ig5mAYefg7IIEgPXIxP
2W7q5mdQugXpVlwNgGxDiAtPhf02dOUiAAflzGWXUysEQN7y9piYSMnqYLin4dg3
vPEZkxqQYrvPIo/e5rAHPDTL2WB1Ng2AD1agBMHjRuCk4rfAPKZnNPgkw6qnEkBc
IxGAnRzg2oEoNcZHiZo+0PK5brjiNkp5UZevxALDKva4LjO17tu2eDZXO/HGWkAx
Oc7Dnz289Dk5cl91nSUa2DrnwrcxR3pH468HVSqa0AVKwBUmhYZe9VB5f3ZJwUnu
990mUkU7hgs8MmbW4uATP/kIUKIDGU+HNp+CLimO1j1Aeb2AkTt/Ku+r4U2uqTym
lWRLxGh7ZLoQNyxE3+W/ZuV94IpRmb4TxxLuLXeOTIyupVfwgFWV8wyyB/WukP1v
d7mf/kKq4iQL288N3BGaV43cqXFHrmsXxpEv+c87zQK48wkFqtDBskfKjQFsxfhE
xUxRF0qFopqXf3KCDAzVhKZhruc6HqJjJOfaQ7pzB3d5lhp868q7JlBDSgC007Y2
2hdJlvn4wh4x1zCYMl9lug1LCt7Vz5sJmbgmDfI+ShNEfY7MJTxF3Joh0gBgUxzy
eLLpaMEXArhDjkk0qdlSviNdLm4D6s4zZjjcpU1CUoAb+R4IvPQ2UGTYaPUkxMG6
WNoyhXpyNsdbUbpBPu3twUVQzz84qE8zl+KGsfHUYfLxRZfTmb7AIvJbxoyN1Cuy
fEw7kxev4xg2ucfhvS2OosqU+Jl5tzGvr3MsI/FkNCjbzkPRQnZklrAcjw843b9e
DAJaVxQjQuzVbRyXK9rx7dOuGsIOKmegnTuhUeTwKi/3mUDfSMPXBCUbcVlvP99z
AFO9WNXQJrCTtX/2ff6ta5cQu+83EFF69feMjlrLaUrQQIiVCClLqAaDRayZqdgp
wAkHrxbv5TeMTB47cDQxFClAvkJEcNfPYbg4ls4Yc8maDsQIpGVO56QHPL1hBRot
Dn8inltE+bb2NNwZc71KQG5oAVXMrMW8S1056hyIQivINNmSt8KtsYihl9cSOz1y
HgGmaP7LlFsctTLWdD8iAHqESMyOlaHpjAeXF62ozT7RwZyfNT6u5VbCcQynTlv2
uEk25f3QBDLlIupA4jaK3Vp3CGppp8vzSIkktb2QDUNzMZNeSoJDEQGOqaYhmO8t
44S8it56YwPAAk3VMWGQyPivFxtbzzTbtzYJDllHJhvn2a50C3BODQu9O3E0fVJ6
yDGL3Cq314bBipvap7AHtQEQEO62xyMGkHpbBah8210/y04zGX0GeTvh4EnVzBZi
54gaj6n6PbA8oN5h51vAtMttL3Vpo+IgRzifNBGRhzE0BODzctJODVkRt8vuIfLP
zr35fUMKYUZgtB52SHKxr93YU/ws66rImTnO93BNOaEtsKSZqeF7122zlReEte4X
JnVARuvH/cxweVOi1oW5sVL3ks1dsKSiGF9F119WtLrui/w7SJDL+aO/YBkzJod6
iGhtbjc2XIAK03ozD0WcWknMYBRaoZ1/5wbbt3nf+vhTPLdAbUaUbF3lKTbE3vy3
SoYyrbmcZ729+V1CxNbBRtth6f66iMsf8kEVB82hnjDWV5iKgBoc9zXigsJFlj8s
ika1uJjM2uNKDFJKmDFU/V0YpMAcshBIngo52khHBAMjqP74fxb6CfFaUgwvo+O6
WWQpgRqEVZ7SkEsMP4ZN6DZ3BQvEwIw+rYLfmhBdKGHdcQ8xUCt98mJKen0lnwaS
1GN9kmh/Q6aWRlvfGQi3iJS+aFYLuNK/uirflnDzvkJg7uyRpUNYjE7ISZ3l/Bo3
uL6Wz86HViqPtxAKcZD+0rrrmYwDZcGz+OWTt+rCtOumA9nIuZC53piU8oQREw78
xji1eZfXy0VlZa+h1UGdmKhBTRbvrDHkt8Xx9VvTJRULjJbO8lskxPIWXJXKYYQ8
R0YE+498vAlT5tPs3rbiRoNO1VYd8U1u6DtzJizCKWTgqbl2QZR/tO3WA5JLtcrf
rskeUnjhI81MukkSIMLKzpiTM8WBdx/0Y4swvvOAvGGo10JeDWRa+tE6kBgRgIGa
kgKZvGwUThu4HBTFpvvxRVFpfkDRWlez3VNV7lHds2SoF3BNI790yy+0pYECA6lt
ABlQjZJpjUK0dClW9wwp9zk6QCecjJKscN80WuGRSWjRC8qmKEBCowWdtf424bBQ
VFXqpgkY905ok2sOeB4W2NGtN5kVhHt/rgx8LzrEyIQ5lc1wLKH0X+9NWyTBBAJt
Os2td1aUzvWA37unM1r4mNvNPPDb5xPZlutMJti1/KNWiC4BdW7fR0Xl4J5ofKUU
sSyhvS94YD9wXRXAKqma5tb/K0PB9bqfmexuFcNhj2ThqvF7R94hIDLVWcbpgle9
N7LtmrV4yzVU+LLkjsv50xTba7u/t65BE34HslVYIDdikNHRPNZkJNqcfBGwfkb9
c2Njr8vfUx6WWqoKc+OPLxJlL60Go+QElKM9QahToKoIS7sOATeNHNEOgjQvttdW
IcTrCz7/OYY4u17R8bPV6fAIEA0VEAanwkqmoE9l8FROxjme5kfN9QU/G5mEHLkV
WJgPEfEnL/8jwAxNL+sejWwqQNv4hzgue1gBzSKSExCidRQnCoGBVT7umQU7Zafk
dEPpoEiNOJAfLsMGg3wOBTeTNld+GeArl8Ioh/fZYICXRqPoNiubj571j07uhDZY
h8rMv3lOF14Y/tjDIS/N0aVRQHxZ0OKZwxwxcawPrjBeEmHI5BSs6kXq0eC89VDD
r4OQrbJkpq5rnPX7D07T+Xu0cP2pMqTTgFwwjTwrB07IhHJZOrvOLo+6sfW0F/mg
orFwLeUWbnhy3u8TiqjSkADdYQcBbIjMcuVwwG2boCFK79fdXnigDg/j+WWSH/BC
Eliad9aCVBjZ/+Pb8SpBIs0T5U+M6E89TYmWM5Ds8zSgHuD7AkqrQ9EoSOlb0q+M
ljSuQVTw3CKQkwgXt3fdXDcqR+JWgKo/6wfJc3/tRpcfTaZhLeOIf0eFSUZODEHQ
3fb/g4xb1utZjNGFJ55vXk4hjxfj1FIkmxKSjF1m7htDz7sxu/CLAtS5mN6RgS6B
BpzM1mPjqBgTQPOo7oS0ZrWh9EgOOY5EY8EgE9QwcHBqDij4X5+rxVsNVSlcbHZM
GIGM9T5dv+bllmc2X75s6kT713sUeb29YLbrcj14lReYaVZIjU5+G1UD23e5Si4r
rwddCthSIM+haB8Trs/nOSwiQ0D2FF5h/53+kjl2UtcIjd2OdD9knGB8sir1b7tX
SeJgCtRb+W6ysPXzqlBFUWA423J6Tldo7kRxMiQYwcQciKbXvS5g5Ui6aoLYOdG8
4v4XmEZ1ZvqItf64UMEO9+junF/pR6+0xo/YvAP89fFcy77ixJFgacjdDySPXiR/
0QD5cfG8AMLHYkoxZ09J7LTrnQwijpH/POHWl7jKwlHYdeytJH47+EFJiDNHQEg9
xSxyaPkC8/iPmkJP1w6+M2d2Aj0rOotVsOVDnChwHgpNFqeJwLraq1GVQSceP/nx
zOHJKXcd5uJ21m9KjBOhRSD18QMr21g9QrdmWTy4Z8qmJzI81pdk1o8ittGXnAt0
cKM1CRcVtstKY6Kh0UA9yZMgnfBlYDVcL0UP+g38sHC5KPCGvA4dtYPiK42igGOd
oRhhFOuYqWT8lZtYo8PVVnC1u655VZTPWez3x3DD5H8Hq7TBwHetl8pPM4wpGY2a
H4Dgk2uRPK5OkXE7uk2F45KysjLspspxYEUuGyb4lMuGAw7jh3v6ZwXytpKCDDNJ
e0l4uLnen6j2rILrzPQdGH1Uf+J2V9L+BPeq6E0h4yc3kvPubtE5jiSJK3EFyZ/K
p6zunT6tRZcIDDVkH37UPWoKxIvjxd/2eDQegtsaCNgcPHgAKejMk5b3Ao3/Jfo+
XjFbBYOsj8S7rQAFkBvU98NgmJ8gEiPSktSv5/Ks192CiC0/m5z1vbC93H40YIgJ
sSFm5+TkHcgQjDuhrJ/vFMAmHn6ysxqtKvv+AxOU9IjQRuKkr2rtc5eRlFZrNfbr
UQoevRoowx60K/Py8UnKUgOKp2Kd2+d08NHC5UJdV8j8HFsWbxRy2WAV+BqSYX7t
6cvtWSUHaqXdmlvAPWv1kP1WjENtSKbT6n6N5tW/Tk84Z11hY5nhDo6M/oETb7sG
rpns42qSmr1+czvGB/abzpLbO3a8uHC0RK8mXL4IflhRJM1fNadeGQ1p5dIya4Jd
7S5LBtukmJI2Q2zHTmydGWVrEhzf53QH6kaA2uRuF0dz/VwK97ns5hWKWdLWvMWQ
6QIUlw3jEgxq5HBj7Y7aZxeiYnDUfaDiZGfgMtVQuFbXnqTSvEaZBxOIdcJaX5R7
eo23tO+yI68ndtW1pQbaaRxEWM5+wsBi1RGWQckkj+kUzOhuPkh342Xu3c71mWPJ
rk29GZV1Y+f7OkzyBk5CdyCg9D509g5opR5gghGdt1dspPkIzyizz9LBVJcY1Drt
C2sOqUWLQWnxMeO3KvIwjnHwetKok57XAU20vSS/c+fO7OPUE/BOQoYeCcQsHIaW
rGC0UZfrLJ425I0KPQXUKRPVCfjH3uWAiCUuP2OFOljJmWYtISDTOqHntksOzg6m
Ri8CHLNPXRmjGRKvOoxdT5XbkeW7x3rtXWKztz1vg2E05wK96P/Ntw4y6Ag1E8Pb
Y4KXyX6aAiLogjOb8zUnwKDRnIHgmTdk+TzyADFZhs/fzEtYuu7eJ9z/3QK6QHXt
+qXfrK+I4s1wlVX3WQ/TO1r63/huemEHnjNhwID98bZjAXSW+KaIt8fo//VycLdg
KMiGZSztazYdr43HeUMX0GvxyISYD4NZi9Xl3tkhkbxbayevw9CjKJSPwgDyfMD6
kG5Y7gSYxHFpCtVk+MHqCglZcDsQRA9jwVQ6i7TR6PZb9KAWmhE2qDtMTxoeqiJo
HagyZwEh2xzQ2Xg6c/4HKiQXaic8fYhJuOWlpLT/qB6UlzAehfYIBJq5Gmio71+6
t+quC5ylkjJT58fWtm0e6T9gAnrRKeM+LZyNnspz+TwXGudRDVMkQK5KIu/w7boK
WU/6F75A9c+jT3Yhllv7JLy7xWy0GoT2OG9zfg99KqAb65bagscq32XyMqqdqj3c
7X0n5tzkFq+mbWBYW5OZX+lkeJe7UABua9WwAoQ9Fz+IKSYft5rOYhy/yfhjtKIR
uuD7ITuhBZR233fDvRRgIVjAsKLO3ufzeDqsNpiR6UFBhoSM7CVnAKr5UB6+jOnI
rV2Pz3VHvw5z8FWqlDD7d6iUl5bUrrdNo5VFxMVWZL4GOP6qlBRDkPdagt8eNI4X
NcbfcYxiFwKrHdNgCQ0MsZIoHBTTDHWXWw47u2E9IpWc0bg7UDD6tGhPcOLoCsey
vee3AovgOo0jFr8vSBAMwxWMBaznz4T9JSOiCzDFm/mF+BQJksX1p5As/rnfk37Z
uIcdP7s0PXXedaYytFRX+0rVNJitcgXZbqzX5JyDNC2nrjO8+mmlrE/lFOo+6SmO
g+ZUfd1kWDHdxqUfGNg35sT2YDm28fQuOb6w2eC1PJ+DTC4Vdmvl2EIYqCmxNLET
+V8NkKJWo+mucKKC+Lx6igkQKtwMEvWGjuqBc+UxDH89ODgFNLWi+59z/6RMvsaI
LCfhANbooups29W5LBGp8fUz8T+5bosJazQWygGeQ+E=
`pragma protect end_protected
