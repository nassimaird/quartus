��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�i7K21ʑyp�X#�1��°�V�轰���z$�����h2��fzT����݈�p(�J,6�d'
�J����0�b�,X�4��a8T��r��$Ԫ��sj�Y��4 N>sɵ�ܖ0q/�"�1}�Y��`GN�Jݎ�<����ԅ���Րה#P�R�,2��rH�	U�e��|4p��2���[1q���B�_�}�yޜ`���X�l�#�l1�X���W/�۔dE�.�H�� X��G8Irs�(�PM���T�4
�.��I�����ժV�6��$<� ��`#�!0��(Â���"�T����u����v�eonA�7D��
dS�(���A亢�L�-�K�01o3�zv�)n��UJ)x:��C�"�V��4�]���1�#��V|&ۗ���	/�>�ϊי[��ƔL��"7�\��iN���s���pe�j��~˯(53�	�p���X�����@�����~�9���u�د>?p{=��;jL� �b'�N��`�|��b�>���{�����m���
����A%E2�2�8Q^����a� �%jU9�-*͑��~0�G��M����&��Xj�EV�2Z�:�D>W��+�����r��?$[mKO�/k(���-���>Td"'��.�n2cӄ���$�TF^�J�n�Lf6�8_�$M���a���+����O
�H��{�Y$JM��iI�(����i,�V.�h�f���C�(9)��F	��^Ȫ�kM_�R�ƞ�D���:HfE,��Ӑ�t����/C�w[�_���aS(c�g�L��=ܣ�X�OCl�>�1�Q��$8�]��$߻�����}�5��&�~�h��A�,�)|�We2 ll"uXk�����Uf]�����z!��O�P���ԅ.sg��6�N�����b�|�TlO�a�&�=m	��]*#��Z��%]/Ԉ���u�K��,�3|�'�l�DD�.gH~E#�SN/Ճ^�٬�I�c�8 7��s��K%)J���[G2W\�t�x	�� ���iT$���[VO-�,����d%�m�8g�Ov����h��?L������+�����J�P����*�#l�>�Z��U��i�]��َ�fa1�$E�����3���Z-�
��r��'0��+r�HPy�,�dT�_.1*�����hvph|��ɯ	3I8u	��K�C������ĝ�ji	G?g`�؟��/��.	���3�b����"ʈ�A��|<2�E�~��1��j(�}�@� �n���>�5�6�&}���|�?�	]�p��4�8�_�����wHd'jt��#��cka�y�;���O�Y�P�+�8b?�����3L��h������m30犪8H l��6���VQܙ�z1�!XP��n鬓�T!��>8�A�Q�Q$�W&�J������<���1�D{�Ý�|��Lx^�6�X��%B�	JNs-�]hפ��>���V�������B��wi԰���`�	uz:�w@n튶P^�1�n�~�!�fNR���?U�t�:�y���\��Cm�-�XZgƑL`�>��(򪳜�����j)Mc��_k�x>Y��C�ѨD�L���$����z,��a�F�-��0��FM�M��a紵�&��I�E���as�87y?��9�����wa}%�Vs�[�O�E��E:���4(&.�/��k���J���m��`���ǆQ��hG5�U����SB9�Lr�^H0�c��Ļ^SY��ׯ�T�0#�V��48M�R�!����5md9� �^���Q����v���Gx1�����E�����6�,x���H��|~�3�V���l�A����	>0���.Dk�Y7�]�ex�8�`)B;v$��)��ʥ��m@6[�Ԟ
)�WE�6��P\���a���88%�Z��|N�C�(!�eVF����oA�E�:�{T�{<��)��C���\Y
����J9��/웰��=�?̏��"~����WB[)%���{���b/��l�B��K�))ծ�.5	�0�g��<��(�K@I�mzu�&� �������\��LHM�\� \�KAq��h,�s���l`�v~$k���<�-���2"��~w�`�Ú�i53B�)�����C� �n��Ȍ,�����bCn�rD�y!�h��c���tO;���1���ͧ o��U1�) -|=J�u��r�����=	�r��³�3@F)��I�V/�fZ?T~�P�L�H����{����+��c���H�B�q`��r~�=�+s�>���t}߶�qVsÕPM8��J;(�"})�E�g���*`��R�ɓ��Mڡ�"�i\����+��t��%�u��wW�Ŏ��&9f���,����� h[i��  �޿/��U��]�{M����_�0�u���K]Z�����G�	�m�	��jjh� ,W����,�Mw��-Z�f����L樳1�4��4cbo޿k����u�g�k����Nq �E/���A� vZ��z���s�o[=�EOJ]��a@% �@ ���Q>��8�o��m�yV�O��;F4x+7�9#�4IR��6�T�#u�ښq�|&��Nt�sU�ٕz�*ﴷX��x�'�*�_(n��I�9����>�Gq�Ӄ)�@�����T��A��fr�wͭ�(����=��I�vp��Ǫ<���a�Xc�M�+@If6C�B�ddea��1�Ϩ�e��O5�sk ���c���ޗ��,zjE��I�	B����F-e��?Z�T9��*�V9�X  z�ս�$}�o>��s�`���>���P�;���i	�.}�ww������~��	�ʻg#!I)��=3DUW�R����Fg��=�}gäHn���B*�
lt�{
'Pl�	��3A3s�;�9��ơS߂7M$j��|��C��xNe�b�@�ֈ��_|��bT�sN�[cÈC ���{����� ���iV7 {�v��Jb�N�T{%2m��~u]J` Uu)�-iŔ�ں#��}"�6�PU�8�h���H���Q4����>��!������z�4N��d�<�)�[o�Й�Jn�{j�x4342=�D��k5$G���@���2�a%��{�x&���&�DGB��iо�:���Jz���kV?����:c��(Y������6�.�g�V slCTb�p��ّD_�����c��2.��X�|9�G��aƙUa�t��`5�<���U#�G�+��`��u��@J�ץ�[uU��3�F�8�ԅ8d��ǎ��$<�Y�O���)�Etq��Z��ki�h�f^��2#�p1�T{��4S�Ac��7J���}�. �0<2��S��HJ���sR�͉zᡰU�:��d����&*�� �H�b�k����~[��<م$_~\��E���K�_�g��x�0���ƞ�,9kr^_uv������d.g��B(֣�J��!Al��пof������pr����+���jģm�̊�X���_������Y.q�,�`�D�o3��p����۱'���Ŋ�L��G[@�q�o�ɀ�F�.�d\��@y�P���3q���� ��c
��H�!E�a�Qı�>�����%5�~��7<�E����0��*�a"�Wk�e)�T��c�9�hY�p�
 �����j���[e(�n�+�~�M�fP�_��Ae��s�s�">�pл��y{�9�6㨲��pp���p'LsB
Qw>?�ʽ����&���41���|R6jV����;2�Jn][����Qִ6\���ib�c�83�1�<
�
�/&0T�������Ω��1!1�`x\��f��1�}�y��N6���L(g7�<��o��@GC����3Z�/�~0�����>ʥ"h��j����ͽ�g�Ԗ�r?��m���&�����5���������L���m3b�0���I����2"��X�!��\�r.����*�h��b��ⷘ�L�6��En.��Ѫ�W`n�&p�O�y'��=�(�姖��G�P|�	����S��8�?�L-I�M>�{+�{�������ڱ��FX���.B�T}��sr�@�<a��{若a���7v�tɎ/[3\��(�s�)k�-jk����qӽ��J�4`�L�x6�N�
���}\�e�JA���?��x�:�Ca��
hs{92�id�(r!l�̃w��v=�E܀����֮h?�8���%��j�AZ��0~�ĭĭ9v���>�4K�-��3�6�>�2 j�p0`W@l�ssFG�K�Y�ܧd��K�nȄ���W�NI��=�4_,r>Y��}���ۆD�{����,����x�#_�Eb�(#Qs�U��𦤎ꁔQUe�,*h�y1���j6x�Keu0y9����nu}�Qm��=S\�D&�d���f�(hC�뢞ހ��$��\�1yO!'x!q9��z$���]6�Q�O�!~��!�9c������n�L�lk�c��i���"0��u�&{�@�1s%�m�r�Q��5�u%{C<�%Z^^}��I��W&���6^��"2��[Tc/P�74Q��M=�
�,[���'\/_���m.vQ"�89Y�eN�wB�$�%)$C���/��E����\�q���r��#�Tvn�pWw��%"贃�7�%��>C
|M�����XP�1����bz�ʩDk@�M��d=�ꝺmiF�K��`0����
�7��m�~
�S0�^�t���hU者��0:k9S#���0t��G'Mx��*Ա�.�ϡ��*�cw)��z��?��c�x�o��.�Cw�p��d	,�L�wL��H�A9�� ���p�^�ȍ�<���Y)����Z��'��*q74�Ë�z��Xc?<�	'�t�e�����b��2O��D����K��w��3[�Q�Z��`J^a^����F��?o��ة�%�_l��]�*a�6��;3��;{�����P��|iȯ)]�ɠ���g�]�� ]5-:�08a�P��G���u���	��u�J�j��@�N:A��(��CVNdָ,���?V��;]�h�"�J��KQ��@�DD�0{�K#B������}�b�J��t�{����d�#��E�6�G���P[ww�Y	���]C��%�0��|I9gOp�2ƈ%�v��M�Ŏ�bq�����ä�q��rJ�eC����{d�^QBb��7��9�� 0��܁����u�R��7����ڲ��"�&�JSucBy����D�$��?��6M�T�i��ӈ.���E��xl���Jh�ǅ�����1��k��hK�9 ��Gk�!��S|y�r+N�;�?�}���#P0:4�N�d�i*�!�p&�D;Pn�)V9⯒�o������J��8|3��gjumɰ�\�ߝ�����Q�M��N���D"�^ƍ�9Vy�(s���M�˱ �9�������61���{��%�;G����8�ZO��6b�S$7�P�D/�yg�����s�h֎�uA�IE�V}gr��
\R���|t��3^y/��xS;��Mu\П"W~ S���zY�KG��d+��z���칰�;�L�u:J�a8�zrff� `�Ņ����d#��8��֒�6N�)���R5����G�/r�lP���S}�C������8
!����+,?���|u���D�)���W��|��u��[<�_Q���K�]����z�2(�f��v�`lG�:�'�tD�{��s���ćh^t4��v����sŘ}��/W�f�Ia��W1�mKZ_Ԩ��q#V`q�ˬ��rs���=�A�r�4E0�},�E~&�M�R��xk�_��8��\��PiU��m���S>��sY�9;B3��d$ߎ��UD������tI��BY�`��4v��;���_gG�X��j�/��;�E���'�;=v���:T��#'ia��o�����{��p�Ha1,G�S�Q�^ބ���&�Q:���W��,�:|�y4��d'Sw�������9���#؟�J�z���z{4�
+�wg!]�M�� [��h*X�̧%�|���6#k�؄��E&�|%Ó�KV+����w/����jL�>�_��t�o��5���Ә�؄�vB�#�$8f8�Y�#� ��CńXh�ξ��{klp�ٺv����K{��`��}�3��,�qN1�� L��Y/\��a�QE�:�U�PJ�w;�ǳ�t�.�R������[���W�@����<��ч�2Y ��i�p�|�G �8+�p��I|2�\f0f�Z�$ҟ=���_n?6U9Is4/&)(y��K��9�j��a	%�V��#�6
H"�N��K\c�Dc�C�v��d@�野JQ���
����I7�hY�j����6�{�鉓A���@�)�	�� �hu8�����Յ���˥۷]�]@�᥇�5�n�SL���A����C���c� !�p�>��6q���˭��\p}m���F��%�*�\�B�y�Pv`K�h�N?*�/fr��1�=�/su_��;ƕK�U��z�.TEv�o�Ii�̀@�����Zu�8}i���"zM���H��Q�*�#y�>��_���Ff�m;�� ap_�ˤR�Kt���t�w�.GKݢ&���F����@8M'�������K��Ļ��T�-������ժ����i@V���&�nw���y�!��>ҫ�S=�+`�=&F/RxX�e�hIw8���6/A��w}p�����i��X�G�!��c��ɣ:��N{lQ�!�������Q�7�V��cl8u�=oC~	��s�	�Ge��(&���2޺�����B�D�F$��<��IB]�|,�#4��Tۢ�p�g�����l�E#$#B��H.5L�� �1AU;t�6{g�w)(KLR�η�����+��#Nn���g��[��!n���([u]��3ĺ/I�	�����j�(��4���/9��������&����R�]闹u����g{f,��/Uc�%)ډ�F���2�I@�$�g\!�w]����0?w������V�b|��ܫ￞�D�"*�㒡����� [g7���v\rS{E�tȔ���ޡi�8�u��m��bv���P�x��r���	T��r�o��4�IZr]��\Hs�+w�8
l^�H�r�u��`[Z��[Sȁ�ݘR_mT���w����c}��n�H[#�H��M�L�Z �)�ZY��/S^��5~���nTdͨ$�-���јX�'8B�m���H��JI�R���/����A�>I6H+�A%�3j��|�Zk�>���i���s���&j3y����g|�#~���3�/��������g�Uos��[E�+� �2��kXM�iB&��e�Js3Ҟ^G��_�Fv�ܲ�Es'3f�HĜ��]��_��K9���8�ˈ�e=�*�K�Z��cl��8
]��B�cuw�v]Qt�)%}� �)�Ѭ��������}�'µ[�W��wG���E�@����'Mz�}�+���U8"o�'',hrAq�΢5�}>��.�S@���R=�XQ�D�o_�C��U�7f�#<ɪ�M�m��,���&�^J���G����
#,���g��߃c�Ф��]~��u#
�l$3q��ğQ���XS�jL��R��49݌l@�������4�:��Y���k_��
ٳ5ОDR�����<m��74�����*��[���	�ߐ�L%tX0Su�[��l��� �_�Ҩ�Cb�P�K��O�~Iu����5��ON��w����[sIj�ri1�y�Z-B�;c	6�1�\����[m��	�Xqҧ�w��}�*�>vXK^R���2��J�nc�U2�[[�8lq�����y��9/����Zj�0Oe�,YJ���X�P᪗R؇L�rH�G���/���檙��L">BbҸ�R�d��s3��Ҡ�u����?صW.F��[ɳ�I�[%�Ě�}J����[���'�[�?v��LF|MS8�8b2"3��Gw���%H6u���/����.�f�X��7Iݾz�%=�d�W��&�$�1 �V�O��H�ND��X�<P�k��_�����3���,�����I�F�"�ߚ��7��	��i�v�ԙh<m�g0i��M9�G'MN�Zx���'�YV�,}�1�!�Y���_�<!� �����q��������.dy;�������B�O�˸�h��"wY�?�G�����l�߭�I�f%H0�z5!a�����JE�V���� N�vc}2&Xْ*�L��{�� w.�/݄뙰�_C>��2�W����n_�_�����ڈ��LTS���2��S|�ME��m�@�&��B-�K�9���H�Ԫl���9.��}9�G���=��;+èHV�}8��:�_�� ��r�����/ö���7d"eiBg�i���L0Ϭ�¿����0��P���;1��p�(���	��%�+ƶP�.�r��s]�@�-n����m�]��6�ܮ���К����+ vw>�l�8@���4�^x��s_��bI��qk!�\\��I4�s8M��,����X�g'���L�!9!��4�󾅠e��v磼:�-*���T*V.uQ�v��Wq�e����hd�b���u�|�~�Y��d]���Z%�*:�dS#�(��֋Hn6�ܡ�n�?^A[�R�T����}�~��C��?[�Mk�}�iE�
fCk5cn��<�5#����"@�$w���>�Gv)4kmJK��_W��?qRػ3�j�*h����G��Ԡ{Q�5j"r��͟	�u4W�A�n��?Z���������jM��J��ߏH7�Z��R�s�Q����9�i�$��E. W�
2�r������8�u5Nx����A��0f^��p����`'"����K��7XB\Q�ƶ虜 U�o������;�9ų6��Z���9��WN ��ɺj��YCXd��fgQ%�}��t�
ؕS�6���6�<�ڔ�]���;��imS��ɇ����}Ed�nZ}�"� ���7O`	�'X�8�ዬ.��uJS���'WA��]F´�x�O�_�s��;���9�F[���f|��!�h����n/��?] ��$r�	��.��e�D��J�U�/O)Ц�[��U�l>䄕�$��o���I�r-��SNVҩĘ��F>i�cv��=.�-E�%�x���}����Q��E�<�^�����G�+�9}T�zI�r� ��6>� j�zo�?J`WR�����8��=�}*�bӋ��v5�0`
U�~֊4�jf:���$��
Y{7_����c�`3�*�c�e�s�޴��#�&�=Ϟҥ���ѹ"�R���<�����W��,�u0�Ə�^�n�l(u��IҲ����ö/��Po���)��#Fj�gp�Bd�D��9�>��#\?�i�W��H���5#Q0���gq(oV�T�o,x%h��Q���gY��ȢM�ŉ�h�%��P;7�{�7;�D�3د�>_�(@�%��/&9�Da�?��~�lRmr��Co1��D��u
��_��TͰ ����"e���s}�Ц0�A�� t�h���gz�����?����{�^������s ����[BL�˄��1��*��r�f~�A�~I��c7?��C�:l�ᬉZ���H���2FܲE)@�e]��"~#���{�t֌���u�l\r]V�v{��hPuH���{ƹ4E�1_4� Hy�Y�r�N�8U�*��G��:�B���AH�t�Y��@�;͈��R%������Ǚ"t����{?�ӓ�0��q�yfT�_���$�Cw�lm���k��'����$x��$W�x\jq�L��A>��Z������2~�?�ǉ�U�s[�E��u���%��R�7�!��h�A�rp��H+����҈�㛲pݎ�X������TQ��Z��Ͽ+s]^y�/6i���3��u�?�"1j�{&c�fvc�[�-�_�S����Z_��o�HeDㇽM�6���h*�c���pގȲ���U�f`,)V��/_��U���68�r��!�h%��#K&I.0��[-��ʝX?θo�_����A|�,�h6_Eӧ'O�P�M9���V��֔h9��O��(ƍ���v���YR+�=��؀�V�Ӥ_���Rc���n�ߔ��w�wQ�ǌ~�0����p(D
�أ_GX�u���z=-aL���H���n��m��h�F�^Gw���6�aq�G�DvD�`�UE	�#�|l. �&�i�`����\����G��g{
sE"��A=AE�T�8}ܤ.Z�3V��L�V�R��������@��װ���}3�Xa�U!|��A�i| F:���W��R�ݵ���Em�p�=�{� �HϜ���QS�P��Է!�������$��j54-֬��,��,w��:�1ɿ˒��ځ|�W-�yku��5�P�ӋX�)�2��Gi�:v���g�ʷ�Z2s��+�٩��Hs:gw�Q贲�]�]��4ax��b6���j{�lVtE"�l�p��65��]�Ⱦ�����?F�e��p��I}�o���f���9��$���*tu�v�.�#Tr_oY�>p��ӄ��:(�E Nq����O�v3f���#�m=�3��1"a����w����.C����L���nǭ��.�j��59YJ;tf	n��:����I;w�٩EP���r�-V�̳=׾X��j6�֋1���9&*R��V�~�Qw����Ǆ���i�Ø^k���M,�$&��\�8��S�K�@!:[��r�a ��z�e��p���׉)��s��>`ă�%E�L�����N�(�5J�)�J)���3�=##�``�vf�b8@�P
I���O0�U��Q�y̶���`�6v5��B�7���9"�֍p� �[=���?h*��*(g-Qk��RW��ߋi�%��k<���3A��|��W�!���?:�Y�(�"�W���z�uɮ���q'rݝb2�>`B����d�qUN=��WN���X�I]�����2�`a����!�s+-R��fx�h�J��&�\Y�����RU�^�E�0
��ٜ�u
od���r��5���z$�g_�U).dt΢�|V�r��@&vD�#B�o[����vf�Px�F�%6ޤ!��K�2����7Q
��c������x\��c�Y�;�)'h\�ȿC�0�%����{�K��F�z��8�Y'��F�ß���\�Fi��L�Q�����7VӐ-:��=m�l�6�H��>s������Ǹ�����2h�)!X`ؽG7�>@�����X^�:'�x�ߘ����A�p7���	GB�����}�H@��� �bT� 4����4By���2����;�*��D׵q�^S�d���y=�'�C��1�� ��o��[�]�4�*�ÍK{����zC1�uN�K�/e�ero�jM��4��l���?F�)'�S��&&�OϐF�aÃ���F��lDo��L"vK�N÷jn:�oH�/�4�K��c��^�Z�w_d��~#��x�𗘧�M�8��y:#�Ʉĭ�V��_�p�s*��y,#�8���)雖�[�Q%��B���l����`�]Wp"�#� �U�J�7� �|�=�7r������ շ�	����7��p�����lų�{���v���A� I��Z����ESd��OP��;�����m�;�c4"�-��������Y
�>���f	�c?����&a¨����#>��3���h@8���s?���BJ;��g�OTׂcx�!��KG�p"s��2{x���k�W`wʊ���*SA�"�C��ʙ�sq��*yd�XGh�W�p<g�URD|̸�@�m}Jw	����v@�1x�<6�^q��*~���qN��<`ٚ�hɃH�"9(Ն��\���� �Z�:�y
�w,�u���e�"XG��9��qf�)�_<��O�!�`z��t�u2e�<�cd��n0=Y���B��?<�O�>ϗ�$(8OO��{�Y�� c$X�K@n`O�-~:J�L���v~�R�f����(Ko7@l&�5�ZJ�]���h����%`������[MKk��&R���;�"4bI ���;�{�hj��pG�}�{򅓸�\��4�<'���m_E �����FB`TW_����9�Y(��c9pU�Nm��������H5����UoB�A��������A���Q�PW����1,
�9Sxfn��魸F�<�0܈���[+	*��#�J��hՕVw����5�Jʸ`z�h[`��=���w��Q�@���� ���R��)���ˌ��g�=@�ך���H+�kԦ�^�o�ڼ�b_��k�X5�TZV�bY��-W� [%�4�s�y����hc� #���_�G�a��Y�v�~#䛄�QV_��S���$�c�Jv��tn����� �c��#)lG�����-�2�z.��W��"� �kX�+���W��/.�`+dC�gc�~O��l'6��kx������6j�\��絆���s��+O{���l�~n�m?ma�k{�D{	}6�,�5f{>:��f/Z���3O@�݋¢��N�@� ��f�]�Hu��V� ��\K0y5�a���F��-���a��g���������s��n,�����yy:��}~=��7e=Lc�S���������-<5|�-2�A_��[�>Y S��O���^i(�cS��y=������w�6���cl���<������b��#�n��0��`%OBB��O���ښ̀��WCRg��;D��\e�Ro��%����C�j��Ҩ��,b��2�nӎ�pE��Z����ߵpN#(��
袾���c�N�������IH�,%�	b��p%D&q�cc;�>+�t�[�)i��҇���)�<���c�~�TY�@�(�M�44���95�4mߏ�w����r~����pږ��#Y���['7m���$��k�2`�$a0�2?�W@씹��3P�=r�h���j�ێ��K��\�<SV����):��, ���@w�
��L��ܝ>Z� dW��:���� ��C�#��!�q`��>�Py ��	*!�W�^�8�'A�'oYh�y���R�A����De���gm|��t���c�]?���6#J�R]̱����ՕES@�OAO逌�7�xH�VK�,/�r5�N:2���L|�bX'���v7]�m�J�� � �j�:vj|B���%V�cˋ�J��/C��k*���V����e�=G`�.IY8X��GO�h��p�4$k:�]Z��3>I���;+w�W9��1j�xnk�u�za�[<��p�H�Վ�����b�bx��0q�Rcd�`	�^}W����X���J g�K��^Mÿ�k!��_6��rf�K?1>�8��N�+<ͭ1R,��3[�46/�w� D���j��D/+����h΁Ŵ���8� ��/�L����YD�ca��1��_R,�%�~��䡭�~��#�! ��bn�A;��[)*�{m�ѓh�<Kxc�ᯕ�v��;xXl��h���7^��b��JҖ����(p<q���d�L�����!�Ʌ���f��+�Y��I9-M�.�D���2D2@'��� %s�?3��i�jiWQ�C���ە�z���εa/���ø(߲�h�F�rcԤ4�x����p=Ήi�酭%Ս��.�¹�������De�Ƽd���r�hN��+?�6N i��~B�Eb�OCG�O[h��f�OUs��9��v�$����o]��7�����^΍;�`����5g��� ߴ�42��������"�V̒?��L2�^��ĘS)+:�#hfӐɱu$˽DY*��M2����|��E�B�7O2^j]'� �`���[ӊ������J2��c�|����o���$'�l�� �ɹ���i�x��uj�_�����|�7�W�����>���Rh���_%	�n{	MN��L��Eǎ.������<R��D+� "���^i �A5�'�Ѐ�K���<������D���ɾ�q2<p�)�7F�<^�}���hh��0���޲��dp:�䮔�$�h�q�~��"&�&�>Z��1+��Ƒe�~x�n V`�~�$���1{A+8��A��?��.�uЇ�mf��"ũ#����ݺnu�V��d�6����^0�&�� Rʍ&F&�N��3y<Q)�� �[�
n7b3	kLξ���̢z�y���U�[� �=|�ճ��?�����e���K�U%���ɨd�R��譪�(����	?�W��Uy3:�򄁚�?�%UNw���_�(�*�2���G�w�'G��1��{m��A7~j�`N�q�F<gR+`Noج�Dǭb��[�t�����
���e��[���궅�ك�Ҝu����f�F,���-���?dȻ��J�B1F;��},���CPD���)j.Tt�(�j��л�3h9r�ڙ����r�����<�6j�[};.HKdº��P�W�a��W���:̑��"�]�o#cQ��ھ��6��I�l��/�Y��$%g��:1�q�>JN�K�U*��݈�m�\�)�U���>�R�T�h�t�7�)�^���Δ3�O�g�lNQm(ԞQ�����ЮD�y#�3켾���d����n�������&���<������
3���=�8����Y�6�i@S����3��Z�.v�1��6��i:^�V�s���S�=o���$q�	�`���`�3�x�#���வ��a�'�i�[g�27b�\�Zf�J���
�Ŧ��CE_,鼘����'n�"�����~�thj�^����Ċ8���{���Ж$q�]�0:b�A?��`�<����?h�O��F?%�9�H��XJˀ[�P�jW�k@��I������=~���"f�ՖP	�.��x��������>����5�Ξ�ǛE��.
���!��xU�1�eW}��JU�s��.!]Vu�ϗ�M{@�Kɱw+!pe�罒�;x�oѴ+<�y��M���I�T�9��a�� �8*�đ^_f��u�˲��}3J����P�5�ޱ 1@��E��IR�hJ�?��&����~pk�3rW�4zI�@ct�'Jf[Н�įc�G��я�2m�T��*�T!�J�gcL)yaCnq\IJ�+��l����Y�I�{��u���XZ�@=?�p���^�I��(�ׁ�/Ι��on��G�C�:[QN��89Sh�cDΪ�Q�0��o3��(F�s���ł�0!��k�DHo���O5������p�H]ݍ�\0��m[��O�� ��&�,0D�>�Ϻ�^Z1�))��?&��ؚ��1++�:6� m�����(�`��/	�*�y:N|�7>���Y�X��f|�'L*�X�Q�`�ّ�}ȯ�J��_DP�Y����Q|�ꓣB�zN�Ŏ�T����͙<9:芅7b����?u�gAw��{�8`緾����bm	�k�aD:����}�V]��1��Cf�}iQ��@��ސ���F�Z<L�/�@5kY�-��t`b�nqD�\k񚢞�J5�ˑ�	���y�#����&�<��4�a���D��z��i,c�	s��!j����"���jנ^���?"}EH�~�;���U�^_f�"���sP�~��A዇�V1l�&�-����,�$M%Z�v�;�*�FI)�q�����	������--4��ϩ�!~��ڂ�d���RiWn�HS���'�*Lͤ��&����N�/�y���z*���B˞���D��RZ����[�y���m�C1YN˺ʮS�L��|�='4|tc��ޟ�7xmN��	;q�5��3E2].⇒9�wF�:����@WJ��ĩIlu�J������'�ߺ���³�^�Q/և�ʆ�Toiɴ٪ZM��J^����F[}�mi�<�:O�� ��"v��1��_�ݪW_�atE' _}����m�Qh�d�bb�����Ռ9W����S�s�<;(rz}�rQO�z#L~Vٹ7$>�S�R���l���!K���~�+JX&[7[`Xs��!R2�/��M�3��L
Z]Zа�Fo�W�PIN6j:����֟�#��X�XV�DM�hV���w���_j���
�T/B��;�lXǞ���`�Ղ��rkS��;�)�g��tS��j�V�����!Ȯ��)��3M�ڕa�A�E[L��x��|h�|6dC��%�푩��V"��MPx�&4=4\�8Q������Q��R~� ~��̿��DD��Й�g6P�����fdH�i�NRgl9�n��	��r|DG/�S�NR~�*1�8��l֕Xby݆�D������+e�餷�#Q�DAFECn,BuH?I��VY��
�5L�����t�4��%����s&|�17~*�����Lt�]�}��um�欺O������&��Z>�A@�
J���ԯR���v(K��M+8�Tq/v���N���;2'�F�#�얉�s�k�0/#��@�1D�����#��ʕ4vd%�ʸ��ybw�}O5����*s v�%������)��8�3����Q�V��%�F�