��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�˅������d�xp� �5��B�{�	e��Hk�Z�徒��{��\�83,�p�)V2V"'������'v�{��A��L�J��ʖsk�eRGAO<M��a.p�b��@�@a�;Dep�r�p	1��"32G º��*ڦ���ƫ�r`�c�}_1������	H?���}� ol4,n����������\p�kх���F�y��f�T%���^5�����8
�2j��pVq��zK۴N��@� 0 �	��ev����m���z_ws�=����#͑��]�Ţ���FC$����
�4o��3[�Y3�v��� r�'��̷�l���S���W�v����E���1��_���Ѵ~���;�ﺴ(ܢ]9�\h-m蹞����3���Q�ó�?�A����Ƶ�̟(|����g��~�Q��6�tg��}Q>�CW��k�9����ΨˡI6I���OS5No��k*�D��p�(ޚ8�5���6����I�0�~����ǏFA�2�;ҩ7^&�'UNg7���ZE(�����
J�E��B�:w���'���W���;/�R��y�p����r��Q���Ĺ�х��9�v|e��E��(h�,k�NNk��xL9ӌe�9:-cJ� ,��[��.����r�A����eA�v�)����8j1�A�ƨg���o��������Ƨ[cP��^��r�Qfm&�ؿ����I@��3Ml����Ɗd/��gčZM��H|,*-�r|��bo{��@C��P�eV�c����C�u�μ0�3�,������N�X�WBC-���2St6�8� �7Uƃ��rX�p����4�P��V 涱�P�n��)\��*՚�S
��V����RO�����d�׾�����P�䈾��*�A� 3�b�S�|�>|0�X���w�g�g=/�CmL�~q��4|S"�p�Ń�%Dd��E���5��@}�n4��`���/�z4�5@���Y���TZ�_}�N�f�%��A͉[	���qw=�Jr�L���=��������n�,P�U+��u��Сs�I�*.D��3����,@_0�B��$�uC����X0佁T3>�?�)hx5���kd�K�H+�6��JЙ�6����B�
������B�Ġ����������,���|p��&n�G"�C@���_��R��7�GGgK�e�3}�Kc�p��GI�X�{�q�W�{�1���;�6:f7���ױ':�ꌤ͆^�q����:��a�<�=.&2O�0�M�L���������6����{�ؽ��)l��2��[F�]��>+���ݱ�S	i���z�J�s2�S�"��P���g�^�޶�� VYe?�����d�H}G�o���������4��'�^.��D���o����o�)3;����é��~�r�&���ߚ`@�o��*b�2.>Vh ����
R�	�����ba�7u@_�
���X�x�
8k���# UMb*	��0���?�6ʤ/z=�f�b�����]o�jk�c����Rӟ���X���z���"���*�0Q��{b����ZqnT��C�T��5�gRy�Meh_��N����9Yy/v���Iw׿��O�'|D���ô��9�L�EdR��w����?��׀���W���A���"[�D�m������L��)$̤Y��9�����A���!� kb�L��5Q�mC�A�XG�H:�e�+���#�w�x&b��Q�2�I#�2��8?�A��5�ӮW�A2G�n۳a��:��8D��kS� ��L�d�oX�锇�Y
2y�q$��"3��1]Xݒ�'mmOR�%����� �
ħM)b���ʪ��+��sc�������r;��E�y\"&x踵��.�BD���z�sJ!�v���l�^#*~��Vf��u�b���9r;�ߟ�^`0�sZ�������fH�lo��ꑵ~��
�����zg�|j�(�`�)�A�yi�W/��^��9� �\ªU�Wa �[�Z2K������*Wˁ?�r.^	�Q��?(��`7�?&�$��KX�=e�	$�UA�
�L�$�[\B��T��~��G;���Rh��ML���7��ܕ+���<|A�rK��B �>�s�>���[Е��2���������=W��r'��C
_v�J1��	��+ =c�˯�qN�)Y*���r��\վ�*�ժ��;p��+B�X8�h�)6��aK��6�Ʉ�=&�x�U)��H���۲��~4�5�J��,;�m�أ���C���L�&�����Q��R~�*��n�L���[��QG�ra_�Zb��LR������=g����bh�E� �o�غ��UW5�f���@�EB5/t�z��V_Kƌ
�R8��wڤ^|�r\]�����>~�"�ptU!�lI�|Vĝ}�&����v���dl�cTH~@!�|���RAZ]�S��T,����E�\�>݃��}�D$�>5&��[��Zԋ��zL��&:C��g�����<3�2z,��M��\�r� v�%b�S��-p����n�T��W+MF7'|X7��]�������/AE��d�"��\�L��$�ɵ��&2��=fFS���}�x�8�jmmȐe�ؼ��L���JtY����OӒ{���v��6R�����._|P�����* で�*��.jL�����bW�x�"D{����k�i؞�Ud� �HPR��)�-6�O�̖� �P��9��l�V(��ݛ�I��j%P<an2!��"~�@}ql��6����`�K���?��4ͽ�ꑋ���jO����������`��3]ˮ.���L�lI�!�tlŢJL��_FF�Dŕ�[�/c9d�7=��I�V��!� �̾�]���E��VcF%M��p���D��[j)��ђ'��X�As�������W��%���%�V9ߥ~D+.ez��F"�EUi(�P%��w����E��=�E2yq�Ә�E!�Ⱦ.���4�xN���O`ȡ6�#$�&E��s��L��c ��}IV�~�jfuQ�Z�B�UJ�F��-��=�{��.h��p�F&x���͔�#�34O��17���k�{�:5ʄwb�F�������pݻ�����rQf{����]�r!)$�Vͼ��ӻǈAt1�0�}j��G/T��<�۩�Y�*=F�lgeP��K6�Tш�*Z��l�E�!9�e��0eǗ��DL9��Zs�!v�
�$�wꩁ����KԓfX4(x(JȰs_�N�����$�����U�?���v�� �ּ�����Ȗ:�kF��k��z�P�'4�#�=�lWl��G3f�,��fB�(�#U|���upR]����\���Զ�[l�m{'�M[U�9�	�"i�j�k=�� ��K�b'^��-*eH����Rm�@��4%r�'��3q�g?dn'�A
��@��&��]{���uVx��I�BQ]���h���U���vn�b֡�|��}����=���Lr��lP\��K����G�:�}���t�>���+�c�)�,][���<�5���,ߪ[�u�ޘ�Y���P��C4I}*&���P�Îv� ��5ZW����,���7�DR�Af	,f�P;>[�>8ФsM��Et9�GOAIO���<�8����z�Y��*�`_1����C��ԝ��6lu�m�QA��"��j4(���&q���
#���s���<�^)�v.�Eg3�0��LP4��N�t΢�]��B�v��inb1Q튳�s�pK���oJ\����AI_�c�v�"S�/ຓ(&��O�;�3����?k�,F��/ �:vs�[l��[Bu���*��+��o�l��YN���n�,O��9���� Mo�>Ҽ��}*Q���q=7LH�c����)���*p�_�`��da�1,9:"7��f1�1k+�@5���S��oM�;PU���9Ve��bYb���#����6-	��.߇��hOUd��Px˸���D:+AKN���OD(��
����!.�}����c�"��@Lϲ~C,6R`�v:��5I�}�e�F��#���y�V�0/��a�j�Kc���uKl5�Rb~\�T�ҋ6���hK�eI
��T���WJ�n��j�c`ӽ�;7
 Z�"D��K.��F��W5+ꌕ~(�������2��֊���w*�0$%��Dw�����P��?�w|d�/uУ�����*=w�_vQ��;)_Q�Kt���3�Q��\}�:)~�]�B�D%�,������/x$'s��(�*�J.������K��A^��"����OJw{��$�7��%��H�D�z1�q�~�!�ư��$=r?"�J=Y�e0�TaG�O�*�h��Ob����:�Ḫ̂��x����2�� ߲�p%l����<�06M(2/VT�w�({�l(}�ɯ�[���e�u��]}�d7�qt�5r�τM���9�ѧ������E)�~n�`ԇ��� @�+���N��8��Ŋ�R��D�ʂ�����[�`�B��F��v�
�S.�1G-Y�P�9�͖�+d\.����pjv.:��	nJ�o��ߗO���x&\D@|��8fe7��?��J��lY�t�=�Q�I	\߹�����j�lǒ�y!�K�B?7�в2U��I�8��s�/B��N��HwsȓSL�Qp���D��Lۖ�(_��?��G�xU��)>����٠����6�뚂x�d�����+orn'>���GS�t�Jp�%�yq_�/0���m~.'���P�:�͊�{}T�m����P�9��������gp��4$�i�%ћ�@+r�*�@Z#Oȅ�۠Ā��{���1� ~6luuV�3y��zm��n������;�
�ư\�0��U����q1��	��N���{�hY��(���p7��
��������D'�^a���^�)���u{�owu�2��� 檬�goxgoQ>�����Xȓv�����r��g�AC�$��e .�a{�����&[}�c�P�f��7ܾ��/�?�ޣxdq6*t�r����'���0�[fi��,�`�q%Pk��`X�86b�
��Ke��)���2C�j�]��P�F����{<w��=�^�t�k�گG��M�G6���J���M��Y�� ����j�����*qW�\�B�ܻyd���$tc�M��I�q�.�l���o��>S�CG�����\i楿���$$�����C4 $N�Г��"p�P�h�6:/\�O�Ռc�,�*�H!u��4z4� ���r՝/�.�h���-���M�K��pI�o�E:��OS�hŴC�|�+a�K�|(|3Y��+�;\.GVOJ����P�H�
�������2\V�DrU��Ǌ����[���z����t���{!�m��WP��#6�zk�8K��������="�����v�wu>�Q"c���#��R�s�t�E���m`����J`���<R"�
�
�Q�W��m%��Y���=�b�3���?�.A�e�4�Sv�̥�4�!��6#z�\���r΃�"#��x;O��ߘ��t�2������&�k�?&�r�7�)���n���IY�>޴�l&�^^�Ww�!ed���S�V�^{���2�"��s�u;�/��y�ws{1�;	c�`᭱;%���i���#ɻ*7���/	d������o ���@�.��Y5�%����jj����d���r[��H�7*�E��~�WlWY�Lf�=��l` B[/��x�mP�S����y��VCF�N`�YTC�J�ۊmb���D��������Z�shS���M�7��
���,���>���AV�[(Nb1j�ٞi,�χ��u�G�uO�u�.̰��L�Go�8��Q�2'==�4<� ��� >	ވ�d�������K�@�Ϯ���	q�ts�E_W�Y0�%����r��5ccWD,	�P�-;>��좘�l���lwG/w�#�ʮ�ZZ���pu[~�%���/�h�e�������O��9��2�ߡ�����@ Y���ߎ�j����PK�w}��CJ]0q�(=v���~��(��0]�F�\��O��x���'� }*"fJ����&�L��g�/`��K�*�TZo�4��W�?��ݱ:e�Q�l��(�7��q{�Ө���5�6�143�^2�!��@8�_䦉���(���Ćѵ����9
9��n�7�ń��ǿ�M�H���XV�~�Z �D%Ӵ@����¸Ғ�ݍG�´�Fk��!�|��$w�c����,��$0'	�8��lK�2z��d<A�����]�;hf}o��4���/ɓZ\&ǌR�8%��z��n}$h�W�?5��Ȥ��C�{be^���g��z�/����y�S����D��T��p󉅢KT�rr1l�:�x?%�1邌���燶A�M�Dkؽ����®c��H�~���2K)8V��$�A84��K�]3.�7��Z*zD�]Y���(�|�S�B��'yBOo�}�֖���|��L?��Lvu�L,���Ŕ��^�,��q�Yi,�V/#o/��?�Y懑�̈������φ2׻H�۠�>���;�:��X%�l�%�/�>ྷ���Kъh�̽I�t�+�hr̈&E�
���r?��O�B,0	�؉+7]ulv[�l�\cϪ!�A����0M�h-7�]kQ}��SN�ӳ��g|�Cf�T�=S���Oa�Eo"���?���o|"��oi|Qo7i�O�E�Q�%��F�6/����Vp�"ZaC�t��k�>�8z�i[n^{׎'J���r�})�5� @5��?ʶȭP���u�����
�K,6sjQ�;����	!���Tc����J������gb2���d�d�Q�S��4�DB��S4 kJ�U����������}����%f��&:����"��²��|��B�'�2<�� v�l�cUթ��JEn�o@�����,��*��AI��Ć�ߤH���B�]��s�_cA��2'�2�,�e�7U�֍���=
;5`��%;���v!+Ku�~�z6u�)/����NL �aQ��RA��/$\K^������*sp��R80�x�{k%kf��?"���Qd@���!��uT=�hq'=�p�%8��8n�L-.;B�[�V��E_�'���yi`��$q��q��Ƒ@�4������!����k����0&��A~Ui�����g��h�zӟ8�C~ą�9�_	��ʿ��c�VP'a�;ʙ����ڭ�AKh����[�����y�ղ�)`:�r�&��k���i��}o?i��l��L<��V���(
[���Ōp����<!M�������6y����0e�ԋ
7��xL� ���-Wm�g!̞-��(��Uz���5kB����ϫ�XЬ3Mʝ��Y۲�k�Œ!�ˈ�%~���!���/xM��i�?�ڋ��9��u�I�ݳe�������5H����_��)gQ�M��
f��Wm����kb�㒕U�9 �W���\t�z�*-Gy֣�iL�سy��%ώ�F��i��G�R�3R��X�EM�ˈ��.��g��z0�����&�Xb�{�m�:�^�L@Ns�yR)'Lw�i|�ڢ4 ��76Zh@�'܀䑣�ɔ���6qi�[J\�h�r<�}�����6�c�?��M��%z�u%Y�YY��+��\�v<��9���o�A�[{CB~���f�?Blx��ߛ����t�	@�C"�oq���=(�i�xCl�ڋ{�LTlh�������"�MaJ�S/W�)c������8��*V� ^ΧNp/�j��������OhG"S�����=.<�C�[����s�ΈUTs�3���v���?����K �cs�85�����{lW C�
����A�p͑W��e� L'���rD&����}�7J�TŹ��Y�K�ف4l���ʬMf0͊�������k��!����2�^0��_=��6f9���}��0�8�0-��J��P�Oo�e�QVj$������8��#���K��8S6���m��p9�����I��uk�6��b�c�p�b���@�V��E���)�#�g��j��7$F�N,6ڄ���.�ߴj��qM��+5X��}��`�I3��c��p�:��H7�P�G��LN�d�\5���tY�秗 ��B\�b_xO���i�U3_��p�M����� &��Aדʇ�s��j�/�s$����wV|�3z@�g�&�T�&�������/9�|CE@>b�R�X�V���@�6D\�ڭ|p߽�L�w�Պ��Ќ�*a-t6c����u��M�ϩ����@�-w�ߟ� �'��fE�d��J�.�� �������G��ױ����lb�5r�@�P���Q���˙�[Cק���u��'R`Pp�ʊj�����{���o7I_R�n�9���Y�E9�2C��l+�ĩz�fK����"?�㎈��^ �CZB�U��1Hc��.[^&U���?��I��X�Q����ً���(�2*Y<�ܶdM���6�JM�|�L��-���g���l�$�Z1Qt�*;�W���%��r�I$���Jʸ�*1�Sg�FS����	&yF!����A�AЄ>��*a�9^��7I������>[ ���ŉ8ҡ�1}돕sI�?��mr� ܫʋ�@9����!Z!P�p�0[��S;��Ҙ<�jM�a���%m��Uh@�5��Xl8;�P��B:-�U��uOLL���e�ue�	n��'BW%�5�h�"4��gp���n�q����M_ۚ]c,7K�؆O� �,[�*���AJ�Q^	|�rɟ����r�}y����=^��&�(
D֍���b�E
�I���ާ�⬨L��|�Od�T�7i�-�PiY�ϖ��򗑖2�ޠO�����4�/��,3-�;
�� #1��X7*n��D���4���ףz��mT�2�f�o��g���Hl��nX�#���Çyk*6/��E�(��O�g����*��8{w� ���h�2�ɒ͂�����Շ"6l�=��~:a�2�H%����V����"-ÕO��u0�7[��ꮶ�|$	�A�d��� z�3a��
��Զ���h
F�@��~ZW������+�ߘ���+�O�k�*B��X��}ƙ��k���[�rU"���������nv��*e�U.����p@H�#�&z٦����_VG�2>�g�������oQspb�`Ele�O�5�0r5����P�}w�y	>�����)�P��iC����I��c�e@����M�Q#��^�o�j{�� �|�%"�9,lI`���s�h`����@͚ ��/٥*��Y��7L!H�6c5�@(2��^�;�@-Oa'�ĺ��}̖�"ҁ��Ep L���\/�!S�!�Ϲ��^��H�Zg`S�����y݄�y����2�oa��s�r�T�A�w�Q��$Q`���Wp#w�F>Tn'�JB��?T�5����C9��\�g��iE2��0��w�-�A��Ur�s�	n��p��&�%:��K���G�<	^�	M��.	�F+�n�(��#:��iY;���y:�+��E�.|��l�X���%fYk�D=}�K�E`�2�M��ƪkL/���f��W8��}���e�n��|oi��^?;�F1:��v��q��x+E�������������c+h��fV��Ħ��4Q��^KKBW	�0H�Y�s���Ѯ�)����0Q�aՠ��b�~�h�^�Z_�x�J6L�;�?}ݑ�b�ҵ��?�${�!�y=�t��q�@z�� �s�1���jh�v��	� �����9�[� %_O�P��j2��Ǔ^�]�W,����y{���X�$ޯ�b�*3pa햁K�u7yIN�P׎2�m(0Y�'#Qqd9�Ed�����i0H�ԉ�Eu��p�>W�_Y�q	K/æ��
?k>���!͌#�D�;|�Jlm�~h���uZbV�|-~-�%\F����O�I>Y�ɻ1��C��YR�����a*�'�{#I�|��P�MJhM�"#��Ӊ����}҈0n��b�W�@]��J���64<@/�$��D��KE��Iž>���Y�H����3K��<L�|M�鹂��&�= :�~�fo�.Gz,uY����T��U�A��4R,5x�p�Rz��U�<�nW4�q�=1	y�Zӵ!C s)��t{�5����7I ���bͲx��A���'X�+�e3��ɤ��$�iPD�]�a�a-�g��w�O}����%�ck����Ye�%��
���m`_X��A�A�W�͝?"e�g��2��Tr�:pa�������3:��(��y�����Oo(�;p�c�ќ���3~��K��COO�C���x'���`$곢T�.���P��G+>{�|'D �h�4o���Z��_��?3ē�7�;7��V.�3�k��P����	Hdz��@b��,�9�{̩��TM�`�ky�8��	�����W�@�F"WԀ��g�â���V��|T�!����-K.1��F�Pe\��_&M����cĳ�}c�!@�!�L�Y_���JՑ�}+*&����n�Ш^ʗ���\I&���P@��ެ;e03�k<��q��~¶ ���n�Z����,����.�H(�_���S�m>m5e˞�D�}��$��<�7< �. p�9�&B%.��{FRk� 7�l?I�ʵ�5�Yy^�d�qs���s�wj��ҏK�cwA����)�xV�!9ɘ��\k�j�hqFY��M./�?�NI���	�*�/^F?����3AX��I`��H��&��TJ(�c<2�C\�>{��**Ɏd�"@5�C7��}�$FA�/��h�tg2:L~���}to�肽y_t�?��FA���#:�V>�V�Y�M�l����rŖ�h�L�-�m):��H�mp9�S���x�P�_�
\F�NH�?��k�������.1�ʉUX�6}�F��
����3g���*�}�3�˳������pf�|h��]���w�J"t��A���i��4HI�.|k�{�����lvt\���z�l�-l���ק�O���=�F�)<�^�.h�d���d�p��'F�'+�\�60�N�Z��'��ڲN;>M�wH�ݻ����+g��\!O��][NlM���'���k��/tw槁8����Iʲ2��#���	,U�Z�k/����[��?�N��K�U����'k����x���(ٷ��k��^���Hf�>��g�`������D>9 �qX������K�tI8�u�.��[7���)o��a�>�$_p 2	(V2�7R���Ε�G���	^%=���>ӜWǻ� �nS�>�H�4U�Y(/[7���KxP��X��/��>�Fk웿4�O(~�%�������m�<�����xb�`VJ��ڔ��Nhp`�:�d�!lP*� NƇlK�ٕ�z-�6x���9�h��P��l���3�3/�}k'O�9b�㖵M��?���z=-�^k��v`�B>�����@�o8�#�4%6��`ld��p���C��'� �4��g��}P#��=b%�R����.Ed��	?#��`�Tм�C4�~ĸ'ES��Ie��V,*r��WsI�m�A�����o"9���t��~���%�F�z;f'������Q�i���m��� `�*!���2�2C�TB@a{�9P
�@�+de;�(�&C�LH��?�����{�,��=��X���_VE�B���.eH{;����L�+I�vS#]n
�>,�b*�l���g���G��J*څ��Ղ�:x\4�c[��a-�(�%�$��Z�B���#�[��X��鹡�����;��T(~�Ex��9���aD�!'\�}k,\+з,�^���I��O_�[NԢ�2�~UzgY֐QQ>�������c��z�be50L��ȸ�D3��u�<Z�P���1.+"_f����U�|���L_鈶ޢ���bq����Iig�}=�4YRa��c�'�~X���zQY+�zޣ��n��bD��� �X�ג�!L�A�M� |n� ����W
b�E��Y����䖶��?+��A+��k�-8�p�S�b�t�'��`�����F�=��o��N�P���ڗ9a���@�4���Td+��C�.����N����}�e>���/�B'!��!�Y��
X��M�K��,]q�/:ha��֓^����Dֽ�39*�>�D'r6ep��Ñ�R���[���fK4�#v?%W��N��H9g��'D�
��'�Bv��QE�%��rF����r�И"k$�&�S��H������X�R����ė���p)g��ө�l'>k���~��)++�6�@��oj[��W��1$���H�G1�Z���3s��@�:�٢ߩҴHu�}t��I��^9 �x�:˵M�W�(�
���y��8t��j�x�E�ړXa�lBX������6?FB�M0💷��_|��y��SHX���;Ei<���y�X1���Iv(��>GS�p����ŗ�2��FA�������K�;~�</�?}�Z��\�Z���1��?���>x%xu��@Kxu�p�H�>p[���Z	>a���߇��3�MI
�)�bJ6w�)�"O���"����"����.�rJ�\
�y��P ��{lM�\V���EX٦�*�*��6Z)�ff8&Eq��r���!LB#<8?�pW�����8z����'1د����WI�m�nw{M��f�>Q��}&.UfO�s4��ve�ױ8��b��{hχ�Mk�c�4��kY~p���WB�|<eǉH��@l�j��免���3H&����>'eiO�<*e*zt�Iy�������+k�_�&��\��,~~��LBk�u΄tQ�J�ܴp"�Ufj�;��
Nq�e��Y�����cB�Z�A�
�p�V����}����q��f�S�.VӃJ��QLu�`��LK:2-®�0�쫨!K�/ <�SZ���h._ ������>�uq�������Wx�5�rR����;���_����zf�YK��^�(R��>e?K�0�5������(������ՙ���`7e�����E9�2��RZʁ��?l\���L��A�qn���/��,�j5������X�'�L����\��[��#ЩaWe�waN:�R:^w��*�4�Ņ�l�)�p�j����9������u����$��$����o#ϸ�,ӳC��3��}@�����V�C�O�7��iQ>οJ��e��Pѣck  �E<���i𧱞t�����4`��$�Α$�i௻��S���$����9��9����� ���P��ǖ��š�����sZ���
)��?\e�O��f ��N��/��a���2��/��څ�w6�y��Ix�ȋ��E���E��۩F�}Q
\�OQ�����'[CH� P�����{R���ј��!�A���^cR����x}f��!��|��f�B��#��.L��:���ZnO�@L{�Ъ5�d�s��q�A�O���ќM������5U	���l�%�c+>E%=���z­���.�Q ϯ}Q�9F�IT�z�hF�oH��K�
��6/�U��8M/)�x{`�YU�x�JEK�I�-�W�OR��P჊ O�d)�O��	|�31��WYV��cljϢ'��ꈱG�[�m� �48��q�D3̴�G�li`�l�K�sH�����:Bi�_��dFnX&ut�a��R1#��N6j(�2���'!w�EUϋ	
_n�
L}^��ʂ�S6���SU�q�p�:%�~������f��g!T:��k< 3a�,��-�3IY��k3z�1O?�(�#h�����
����J ���G�W���)�$i�Pz�X�9�R0`��&�Һ[��^������YO#�C+�Ogy�Sc�H��ob3۪��Ƕ����*��yQݽ�k�{Ԩ�<;"��RY9d�Y�����?sL�k:�}N�j�	E�T�/��ec��B`�qsh�oJk�N���겠@
a������	���6������&�Tҿ,��^����B=��K@�d��$"uV�S�ܔ��O0I�b�]�y�����9R"�~���uE4GyR��	�:�sԜ����x�pi,�f~��zB��H��-�~g�|�u��Al���Ga^E�GtQj�Vht����		nG%Y���R�~���q�E�x�7�&e�;D^�Mt�,�AL؜�Ɂ���pL1(�J�_T�Q� X�_����X�Bg)�l
���A��|��6Qq
;M�b:��F�)����5��6Em�=p���ܲQ�@`ܧ�=2�Y���Yd2���K�	��<����\!{D��Ew���UB���{�uh�+$���;w�NK�2:ٰ�S�p��g��25�c��U��7ɼ�>`���p�φW�Ar��薟����|���B����}$J����ʰ%4�Vi��k�׊���ܙ�m$�c1�:�	�_�(��kJ*׳�[��ې+�KQ��9�3�M�,6�)dqX$0 E(�r�,��ZNf��;Nܚ�FٮF���CQ赐p�P�	;��O&T;1+�~��'wв:��MP��� �x�}��ص����C1�&��V��Վűz4���c��JIu}�ѿ �k�p�ƽ$j���w�
X0\�Y�۽2�*��(��<�%!���������Pz�`^�:0�,&t�s l(��.�}�MR�[�oEá����"}�X��rzk��E�����x�8��J�վ�(Ha�q�Ff>S���e��ٛ�W����n>Hh���B������'�e�ʝ��ę��2�_��əp@i��aw[���gM�p-�̸F�:K��"��X9����җ�[u�M��@��Ҷ��G�/}8���sdGtϙYt�^ו11Y5��#C;�{�x����?�]�A@.KH���N������x�Pr{�)<o���	`X���F
�柰�g�t9����s�qpٲ=���B��Q��RZ-6zVjn:�V����J�2 �V���������UeIj�<��%�^Ӧ�`��xH��*z�
�p�p���{�q�~*V���q�� G�3����
��X��_@C���&���M��g..�V��hi,1�+B��-��V�0�������e�u��𴯰�o�kDn����C2�����?>���K���$��6��O����7�ݟؐ�111T 7�gM5L��w������(>���t;)����A �*nь��z�n���=Q#��4�����|�3�:�|�����z"��������'W�51����\o���l�<�a��0C�y�]�f-�-�T��_s`0oR�$w��9-�a�4*�����X/�${�PyԺ\���HB���~��o̸{�,�*�����ی�ks����}�g[��h-��3L��ײ��T�����h�F�P��>�I��߄�Q��[:���`�n^�s�r��q���4�4ݛ��	�|��CH(���.��Q�-��x�>�=��^�p@ɴ@�gQ���Rߗ���]��+(q�^�u�l�%��%���I���~�y������M)�T���hj��xr*��Q�t��}�YTm#%����)���p#�.��C�߮�?|�Ϩ5�3�&>l�帠�&;�t��t9�U1Vu $T�@5�_�H�W�m�e��&"��'$�����cQ�;̜.c�7�n�o��-�8����xK��Q4�w�&�����Q�+�S��u��a��{�k��#��eu�O�1���n��Є	�G�H˖\n�EЫ^aP~K���z��^�^��?�	C�Nr���t1:��gТv�yx�����F��=��(Ln�Ӣ�
.<��KXP]��,R�?���$+�f^9d�0�������(N�N�me���A�)7I7�`N�'$��x z��Cb\��N�2��]=~(K�g�@��I��7AZG�hӥ>6�E��)�m�?�RwQтN������C�q()7�)�=�'��ZT��y��d��L��U�0`fLO�5���gc�?�ư��$}�A"Sgh:���6ҬE$��7�M��g���v|3�2���,�NI| ����fHC���'3�o}�aS��q�s����֒k�3>RYO&��T�v�+���r�n 0�3�U�9-\���l�@3ԦE��C��ITI)f�����y�8�2 �����<�q�fy�i���*W��[�m��N�ܓ+�P�_cK�'	����W�(�i�C��m����\��9g�W�a`P�j����k�TX�cm���mV����u��)�6�<ض��R	�[�9_�y�r��kb�X��x�n1a���N+�V�Փ�� fAL5}<p:�$�"h��B�uMH�����u(s5̆��U뢪�����փ�l��ї�AA��Go'��y����Ba�qj�N����q8*W����ye�8�t0~Eq�?^���� ������e��'8���oyfa%p� ���]D�����w+�蝭�&��r�>���ld� E@v��T�j���"�����<�Oz9��( � ?��.Lۧ&ᄥH�\�����&C�<��M�
D?�Uq ��B��'f�ւ����t���rHx{�[�+���{K�3�|s��Y��!MC�ó�i�.��r��%_�`�
��۷#b���ٚn�1�)^<�Q��m�L����F�L\ܙ�J��+��������R\�V�`�#X�%˃�{���oN)�e��=��A�GG\`C��Ԧ�
)@4��N|�ۇ����@-<��r&�\�2��E��}��U�{����iEH��s�d� �~�*a$y�Y��0'a+PZrX̯�НN���M�R~��D7*�*��n�~?�aR}Il�7��А �5��a����)zD_͔V�h'-tV ���߼��"S�q�k�{���2v��w�غ�ѵA���̀e|դ{ST���L~0��W��>kP�U���t���e�y#R�?�����et硛.�.mv���Atb�\(?*�t\@�G����v�@�j���y�i攇�~�79P?�0KQ��c*���x`p�biX�&Gc݉���5E��,�BVR逧V|p�RS,�ƹ��k�ҐH^�/b���G���Az�H§j��+C`���hH��u�l���U�I�|�j'��N�0� �}LpÚ�1��N Y�3������]�8F��Σ�r��^�4�j�7-�?��W�X"������(!���V����-�J@!�R�~�V{�s������@g*�l*�_期�Ϗ��|l�0F])j)"g6`zKk~Qx�nN��"5،����g,����I�ڜ&�Tq��_Y���P�
�cBO�{ ���or�$ݣ���5
�]敋Fc�f�o��]�'h��yMv�1f<��6c��k�����GV��0LN^��0Pϩ�UNd�Rq-2
p*��7��E�*��=���Ue�Z}U}:��`��6��~�d��Eeya�0��@���>�,^p8�gl6Rv� ���y*���G�^��St]Y�&����XN%-�D�H���ګe�����{fu�7���O�7��z�g�[4�>�	��Ym���6��̓F�:|��l��HP�tŗ�J?�r�B��� ]�����h�lriF�������Z+��'�$)J�O���a�5��^��ܰ����Lr�Up��(]��l�]T�>��I�Dq.�}��#Tc�'-���?X������}��zwz�Hy.��W6��#=�7@��.�k��0u{,�[�NΘmC�3��7�/{��*XB*�ڂ��p��H�9���&�.@�Ұ�pU-�%��njC#-�oY�,H���cD�_V\S�h����HEB?�+a"��"䌯̫-*y��8��lF�:�voh�<��gښ�Jk�P���5hO�B-�m��������w���S�C�{*�O5�Hh�$+P�Pˀ�[����j���0�v��b�)Y}������7���� �}�N���"R��Z/'������ M��Q��d�,d����)�Y����Y��Hv�7u�Nׄw�^����Y�`w+�}+���v��:���e��8�8ڏ�+��xp:��6{p�?ܦ�vZ�j��ΐ�ˏ���/�)�g�����ƛJ�d�)H_�����?�Ig�P�J?�`�`A��h�;���U=��,�Z�F[��rZ�7��%烵���ق��\\ K��E�Ά���Y�Cc`�9k�H֋FY�[�>N���e��#��gz<�-�!���1����2I�������n1*��b�%;��k��;0��h��?�����z	l��Ӎ>|ASvi���Ə����yn��n�w��mD�I��B
��/
�����D��(�W�T������s:|�7��v����>�����Dx>مX�����G�9 �}�j��t��׈�V ���褥	,0=���3'(���ŷEF��9�\��tv���F�j�j�����/�T��k+�܌�F��5�n����p�y�	�F&��3������	F;ʫP� ��n:mCr����O��Ry؇����4�S�;=����K����xibW`�M{d0���1���I�-!���}ͯ�z �f,�g�:E_D)K�?c��+�Q~�fATc�2p>��� ю�9L�E,wZ.Ib�m��É�Y�S�UU�E�B��΃0h�ʂ}QE$;��钢h�p�#�h�?���Ǚ�)�0ؓE�`o��^0W����n*�a�P,����7{EM���0k��7�lo���$�$&}E��W�b�P�U���9~S�O<Uqh|O>�T�٠J�w#6�B�J���N���a\��Dxip^�������o����� ��$7��u�FV*P��ӽ�
���G��:�c5�dX
[/o�i�l5W�ed	��Eܩ����}༮K��;ә�zT���Fxb��~;X�N-�(�W��,�.�d3/^�m-JX�o����&�[��V� �R�(g7�+����0+m$�2����f<F�ZB�귁؅��?���˽�c�?�G���2�w-��ͨ��9j�V���Jw�AŘ��]K�f
��Ot�_2צP�����	�8���轾�
��r�ҞLw?6 �g邓h��E_�'���DwsQ�y&�Y�o>1�����Mv����G���й9ɳ_�;��">�bи��F�1�v~yik������f��^q��:��o���[^�\��42�E�q[�Wނ��o"����]P���?��l�X�?�RE�;�'�_��εi���l�����~�)�!ׄ���;oSd�+sc��/������!�y@ՕQ��
��P�\��a+��.�_9c4 �q$����'�E]Ċ�}�R�TY�q1�}�*�Ȇ�ބgu;��@Єt����nr杲��߇N����<�����u1��O�ü40�A�ީ����6+v
ت�p$~��QB�����+F�L��:�Kd�ʿ��\�R�S���P�w�Cu�{>��LQ���;7d�I���p[���5��.�mjǗ��/�=��)�e/����$_4�r9?r뒳~q͗/�wq�BN�M��.ӹ��vנ��5���C5���X��Tk{�=	x��U	T�U�Y:�z��P�99��8���oo�r��)G���l�&�5N�q����>�Uk3	�~�1n������l���Tp��|b&��^T��7
�����XXb���J~X�eq܋�K{۠-�������Vc��r�7�>�=��K̖F�0,�� �b�����NS<�ǭ�MFD`^1���"�㹖S߬��3�21�Ѱc�����&".�W���6�����ZWcnN�)�Ɲ�?��>y8���@��J|�����s�Tg-Iu-G=-�H�0 ����{�s(�{�r/ZQ{Tğ���ڞjx����d�6�&�Z��M�g}ӗ�>���(n�r)���+��Yؔ���6&-I`�+��^z>�ބ�4�pr�ɉ�|e���x���VBg��Hx9~d�z��ٟ4����v��Ɛ(u|B_����&�H?�`�u\b�`@\��c~��F��k����jĠ��c��&�L�;SQ��\��A�q6��3F,�=�*�d���E���5j%_D6%`�v"���n�����H	9�+QR+�DG��C����.���0sj��e��J�|�6r��A�%1�n��?�M<k��7p�;�nh����i�'99w3��ޘ
Zj�=�3�a�_���\iw��R�a�K%��鮂����u�_f��7��U��\����"u�_?jd(sS&�~��K�� ��t�}�����ֵk���O���(�w"-�x��߼�Z�Ԋ��@�~(�q�h���[��5��a�[�1��$��T�u�5#�MT�*���O�I��ZǍs�҃XH��5ɹ
�E<K_y��:�:������T�tz�,����ES������9�F������&uA�S٦��+q�J�Oz�0P�/b*�L���h2L2&�s�-�z�d=��,���g^8 Ꙋ�i�o8��b��(:���5YQ�l�rE�OJDT�W�f���|-pb`n�e��5@y��WC�9�+0Ou
e� �'�M��B��Y�:���%��6^tμ��ێ�K��H��+0�q+��u�Tf��FV̞eh�褈�C*�|J�)_v�S���@��)��٠�=�f�]������кر��ɖJ�a�ӎ��d�ç�� qW<�'�ବ�)7�*�'f�r�B��Ki�M�)A=f�o^�&�w`	B%���U�T��%�U?Cl��Ox6���v��M�Y���ޒ2�0��1�F!a�ԃv �J�(�q�ބ�G�B����|@�j�|R-����o��<J�i:�|}�\���e�T�!�ܽ������Zb��p����a�H�����%���rR��M��S�/AC�4s�Qv�bF�L��D���dL�Ċ��ܫ�6�Q��gm{sUK�j%�@�<t7ۘ�UW>[@WGq�a�����GS������q��F�ۡ��2�٫��W��\G������8V�)@��~W:��],���IqxTl+Ǚ�ս)>��:f��$�p���� ��W2�p
�6C��w���}E�W���ȓ��'��&l,]�@͡��Y��ޖ&DFBH�2��� �g��V��$)_���C�z3���ç?��3�(�u���̔�˸|&h���m��"�Pp��$��C�3�|�A���=g�G�v�����Ct�A��[K2�j�z����2�\�*�nh�zV��?R��Ԩ�n�&0�Mpi�x6�u�v��/����rwT�>9�n�K�r,%�ć	�Yt��!�|���7z~`�m����{k� 2=+�B�����#,މ��oI�K|{�[���8��p���kR}��zI�.Q���n+ɒ�~���|m�	?/Ӯ��>+�Zl�]�t~�sˌȐB���g���H�j�~�i�%�tN�x�~'�K��S%"�%�;��g��*����`�������6�/K�nnZиAjC8�x�7RF��<��˄Q4��5ߡprn���m������C�zz���������:���U$D�`�k�*μlt���^+��"��V�u|�z�ʖ�Dj��Qj0"���,�A�ih�C�D�0㚮�t�4�Vb ��,�T�VT�sb-לJ�_H�����rK1E�\��7�>
�O+��ٸ��LtǞ��Q�M~:,j�p5F�Ŝ}OfG^��n��{����M����N	��,�(D*���Оݼ�R�Bz&�n!Y�G&�ȉ��@��Ek.*���^����H���2�����*|���I\�&WG�r�L�Mcвw���e�����s��m旳N���JU���cK�JT�H�gY)�[��Bф�,�y�a0Os,��HdUP����N8w��|R#3��yR�]�m�!�g��<�m�����OȲ�խ��p�c��/�-�˭/�(3�0�v ~�`���9In��&�b���� ������y�Q]{wf!�}p�n�7=�<T���`+�)����^�P5��B���ކ엺�p���Hm�lũ��@��JRe�ܑ-�vv�><U��b1<=�}�#����&�|�����iR%N@�_y����l���\�A�0h��^�.�HІ���n�A|#�G�zc�&��&|���5~h�@'�����~QSZsg]�lɽ� I2�P�=���Gu�'��z��*�̓�LN�J�@]�<0���^���e	�p1C��� �Hi�� �x�,<R����*��j�+D����{kФ�W�����!ۺ�~C���	��I� -Ɗ�f&6}�M:u?_�(V�p�Fi ��3�~��n�s�����63�(�/��$�x��_��Ȋ�qs[�熜8� ��/���d� ���/Õ9K�RJDJ}�
L:��	��A�#��vH��_1��?X�����GFJ�8$<���7v���UPg �ɵД�v�$<3��z�u�ä�+Ӻ���S�4tr�̕�zMP��@ɢ]V�ο�jyv���"�<Q �K"���w� ݥ�|�mZk�S@����5��9;x� �K;��28�!����G8��A�p�]t�9�Hd�n����H胱YW_b��Q�}��ǗP���s���,2���la�;bD���'��,ݿ���5���݇���i-���x��!���L�6�����)�B�L:u`遁�
s
��D̓`�p�ϥҮ��<`�1�z�C��N��,��J��:P#x��NlL~�(e�m0m�G}��֊��|B���NIåv.3-�Q%)N������F��2�Yi? ��1�U�K�8E��q����]���\�VI?�3~�Y �r�����*?RZ�ܰ��&A�k��cH��^I����n�9����X�6,,I��#\�?�[�.6��)"
;&A���y�X��}��m��A&���y1����
q��*`�=�.��-G�ӇFz�cV!D�
[�� 9���'YA��nat��� )��� 4.����b�Mp0�#��4��	ھ!{(�m��V��qEm��(j���̀쭷�l]ww{��-1]��8�cl��!�Ao�� �鼠�S��a���<�s�(��U�r�����.s�ɋ�SHK�%��w�LS�"8e;�_1<�"6�9�7{E��g�|��%1�����L����@f��6P��a�$�n?1�1�@��w����v�NT2��t��L��2�G���mό�B�:����w�7�)���J�3������)>���⳺���'k��ꀪ�Q���铱/��	YΦ�����'�hN�Н!r3��R�v�b�X�nn�&GNOu�Z�:-\E��rm��M`ô�X�V�X4S��5�mҐA_�8�)��zVzv�i�:��W�
���w�eG�9��#�
�n�(����`���Q�����6
!Hoea���X�n��IeZ�%�")� ��?���D�ސc
qjM�����:�ν���;^,�L׆u!y�ە֝��0���%^БH��ctE3�|��Ǩ���v
���;�Qo�ÿ���*|+Dϐ��lA��������j��ds�N��a���E�f@߸���P@�*��E9����"8���<1����D��2�Q��ɭ�'��q�c�'@��H�4�%�Û�3��	'pd�S�7d^L���K���AcA�a���u:6�b�X���<-lEE)������7
��k���
�J{���(T�]%^��2,�h�9:y���O�"b]E�����#i�7��sh���y� .��$`�����Ic~ȓ��d��5շӖ�[�
�|������_J����[!ZU��_���m�$��^Q�@��o��wM��}�o����х$���{�q컪x�����)������ƶBad�/��S@��Y��90o��z��Q�����k����ϳ��Hr�7�K�?��$��mE�c�%O/��r�+��`��5P2! ^D�X����+�?��W~�@o�B!�o��ښŨݚ8���G�*�yyڋ�8:���^w�u�H�4�U`�r��Ɲ{>��運1l���s3�J�]�-��}�κ���m� ��W�/h�8Hҳ�y����Ao�~�]�6s�[>ő��I���9&Kd �/%����֕X�^g=�NV]<���L.?�����։��^�1����ar":* ���lac�H����+iu���%�dzY�]*V�8��#j ��D���%���v��/wǌD�k���|,c��qϯ��[�hE��2��7���l;@h+_�r��4��da��Y��X��"ʍ��2��?�B���'ag"��-�G�D��n�lމ����j� #JL��|��me�2�"�>�d�g���^�\ ��'iJ~Q5���ƜD���<i����Q8�uY.�t��?�L�r��s��gZPgcJ�$Rr�=�m�9�K�π�)�.n�a}�u���N�4�y�uUs�1��������`����7:��I,ey���ߨf�#��o?)�ܲ�\&�嬽�ף�f�X}Q�����d���]3&9^��k�i
)(�m�k"u��Wʹ��� �����U�Ʋ,�H���o:�k��~������R�|��u�'�=�۶��q������4��
NCr!%0"q�7	I��������v��/�>rA��|�	%>EJCf7FP�C��Mpt���vx��io�K	�;wS�R��A����czWٶ�&�5�]�V.���ݐ�İ�l}�bƭ�|.��^��7O��~�s�5��=,�۸(��UZ��s�۰+�u�mdcnufq5wOTa�B��s�$AL���G�(~��Z�=�l!uC��)�jҞÞ�_-T��6��x؀jAC�J���rfD���eD91�z��E����r����D�?C7K�fx��p�,��V��Ճ�L�^�#��.���,� m� <U�,/�Erd��?::��]F��Af�,0��d��B��jobL�Kt�Jw@
c7AM��.�Yv�	���}cE*�/�5+>���h`<Ȩ�0�k��v�\���+'�F������eY�H.w�����>�&�n��M�$��?��2��=��Ê����T#"{�]�븘b���ͫȪ���lm�ߓm>�^���PKem4����k�0� �u� ��UC ����fc�P%ߴ�����e�x,��U�������b-���� �AW�(d�ˆn�H�U�5��*�ɏ�#�`�Lj�>��b����x���z�B���',��H��CRIdgG���rF<�fx�2�����*�D�a�����lJB)�4ahY҃�9G���he������'�JF_�����<[� f0/�k�v}�Heg��Q����5��fW�n�W�יZ�HΘ�� {9�pwzt�p�g@�"�?�KDڀp��}|e��~��j���Z��|�oc*�Y�T>X���#p^k	1t�>Ɂ}�$S׬ӈcN�+�S
E�{��1�7֨�w�Sd5�f&��z�y���mM���\��K��&"Vmf�3��a�*4yQ"��gH0�DX��]��8�ԋ0�ӱ���8Ӻ�
�I�^�n?إ�S�.T����IAAeO�i�8C
�Ӿj�|�9O��;_�`@ce����˂6IY�*��W:�������"��eO��G���B��t%G�})p��HZ��f>�J���<(�އ�P'��{`�E?r&Q�A�/Õ�-c@�.�,����t�i)>l�J��(�S���XXz�s~��ޯ�}�;��#`���R�gn\0��6�K�	��$���!�q����Ⱥ��d@��O��<��`���ǩ���X�P�\�X�A���;܄��̌��4kP����a��I��O� @[D����֎E&�>(D����gw@���}y7X�@��3�x�Ix�8�l>�v)��Z�"$|lL}�\��M����u;4�[A�h�S3`O1�я�8Cɋ�Wٷµ!�3�/P�Syū����>�\�J�d^�|4�R�ʜ�zuH�gKW06^���k�k'I��o5ٴ�᯿~0lV"Ev-y��ǲ�Ҩ�`��J�;hL�{�s��uE��>F"G���(��g��8�l���h��F�.�����%����kǥ��~[�{ __���T�߳S��G�r%*�cح���������/;O�\���|#z?!EħL��u!o�3�Nl��h��ܗA>�I��h�`X]D�/��]����,��xK�ܹ�.���i�zb�����IХ�-<+���X�'�.9�{Ǘq}��c-�O*��`Y�7��P�`�Bj��
=4O'6��{��>��2!׿΋�f�#�|��*�1�����𢥙S��B�#��fG��)�W;�^��$�A{�G|�������%���%��ov(h�;=?�.�H�B�b�����7%:4�� �l�&UHv%�%�����$�B=�1[�����w�"P�/��ʹ>����� vtf�LVM[��q��s4P^0F&887��UJ��6C~��>�ˈ!e�K�`�&0J1���vEɇ�U7?S��
��jd�s*At���X�u�J�jo�Z�CP|�U�� �+O�9��'��]+�j5u@ :4yDܒ��ʜ�K��cR����%s���M�%d�^V�֞���[:n1���z#9ko�2ܻ)� ���S5LDµ��G����@��!6���⸱hfV��=C��I��a�`�j�e	0O]��b�Y�@A |zvT��(�ߪiSܸ��5_��:!�3ʾ��F����l�>A4�D�iHl--;Y�F�����a�wӑ󛏡q�?�wOQ��u�G�pl_���9:F�
	1^��\�K�2E�F��9"�A��ԯ��(Lq�.�j�p����a���{��~Hx�I�^v�G9���Z�ko"��O�cc�Y@�خX۫e����kؤ��D���걡������#�Ԉӈ**]c>#1d���7��:;�����nh[��&0�U-����(ݧ���yn�;�J.��2�}��)���ي�����PT��.� '�<��E�@���5#�)��̺�*�K�_F���;�A%�wQ�ߓJG8i�(�mfT�L�M����/�A,8���!���U-����Щ�X��j��i�2a:�/)j�jI�G�߼@i�Xʜ�u�Q)��a��g��m�Ʒ�� ���.A�w��;�
d� �Ρ0�ϫ-�5�_�,�W��,�k���X+�����bϧ�4$Ŭ�<���0Fz����v�2x��X�ے�E���8���j�kMX��sc@h�>��4���S�����]e҅�`�&ċ�<������}ò��3�kH�Sź������n���S����/1С���9k�C�����g�(w���+#���A����Y����
��+��<��V��;&F�y ��c,�d����K4��Yь�M���B�݃a��䖐�M��4l0I�ٵ��M��*nn���P��MA��K���{�,n�� �7I��v���Y�YD�](�7 ]��!˅�r��nV��@���0�x	��VYQX��x�sf�h�̠�ѽ�,#G�a��s)W#m�<�dX��{d	l���~npI��z�;~S��J(�ai���6�E���9�`��b��:*����X����R�ѫ�+N{�:]h�tr��i:�g��]��q�fŕ{����{rgN�w�n���U'Z��%��:��A�����$��Ay�*:�ǱFY0�E�ux�bEU�G��~�X��[F��'6$��?�Ub.��y4��Nk�!������U�4�;��P���t1D$�q���> ���'���1zo�2�tn��`��8p����Q�"�;��tV��Uԋ�aׄ�ihѕ�u��@�&{��.]��+�;8%g �>ԲvB��0kML�P�pa	I�Cx�)|N��mGf`�01퓌N��Cb��c�h*�,�$�:٫#�/�{sxaӭ�V��!�n-�Eu� W�&����B\M F�����-Y�]�-��7D`.�s��v����[���.�{��7�m�f���5c�� M�v4�k�����
F��/Qp;��X=�
d�L���XB�1v�
����D�J$P-gUd��x�g�� �,�x�������fc��z�g��g�F"���կ^����.q�<.��� {�~��_�
v�P�S����&����$��}a�,��H��=y��� ��U7��
�.��eݺ[-�o��XN�z� >�f=ʋ�������:bGIdر�ѯ���������`�y���z���I�4���ԉƲ������� �
� l��L�ٝ����s&�8:OKyc��%G>�̶WW]lt���*T]��?l�4"di���9[��;�K�fx�yy�/N��;�z��U`H×Q���LS�-Ā����hO�`��O�f�R�hT��n�F@���O�F %"��;���k"��=�,ߧvHY� �oRq�,<��əG��`��\#M|�� #k&@u=�#�?��6i}p�������lsb���*Q�}@>�,r����5�M�N�B��u��H� �1�#�f��#�+�Z���@Xk�����K�"�7vj�;�y|d�{-s�;M�j�:��}R)t�^�������7��)����p ��[зϯ����I�(t�kܸ_b��u�\ϕR��6
�rӊ�Gb��7�+s�:
;��9o5�g8T���.` ��.0 7R6z��yZ���l�[��c�Vo ���s�l���2Y�����z8�]�m9x9���Q�\`h�+0�N