`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JyEBFm8DHF+LFfXiJXUr1tZt8HBDBj2iRfqrs0ErAkMOeEW2B43kFPJwpqHZ8Spn
I8FBdPAHr0SjaDsJ8uCQkZDak7qMRY9cEqLE0eTjDVW17UmbzAOphu6IqDu9733T
ccv+UDwT0CZWeozJHhcvvLEl0ZpfoOt5y4/5uW4tg5c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4128)
GRTUKhdFvhVRvDXu+LuKhAfWUV0z5KdRhmkroouU2fKRAFHgyvP7AQFv+lD4Sn3o
sjebk9h6ETUqVJDlhQMKTuRZ21OVOMdmlCahhxI+c7Mm3yZazh44OIa137Bl6lyF
Z+96+5f47EbpM2qKryCh3+goEu6lVzKHUTOPfReGOIh5HOrTjRXE0435bN7YCIQf
JZBK9A6lyq+T655wb5WXYh9DibpwdmYuPfcFPIIfX22zIfm+itf86qW6HAX196Xk
W5loqtJhMZDTfQJ77c9LPobSe6E72ZjNgEe+Lk32ruu2C6YPQNXN9NzfihZBirc2
E83+Akhog+Ep437UFqQomy5xy5z2tMzWm3Fk5tnY65nQ8XrjyQOq1K+yB1B5QEbw
Shy7WP6yS5sPvlx3FHidtUxWDAMLK4Xp5X+XsL8Xt/rYPqySlxCqU1MCUdREITaD
XnT6qNpGrcv6DJR2vKx3mUvG7pxY+trGRdrpljL5rDjex+zvJ0ux+Dk/fV5jrqlG
V1C5l0sNStB/uV2VXUHNl20QyuuYEaDrKSibGQtDYIRMZtTXo45l3P90FzBWTZPV
+1yOx9SugLKZ7B6XErhpGkFDUiGw+jhlnQYan0Egz0qsA0R0yRT2re4tmF99mnJa
gSS8zRpHit40bU+pudDOFGFycBlkhon+f3Cw18tMnlqwMUUHRrxe81rD/VFbbyD8
irzLENNdbMaXpF1cQ80c5UZ5Lnp4Xz3YztSn4fFslHpOUxHz1rW8rnAklls2AJbz
lP5xJM5WV1hK7WMbCiwFuRGbPIcnAQiBjOrX4qPmX4xwmmgMu94TMa21yUNJp14Z
4oDVRBiRY2E3Vm8L5KP2U3sIfryExMYz3g4R5WQGQ+Io052sjddUxa1jjcINxtWK
bFSQfMNEP5jRKkJyoR4npbaYPjCKUjcah2W1xh9I+mmiuiK8mMuSqmi74g/rcTVQ
iZkmKRYySOpZ+D6Nd39skXLcWTxVx8LbsJnbDglTVrrX0tZLZF2SuGx8ETrT8543
Q9FOmIlnxaRI6ZJ2qSmY84DE5ZROX8T8opKQZekNttbYxDxZJMa+8iYJyqZ/Xv/B
16ciZ7kfA3XZhilC6OPrGeZZOvFcyK5e1VuRx/09xCIoU60MMdBvAqeWanuqdjnB
ilF6G8a6HXJRLnjN24IGOvUXuCsjq0soE5DYcbZ5UQDHKRroQYL9PxXlhVp+bsKv
2N4ZMCP4IIOKS4npu6VM9DGp2wDKKWxwzKs4qTZ3LY3yEkSTOXsbWpF0wxVRk5n1
jUYTEMQp6SqiYqtTGqg3xrXHi1Jv2NQvLKRY74JlgKCkTbmd6926x0004XvwYfFe
q/yoZAkexDkeLJIqAUjP47H4PAGPgiV+YFvQMJAOPzco7sdJn9WyFBaza0bNEKhE
YfEjv8POcf3WjpbDHlr4eeyFu14iVlL6OjaGaiVBTZpVndA0HwjwbkF/4YCRfPEk
rJzaZTjtvzQ3anclW4TvslXfVXr46D02oOv9duLS4BbAyufvREV5meEgYuRGlCDz
9vU24ufwXBueho7+0N48q8b9rPElkQE08rx60mL8ghLn+HeriDNxV/Qk5ulKm0Bz
SgFEiexfOg5kFvJkrKsnW6X27oeUabyDWzU2dtRY6639ozBlHHItZx7Y2BofQkyR
E3khS6MoF4kO0gVkiHlXNARgqe0oWDNrsL/2bafsFv0GAUdYLd/ifAVTR2fiNO+5
XjNgfQdmp7rA/yJxZHPY4DSp30v538uIcn8h5jpo9eMp99tobeCi1Z97OMaeyo0j
gLIfaeUr366ZyiIKEhtGLiviF6lniuermleM62jFAqrPTql6wBDy5+6KXOqJRBFH
lHgcMOBp5cyFQck5fApiK+Xxhh/oFA9BW7RgQD8YeDpRXDkZ1DiFasYYOQPVawVg
J1bV56cAHESIrSSl52A3KacWxAi9mcFOb/hly32TSyDGtHRX2lv9ddVbg+3Je2F8
kOJn6mxyUVGE4EZGvARcfiufmAaLmkWRA6Phn+LyZe+N+0tdJDFPaRizdhKcaXoe
M44bobQiTFoAV7uxlX5yP3py2q5ZiN1rgEGmF7flYzyriiXzjYZUonCPF4AkX4cy
jVoUMHNP36n/42Da/hbeV9Rsl6Sebxg1K5LK8P4gAyC7tns6gNUHCvFePQFCD1jJ
9aEMLgQWlOCaDJlYL2w2pxM/Mca+TmgGVFWygBDLV2L3KkSlzqzvu2tkKEN9b85B
4tcnuRXkewnSYqMcvsW+ynab9LvC+n13dBBG3kwnvdaaJWy+RwfSOJBZu4lkwG6N
TR76GA1MDtTZwmXhLN+uCsulUN5vMgoEiYWaJT9Mm/5+FEcayBcBeudu56vRNblM
0T8cI0TJh2QO+vELyXd/xZ6XfqMYkxrYYXTtZBRNdXUOiOisF9Yd9u63JlwPHm4z
OKrFfm5X8I5yRzIz/nOyPHmV2a+FPKbqpNPNndylYwawh7QMU/J9BEs8y+IPzQKM
y3ywQP9YoTBcqWvoqoQ2fl0VYEzlniAvYO0UvCpJtR2e+/M9iRozzyxTJt5yuhtA
ZshMxfb/Vkx5HrpxTFE9KFBkZLEhF5z2J3K3LTrZuOGIRsSPOsXYHb0fGdpDFQZJ
Y1TnKBq0PjXN3oSZGIscijikgnl70djXEHamWqAOZZX1JthKn9XjgD3RyYX5l7lS
1sb75H+aCul57TPZvoRkPreayBzo9iKA665X5s2FIhVDG9Z1qfLLp4du5opRhzkb
NfKz2IPcjJNJbt2EdeQVcBdoaya4vmiZcR0f1/AtYOzqdjzERSSecqkEO/G01/ij
J956nf4pmxSB625ZnoMnZz0Oo8Zj2Hx+2XBQMIuVhSx8DBITf1hGeV6iXH7p3G3d
Eid9u9AJEZhVKiznBHkx5tlryvNRRgzbKzoySHetsPGyKRKde6tQDeUAZp/05OlU
GowWqZNZqvXJc/1HPGRe36MzMza7YOl/HUXEwVkCNjv7dI3HauDokD257gFOoC7D
WfI2HwLbjsD4nWZc16bsuDsuUkyfinV/c5v/xGM3jXHQ6uZzcburS46oaUQEJCo6
xxEDYT9oPrylJx8y96WBRoo4+e8MpOTnNmBuYcAHCt7N54thIX41wCEGilu5Z6UC
hbyPpx+JNMaGNjEWqZ8j1g7za+I91HdM8D2oKhrGFtgsRU5u5q595EtSqANcA0G1
py3Dir8O2RSZOycjXjRVCW5C2HO63hOWPZC7j1lgp5R77T/qhSh9p1eZbbTs1Md3
utoBHgzjhHiq4XUpwR/lZwfDNJCLwlDxRJvvGo0iAv7nM4DPVRCniBskEOJQ7Qks
0qLym75qPgyJ+cAtRnJzBEhHdW9vGLR1eiw7YWZdHfoxmEN7kB32aj9PzbyFcIDh
JoMru31FrfqWzTvslpWDYwGbr4qp8HAC+/yrC59744q+9j+myB/PMPwl5WgoBQLk
+FOJ/a/fuqyfJUIVMugbO9foJRakE/AcdBPT4sGdQfbz3e8HvIzWNijvl5E/PTc9
mOTzL5wEjc9v988VRiyQbOd3FEMRCNsif+gjXS73I4GTti0KBg5/xOSxj9kxvFs1
yCmyBejoPUoo0PlP/GWUmRaO5bqi0AYJjVXT5U4JLhhDZlTI1xp1XmtiKQcvfF1B
ZR2Lwy6PAjMKOu/erQJmv+Y3W1S1isk/aaNIu/KRv0XWW10CnmUH0XLQnrzO8VC7
pvFCKoBL0AEtzAmfbt8anj8shAE/bUt9EwnoE/7DbMsVqNWztRAqEusITCCsxWA4
sVBO8poaL9frnCr2BbMBewJ4zBi0h6MTfFYcnN0E9+1vmXFDP42Q+g4zavhoHMUo
PeK91UhX/CDQrQdOjg68tXh8fcPWSuumAw/jVFbOlM93EEUeZ+5ES1cwYNfIQNxR
hoS0mTSU1ZNUvjIXIWgoIS69lK1Na60I40GGNY9gzeYNzeKwHVXWtEcTrTM2xCqw
oPUH6+o34f895WPxsesOWSo99PWNSHz7SIZwNPtIB6IBhqm82QMJctK2/Dud4WSC
t+3lc1G6CAl1k729d7Ex0npdIHTFUS1Oay/RbR+Hd7c2EwKICletwA2/oeVsKhrx
CwPMK2DITL8HgoUfkW3NV7DKqS1CSvY2vLUsz80Z9yuDgLJsNqTR7NHbN4LN3Ar+
4/eh7Vgv9PdnAaWaQEVTWOFJ/xqBRb/BgXKHlLOHuBJmUTF9KswFS9+efuRE/Ge6
hU5SgRWn++A5zGR2OZbmGo/xC0q6HjA1j5G61QfAPS13mu7HcdWEeK5tDc6PNH7d
kWrKyUvlNNokB5rQTqHaYKX6SUxeDW0ZKsZRK0r1P8uvZP+sSI+kHQhw6Zyv8ls5
aFI/oEb3K203IYkdEUjyz3aWJTRkwR2h2mo97eIokEzc/Gd/ZliORAotBwG1dPua
MRaULtZGdmnvlhjxSrtoplbDeDf+/IAjbGaEb7uaLV7UgH6s3NayWS5hCqO+3+2C
qBNXOcoNkr849bnNpsjRzwnWVEDPfVKOoUI7PWoj/na6F+V2TyKceTecZIUwBLK5
ZMpbwa42qvuUgycGsEao+9CNb6x7IkjOTdPY/kLTtMA4KSHrpKNo+B+JuxZd1wq+
PIm5c5PP4nwgqgZlrvPeySQr5SmgweCs4l/nEfJq0XbCgyNCx3RQc5oGyXF2ITxv
f2FpTd+1cXcpYEwo/qMv36CEDBCDaHEqN7CGg2QeRHPXXaa5GBRapFyCOMp6wOg+
dTD33Gy4b9KE/XK5f3NiuvaXMl17EehfWF7bQpcu6riq7/FdtHfLL6c4+UXEu+pu
Vd7SHXh0SNIH1EyF3ofJWIF3cQg9cf1oqmXpzMBGimKmsO9RAdQ4QHViNSHtJNi2
vxkScPV32VYNL7Hx+x/kw+JzrrO/+mU9jnOktYpBCi8XRl3K/UVo7L5oW8mlhOz2
POHoDCpA/Ai/6SmhtTfmThF2Bmc6t0FIsZZ+orLDXaOCpsXdtR7TNdoxiZpMslpK
s9kKmEK+ZjbRWiHnwXaLSG6CNaTxlU24GvnAkg33JfM3Uom+qnV8Iwda7gNHiRXe
hQG1lQntNAGopouC8jq8cNKpEAUR0buJfp36YCHvCRXYtuMycuq2Ls3Ir+wyI2Zg
6KE/7INA9OlL3Bigr7GD1EwNteVyz4xZp6LfEXhgyI3boYHSciKweIxGoH0e8fwq
Am+vv/LaUQthRwdQc0xcSb5lxEIVKSfc6t22y2kJVYkZMm6KjoCtzgDPirU3DCWH
8/S4X6yH5rbQ4jX6PjYN6bbYYT1F3QvsDEvHMnF42bCFadJcb6IwFp87fxQUQLsc
IzYCvXngp1dOb5ddl+ykQ+3ISNQIhLesko0K9pIEzxgTTCk1mwqthM7TStJe3EVX
7c7HV8KQf8m9Fp+vrln3hJJQpi2NCql3QBn7pB9JpCdGfEWdLp6n8MwekMKz6vbL
/0Nt2C22/yfbJcbWB2cryy5dTBR3SHNS1/AdOLXHvgZP2pDZOX8VQBAaq/NaqIkU
`pragma protect end_protected
