-- niosvprocessor.vhd

-- Generated using ACDS version 23.1 991

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosvprocessor is
	port (
		clk_clk : in std_logic := '0'  -- clk.clk
	);
end entity niosvprocessor;

architecture rtl of niosvprocessor is
	component niosvprocessor_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component niosvprocessor_jtag;

	component niosvprocessor_niosvprocessor is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset_reset                  : in  std_logic                     := 'X';             -- reset
			platform_irq_rx_irq          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			instruction_manager_awaddr   : out std_logic_vector(31 downto 0);                    -- awaddr
			instruction_manager_awsize   : out std_logic_vector(2 downto 0);                     -- awsize
			instruction_manager_awlen    : out std_logic_vector(7 downto 0);                     -- awlen
			instruction_manager_awprot   : out std_logic_vector(2 downto 0);                     -- awprot
			instruction_manager_awvalid  : out std_logic;                                        -- awvalid
			instruction_manager_awburst  : out std_logic_vector(1 downto 0);                     -- awburst
			instruction_manager_awready  : in  std_logic                     := 'X';             -- awready
			instruction_manager_wdata    : out std_logic_vector(31 downto 0);                    -- wdata
			instruction_manager_wstrb    : out std_logic_vector(3 downto 0);                     -- wstrb
			instruction_manager_wlast    : out std_logic;                                        -- wlast
			instruction_manager_wvalid   : out std_logic;                                        -- wvalid
			instruction_manager_wready   : in  std_logic                     := 'X';             -- wready
			instruction_manager_bresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			instruction_manager_bvalid   : in  std_logic                     := 'X';             -- bvalid
			instruction_manager_bready   : out std_logic;                                        -- bready
			instruction_manager_araddr   : out std_logic_vector(31 downto 0);                    -- araddr
			instruction_manager_arsize   : out std_logic_vector(2 downto 0);                     -- arsize
			instruction_manager_arlen    : out std_logic_vector(7 downto 0);                     -- arlen
			instruction_manager_arprot   : out std_logic_vector(2 downto 0);                     -- arprot
			instruction_manager_arvalid  : out std_logic;                                        -- arvalid
			instruction_manager_arburst  : out std_logic_vector(1 downto 0);                     -- arburst
			instruction_manager_arready  : in  std_logic                     := 'X';             -- arready
			instruction_manager_rdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			instruction_manager_rresp    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			instruction_manager_rvalid   : in  std_logic                     := 'X';             -- rvalid
			instruction_manager_rready   : out std_logic;                                        -- rready
			instruction_manager_rlast    : in  std_logic                     := 'X';             -- rlast
			data_manager_awaddr          : out std_logic_vector(31 downto 0);                    -- awaddr
			data_manager_awsize          : out std_logic_vector(2 downto 0);                     -- awsize
			data_manager_awlen           : out std_logic_vector(7 downto 0);                     -- awlen
			data_manager_awprot          : out std_logic_vector(2 downto 0);                     -- awprot
			data_manager_awvalid         : out std_logic;                                        -- awvalid
			data_manager_awready         : in  std_logic                     := 'X';             -- awready
			data_manager_wdata           : out std_logic_vector(31 downto 0);                    -- wdata
			data_manager_wstrb           : out std_logic_vector(3 downto 0);                     -- wstrb
			data_manager_wlast           : out std_logic;                                        -- wlast
			data_manager_wvalid          : out std_logic;                                        -- wvalid
			data_manager_wready          : in  std_logic                     := 'X';             -- wready
			data_manager_bresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			data_manager_bvalid          : in  std_logic                     := 'X';             -- bvalid
			data_manager_bready          : out std_logic;                                        -- bready
			data_manager_araddr          : out std_logic_vector(31 downto 0);                    -- araddr
			data_manager_arsize          : out std_logic_vector(2 downto 0);                     -- arsize
			data_manager_arlen           : out std_logic_vector(7 downto 0);                     -- arlen
			data_manager_arprot          : out std_logic_vector(2 downto 0);                     -- arprot
			data_manager_arvalid         : out std_logic;                                        -- arvalid
			data_manager_arready         : in  std_logic                     := 'X';             -- arready
			data_manager_rdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			data_manager_rresp           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			data_manager_rvalid          : in  std_logic                     := 'X';             -- rvalid
			data_manager_rlast           : in  std_logic                     := 'X';             -- rlast
			data_manager_rready          : out std_logic;                                        -- rready
			ndm_reset_in_reset           : in  std_logic                     := 'X';             -- reset
			timer_sw_agent_write         : in  std_logic                     := 'X';             -- write
			timer_sw_agent_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			timer_sw_agent_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			timer_sw_agent_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			timer_sw_agent_read          : in  std_logic                     := 'X';             -- read
			timer_sw_agent_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			timer_sw_agent_readdatavalid : out std_logic;                                        -- readdatavalid
			timer_sw_agent_waitrequest   : out std_logic;                                        -- waitrequest
			dm_agent_write               : in  std_logic                     := 'X';             -- write
			dm_agent_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dm_agent_address             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			dm_agent_read                : in  std_logic                     := 'X';             -- read
			dm_agent_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			dm_agent_readdatavalid       : out std_logic;                                        -- readdatavalid
			dm_agent_waitrequest         : out std_logic;                                        -- waitrequest
			dbg_reset_out_reset          : out std_logic                                         -- reset
		);
	end component niosvprocessor_niosvprocessor;

	component niosvprocessor_sram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component niosvprocessor_sram;

	component niosvprocessor_mm_interconnect_0 is
		port (
			niosvprocessor_data_manager_awaddr               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			niosvprocessor_data_manager_awlen                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			niosvprocessor_data_manager_awsize               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			niosvprocessor_data_manager_awprot               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			niosvprocessor_data_manager_awvalid              : in  std_logic                     := 'X';             -- awvalid
			niosvprocessor_data_manager_awready              : out std_logic;                                        -- awready
			niosvprocessor_data_manager_wdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			niosvprocessor_data_manager_wstrb                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			niosvprocessor_data_manager_wlast                : in  std_logic                     := 'X';             -- wlast
			niosvprocessor_data_manager_wvalid               : in  std_logic                     := 'X';             -- wvalid
			niosvprocessor_data_manager_wready               : out std_logic;                                        -- wready
			niosvprocessor_data_manager_bresp                : out std_logic_vector(1 downto 0);                     -- bresp
			niosvprocessor_data_manager_bvalid               : out std_logic;                                        -- bvalid
			niosvprocessor_data_manager_bready               : in  std_logic                     := 'X';             -- bready
			niosvprocessor_data_manager_araddr               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			niosvprocessor_data_manager_arlen                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			niosvprocessor_data_manager_arsize               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			niosvprocessor_data_manager_arprot               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			niosvprocessor_data_manager_arvalid              : in  std_logic                     := 'X';             -- arvalid
			niosvprocessor_data_manager_arready              : out std_logic;                                        -- arready
			niosvprocessor_data_manager_rdata                : out std_logic_vector(31 downto 0);                    -- rdata
			niosvprocessor_data_manager_rresp                : out std_logic_vector(1 downto 0);                     -- rresp
			niosvprocessor_data_manager_rlast                : out std_logic;                                        -- rlast
			niosvprocessor_data_manager_rvalid               : out std_logic;                                        -- rvalid
			niosvprocessor_data_manager_rready               : in  std_logic                     := 'X';             -- rready
			niosvprocessor_instruction_manager_awaddr        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			niosvprocessor_instruction_manager_awlen         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- awlen
			niosvprocessor_instruction_manager_awsize        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			niosvprocessor_instruction_manager_awburst       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			niosvprocessor_instruction_manager_awprot        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			niosvprocessor_instruction_manager_awvalid       : in  std_logic                     := 'X';             -- awvalid
			niosvprocessor_instruction_manager_awready       : out std_logic;                                        -- awready
			niosvprocessor_instruction_manager_wdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			niosvprocessor_instruction_manager_wstrb         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			niosvprocessor_instruction_manager_wlast         : in  std_logic                     := 'X';             -- wlast
			niosvprocessor_instruction_manager_wvalid        : in  std_logic                     := 'X';             -- wvalid
			niosvprocessor_instruction_manager_wready        : out std_logic;                                        -- wready
			niosvprocessor_instruction_manager_bresp         : out std_logic_vector(1 downto 0);                     -- bresp
			niosvprocessor_instruction_manager_bvalid        : out std_logic;                                        -- bvalid
			niosvprocessor_instruction_manager_bready        : in  std_logic                     := 'X';             -- bready
			niosvprocessor_instruction_manager_araddr        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			niosvprocessor_instruction_manager_arlen         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- arlen
			niosvprocessor_instruction_manager_arsize        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			niosvprocessor_instruction_manager_arburst       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			niosvprocessor_instruction_manager_arprot        : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			niosvprocessor_instruction_manager_arvalid       : in  std_logic                     := 'X';             -- arvalid
			niosvprocessor_instruction_manager_arready       : out std_logic;                                        -- arready
			niosvprocessor_instruction_manager_rdata         : out std_logic_vector(31 downto 0);                    -- rdata
			niosvprocessor_instruction_manager_rresp         : out std_logic_vector(1 downto 0);                     -- rresp
			niosvprocessor_instruction_manager_rlast         : out std_logic;                                        -- rlast
			niosvprocessor_instruction_manager_rvalid        : out std_logic;                                        -- rvalid
			niosvprocessor_instruction_manager_rready        : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			niosvprocessor_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			niosvprocessor_dm_agent_address                  : out std_logic_vector(15 downto 0);                    -- address
			niosvprocessor_dm_agent_write                    : out std_logic;                                        -- write
			niosvprocessor_dm_agent_read                     : out std_logic;                                        -- read
			niosvprocessor_dm_agent_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			niosvprocessor_dm_agent_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			niosvprocessor_dm_agent_readdatavalid            : in  std_logic                     := 'X';             -- readdatavalid
			niosvprocessor_dm_agent_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			niosvprocessor_timer_sw_agent_address            : out std_logic_vector(5 downto 0);                     -- address
			niosvprocessor_timer_sw_agent_write              : out std_logic;                                        -- write
			niosvprocessor_timer_sw_agent_read               : out std_logic;                                        -- read
			niosvprocessor_timer_sw_agent_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			niosvprocessor_timer_sw_agent_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			niosvprocessor_timer_sw_agent_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			niosvprocessor_timer_sw_agent_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			niosvprocessor_timer_sw_agent_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			sram_s1_address                                  : out std_logic_vector(16 downto 0);                    -- address
			sram_s1_write                                    : out std_logic;                                        -- write
			sram_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sram_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			sram_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			sram_s1_chipselect                               : out std_logic;                                        -- chipselect
			sram_s1_clken                                    : out std_logic                                         -- clken
		);
	end component niosvprocessor_mm_interconnect_0;

	component niosvprocessor_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component niosvprocessor_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal niosvprocessor_dbg_reset_out_reset                            : std_logic;                     -- niosvprocessor:dbg_reset_out_reset -> rst_controller:reset_in0
	signal niosvprocessor_data_manager_arlen                             : std_logic_vector(7 downto 0);  -- niosvprocessor:data_manager_arlen -> mm_interconnect_0:niosvprocessor_data_manager_arlen
	signal niosvprocessor_data_manager_wstrb                             : std_logic_vector(3 downto 0);  -- niosvprocessor:data_manager_wstrb -> mm_interconnect_0:niosvprocessor_data_manager_wstrb
	signal niosvprocessor_data_manager_wready                            : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_wready -> niosvprocessor:data_manager_wready
	signal niosvprocessor_data_manager_rready                            : std_logic;                     -- niosvprocessor:data_manager_rready -> mm_interconnect_0:niosvprocessor_data_manager_rready
	signal niosvprocessor_data_manager_awlen                             : std_logic_vector(7 downto 0);  -- niosvprocessor:data_manager_awlen -> mm_interconnect_0:niosvprocessor_data_manager_awlen
	signal niosvprocessor_data_manager_wvalid                            : std_logic;                     -- niosvprocessor:data_manager_wvalid -> mm_interconnect_0:niosvprocessor_data_manager_wvalid
	signal niosvprocessor_data_manager_araddr                            : std_logic_vector(31 downto 0); -- niosvprocessor:data_manager_araddr -> mm_interconnect_0:niosvprocessor_data_manager_araddr
	signal niosvprocessor_data_manager_arprot                            : std_logic_vector(2 downto 0);  -- niosvprocessor:data_manager_arprot -> mm_interconnect_0:niosvprocessor_data_manager_arprot
	signal niosvprocessor_data_manager_awprot                            : std_logic_vector(2 downto 0);  -- niosvprocessor:data_manager_awprot -> mm_interconnect_0:niosvprocessor_data_manager_awprot
	signal niosvprocessor_data_manager_wdata                             : std_logic_vector(31 downto 0); -- niosvprocessor:data_manager_wdata -> mm_interconnect_0:niosvprocessor_data_manager_wdata
	signal niosvprocessor_data_manager_arvalid                           : std_logic;                     -- niosvprocessor:data_manager_arvalid -> mm_interconnect_0:niosvprocessor_data_manager_arvalid
	signal niosvprocessor_data_manager_awaddr                            : std_logic_vector(31 downto 0); -- niosvprocessor:data_manager_awaddr -> mm_interconnect_0:niosvprocessor_data_manager_awaddr
	signal niosvprocessor_data_manager_bresp                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosvprocessor_data_manager_bresp -> niosvprocessor:data_manager_bresp
	signal niosvprocessor_data_manager_arready                           : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_arready -> niosvprocessor:data_manager_arready
	signal niosvprocessor_data_manager_rdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosvprocessor_data_manager_rdata -> niosvprocessor:data_manager_rdata
	signal niosvprocessor_data_manager_awready                           : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_awready -> niosvprocessor:data_manager_awready
	signal niosvprocessor_data_manager_arsize                            : std_logic_vector(2 downto 0);  -- niosvprocessor:data_manager_arsize -> mm_interconnect_0:niosvprocessor_data_manager_arsize
	signal niosvprocessor_data_manager_bready                            : std_logic;                     -- niosvprocessor:data_manager_bready -> mm_interconnect_0:niosvprocessor_data_manager_bready
	signal niosvprocessor_data_manager_rlast                             : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_rlast -> niosvprocessor:data_manager_rlast
	signal niosvprocessor_data_manager_wlast                             : std_logic;                     -- niosvprocessor:data_manager_wlast -> mm_interconnect_0:niosvprocessor_data_manager_wlast
	signal niosvprocessor_data_manager_rresp                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosvprocessor_data_manager_rresp -> niosvprocessor:data_manager_rresp
	signal niosvprocessor_data_manager_bvalid                            : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_bvalid -> niosvprocessor:data_manager_bvalid
	signal niosvprocessor_data_manager_awsize                            : std_logic_vector(2 downto 0);  -- niosvprocessor:data_manager_awsize -> mm_interconnect_0:niosvprocessor_data_manager_awsize
	signal niosvprocessor_data_manager_awvalid                           : std_logic;                     -- niosvprocessor:data_manager_awvalid -> mm_interconnect_0:niosvprocessor_data_manager_awvalid
	signal niosvprocessor_data_manager_rvalid                            : std_logic;                     -- mm_interconnect_0:niosvprocessor_data_manager_rvalid -> niosvprocessor:data_manager_rvalid
	signal niosvprocessor_instruction_manager_awburst                    : std_logic_vector(1 downto 0);  -- niosvprocessor:instruction_manager_awburst -> mm_interconnect_0:niosvprocessor_instruction_manager_awburst
	signal niosvprocessor_instruction_manager_arlen                      : std_logic_vector(7 downto 0);  -- niosvprocessor:instruction_manager_arlen -> mm_interconnect_0:niosvprocessor_instruction_manager_arlen
	signal niosvprocessor_instruction_manager_wstrb                      : std_logic_vector(3 downto 0);  -- niosvprocessor:instruction_manager_wstrb -> mm_interconnect_0:niosvprocessor_instruction_manager_wstrb
	signal niosvprocessor_instruction_manager_wready                     : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_wready -> niosvprocessor:instruction_manager_wready
	signal niosvprocessor_instruction_manager_rready                     : std_logic;                     -- niosvprocessor:instruction_manager_rready -> mm_interconnect_0:niosvprocessor_instruction_manager_rready
	signal niosvprocessor_instruction_manager_awlen                      : std_logic_vector(7 downto 0);  -- niosvprocessor:instruction_manager_awlen -> mm_interconnect_0:niosvprocessor_instruction_manager_awlen
	signal niosvprocessor_instruction_manager_wvalid                     : std_logic;                     -- niosvprocessor:instruction_manager_wvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_wvalid
	signal niosvprocessor_instruction_manager_araddr                     : std_logic_vector(31 downto 0); -- niosvprocessor:instruction_manager_araddr -> mm_interconnect_0:niosvprocessor_instruction_manager_araddr
	signal niosvprocessor_instruction_manager_arprot                     : std_logic_vector(2 downto 0);  -- niosvprocessor:instruction_manager_arprot -> mm_interconnect_0:niosvprocessor_instruction_manager_arprot
	signal niosvprocessor_instruction_manager_awprot                     : std_logic_vector(2 downto 0);  -- niosvprocessor:instruction_manager_awprot -> mm_interconnect_0:niosvprocessor_instruction_manager_awprot
	signal niosvprocessor_instruction_manager_wdata                      : std_logic_vector(31 downto 0); -- niosvprocessor:instruction_manager_wdata -> mm_interconnect_0:niosvprocessor_instruction_manager_wdata
	signal niosvprocessor_instruction_manager_arvalid                    : std_logic;                     -- niosvprocessor:instruction_manager_arvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_arvalid
	signal niosvprocessor_instruction_manager_awaddr                     : std_logic_vector(31 downto 0); -- niosvprocessor:instruction_manager_awaddr -> mm_interconnect_0:niosvprocessor_instruction_manager_awaddr
	signal niosvprocessor_instruction_manager_bresp                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosvprocessor_instruction_manager_bresp -> niosvprocessor:instruction_manager_bresp
	signal niosvprocessor_instruction_manager_arready                    : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_arready -> niosvprocessor:instruction_manager_arready
	signal niosvprocessor_instruction_manager_rdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosvprocessor_instruction_manager_rdata -> niosvprocessor:instruction_manager_rdata
	signal niosvprocessor_instruction_manager_awready                    : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_awready -> niosvprocessor:instruction_manager_awready
	signal niosvprocessor_instruction_manager_arburst                    : std_logic_vector(1 downto 0);  -- niosvprocessor:instruction_manager_arburst -> mm_interconnect_0:niosvprocessor_instruction_manager_arburst
	signal niosvprocessor_instruction_manager_arsize                     : std_logic_vector(2 downto 0);  -- niosvprocessor:instruction_manager_arsize -> mm_interconnect_0:niosvprocessor_instruction_manager_arsize
	signal niosvprocessor_instruction_manager_bready                     : std_logic;                     -- niosvprocessor:instruction_manager_bready -> mm_interconnect_0:niosvprocessor_instruction_manager_bready
	signal niosvprocessor_instruction_manager_rlast                      : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_rlast -> niosvprocessor:instruction_manager_rlast
	signal niosvprocessor_instruction_manager_wlast                      : std_logic;                     -- niosvprocessor:instruction_manager_wlast -> mm_interconnect_0:niosvprocessor_instruction_manager_wlast
	signal niosvprocessor_instruction_manager_rresp                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:niosvprocessor_instruction_manager_rresp -> niosvprocessor:instruction_manager_rresp
	signal niosvprocessor_instruction_manager_bvalid                     : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_bvalid -> niosvprocessor:instruction_manager_bvalid
	signal niosvprocessor_instruction_manager_awsize                     : std_logic_vector(2 downto 0);  -- niosvprocessor:instruction_manager_awsize -> mm_interconnect_0:niosvprocessor_instruction_manager_awsize
	signal niosvprocessor_instruction_manager_awvalid                    : std_logic;                     -- niosvprocessor:instruction_manager_awvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_awvalid
	signal niosvprocessor_instruction_manager_rvalid                     : std_logic;                     -- mm_interconnect_0:niosvprocessor_instruction_manager_rvalid -> niosvprocessor:instruction_manager_rvalid
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest          : std_logic;                     -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal mm_interconnect_0_niosvprocessor_dm_agent_readdata            : std_logic_vector(31 downto 0); -- niosvprocessor:dm_agent_readdata -> mm_interconnect_0:niosvprocessor_dm_agent_readdata
	signal mm_interconnect_0_niosvprocessor_dm_agent_waitrequest         : std_logic;                     -- niosvprocessor:dm_agent_waitrequest -> mm_interconnect_0:niosvprocessor_dm_agent_waitrequest
	signal mm_interconnect_0_niosvprocessor_dm_agent_address             : std_logic_vector(15 downto 0); -- mm_interconnect_0:niosvprocessor_dm_agent_address -> niosvprocessor:dm_agent_address
	signal mm_interconnect_0_niosvprocessor_dm_agent_read                : std_logic;                     -- mm_interconnect_0:niosvprocessor_dm_agent_read -> niosvprocessor:dm_agent_read
	signal mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid       : std_logic;                     -- niosvprocessor:dm_agent_readdatavalid -> mm_interconnect_0:niosvprocessor_dm_agent_readdatavalid
	signal mm_interconnect_0_niosvprocessor_dm_agent_write               : std_logic;                     -- mm_interconnect_0:niosvprocessor_dm_agent_write -> niosvprocessor:dm_agent_write
	signal mm_interconnect_0_niosvprocessor_dm_agent_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosvprocessor_dm_agent_writedata -> niosvprocessor:dm_agent_writedata
	signal mm_interconnect_0_sram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:sram_s1_chipselect -> sram:chipselect
	signal mm_interconnect_0_sram_s1_readdata                            : std_logic_vector(31 downto 0); -- sram:readdata -> mm_interconnect_0:sram_s1_readdata
	signal mm_interconnect_0_sram_s1_address                             : std_logic_vector(16 downto 0); -- mm_interconnect_0:sram_s1_address -> sram:address
	signal mm_interconnect_0_sram_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sram_s1_byteenable -> sram:byteenable
	signal mm_interconnect_0_sram_s1_write                               : std_logic;                     -- mm_interconnect_0:sram_s1_write -> sram:write
	signal mm_interconnect_0_sram_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:sram_s1_writedata -> sram:writedata
	signal mm_interconnect_0_sram_s1_clken                               : std_logic;                     -- mm_interconnect_0:sram_s1_clken -> sram:clken
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata      : std_logic_vector(31 downto 0); -- niosvprocessor:timer_sw_agent_readdata -> mm_interconnect_0:niosvprocessor_timer_sw_agent_readdata
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest   : std_logic;                     -- niosvprocessor:timer_sw_agent_waitrequest -> mm_interconnect_0:niosvprocessor_timer_sw_agent_waitrequest
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_address       : std_logic_vector(5 downto 0);  -- mm_interconnect_0:niosvprocessor_timer_sw_agent_address -> niosvprocessor:timer_sw_agent_address
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_read          : std_logic;                     -- mm_interconnect_0:niosvprocessor_timer_sw_agent_read -> niosvprocessor:timer_sw_agent_read
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:niosvprocessor_timer_sw_agent_byteenable -> niosvprocessor:timer_sw_agent_byteenable
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid : std_logic;                     -- niosvprocessor:timer_sw_agent_readdatavalid -> mm_interconnect_0:niosvprocessor_timer_sw_agent_readdatavalid
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_write         : std_logic;                     -- mm_interconnect_0:niosvprocessor_timer_sw_agent_write -> niosvprocessor:timer_sw_agent_write
	signal mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:niosvprocessor_timer_sw_agent_writedata -> niosvprocessor:timer_sw_agent_writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal niosvprocessor_platform_irq_rx_irq                            : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> niosvprocessor:platform_irq_rx_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:niosvprocessor_reset_reset_bridge_in_reset_reset, niosvprocessor:ndm_reset_in_reset, niosvprocessor:reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sram:reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [rst_translator:reset_req_in, sram:reset_req]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> jtag:rst_n

begin

	jtag : component niosvprocessor_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	niosvprocessor : component niosvprocessor_niosvprocessor
		port map (
			clk                          => clk_clk,                                                       --                 clk.clk
			reset_reset                  => rst_controller_reset_out_reset,                                --               reset.reset
			platform_irq_rx_irq          => niosvprocessor_platform_irq_rx_irq,                            --     platform_irq_rx.irq
			instruction_manager_awaddr   => niosvprocessor_instruction_manager_awaddr,                     -- instruction_manager.awaddr
			instruction_manager_awsize   => niosvprocessor_instruction_manager_awsize,                     --                    .awsize
			instruction_manager_awlen    => niosvprocessor_instruction_manager_awlen,                      --                    .awlen
			instruction_manager_awprot   => niosvprocessor_instruction_manager_awprot,                     --                    .awprot
			instruction_manager_awvalid  => niosvprocessor_instruction_manager_awvalid,                    --                    .awvalid
			instruction_manager_awburst  => niosvprocessor_instruction_manager_awburst,                    --                    .awburst
			instruction_manager_awready  => niosvprocessor_instruction_manager_awready,                    --                    .awready
			instruction_manager_wdata    => niosvprocessor_instruction_manager_wdata,                      --                    .wdata
			instruction_manager_wstrb    => niosvprocessor_instruction_manager_wstrb,                      --                    .wstrb
			instruction_manager_wlast    => niosvprocessor_instruction_manager_wlast,                      --                    .wlast
			instruction_manager_wvalid   => niosvprocessor_instruction_manager_wvalid,                     --                    .wvalid
			instruction_manager_wready   => niosvprocessor_instruction_manager_wready,                     --                    .wready
			instruction_manager_bresp    => niosvprocessor_instruction_manager_bresp,                      --                    .bresp
			instruction_manager_bvalid   => niosvprocessor_instruction_manager_bvalid,                     --                    .bvalid
			instruction_manager_bready   => niosvprocessor_instruction_manager_bready,                     --                    .bready
			instruction_manager_araddr   => niosvprocessor_instruction_manager_araddr,                     --                    .araddr
			instruction_manager_arsize   => niosvprocessor_instruction_manager_arsize,                     --                    .arsize
			instruction_manager_arlen    => niosvprocessor_instruction_manager_arlen,                      --                    .arlen
			instruction_manager_arprot   => niosvprocessor_instruction_manager_arprot,                     --                    .arprot
			instruction_manager_arvalid  => niosvprocessor_instruction_manager_arvalid,                    --                    .arvalid
			instruction_manager_arburst  => niosvprocessor_instruction_manager_arburst,                    --                    .arburst
			instruction_manager_arready  => niosvprocessor_instruction_manager_arready,                    --                    .arready
			instruction_manager_rdata    => niosvprocessor_instruction_manager_rdata,                      --                    .rdata
			instruction_manager_rresp    => niosvprocessor_instruction_manager_rresp,                      --                    .rresp
			instruction_manager_rvalid   => niosvprocessor_instruction_manager_rvalid,                     --                    .rvalid
			instruction_manager_rready   => niosvprocessor_instruction_manager_rready,                     --                    .rready
			instruction_manager_rlast    => niosvprocessor_instruction_manager_rlast,                      --                    .rlast
			data_manager_awaddr          => niosvprocessor_data_manager_awaddr,                            --        data_manager.awaddr
			data_manager_awsize          => niosvprocessor_data_manager_awsize,                            --                    .awsize
			data_manager_awlen           => niosvprocessor_data_manager_awlen,                             --                    .awlen
			data_manager_awprot          => niosvprocessor_data_manager_awprot,                            --                    .awprot
			data_manager_awvalid         => niosvprocessor_data_manager_awvalid,                           --                    .awvalid
			data_manager_awready         => niosvprocessor_data_manager_awready,                           --                    .awready
			data_manager_wdata           => niosvprocessor_data_manager_wdata,                             --                    .wdata
			data_manager_wstrb           => niosvprocessor_data_manager_wstrb,                             --                    .wstrb
			data_manager_wlast           => niosvprocessor_data_manager_wlast,                             --                    .wlast
			data_manager_wvalid          => niosvprocessor_data_manager_wvalid,                            --                    .wvalid
			data_manager_wready          => niosvprocessor_data_manager_wready,                            --                    .wready
			data_manager_bresp           => niosvprocessor_data_manager_bresp,                             --                    .bresp
			data_manager_bvalid          => niosvprocessor_data_manager_bvalid,                            --                    .bvalid
			data_manager_bready          => niosvprocessor_data_manager_bready,                            --                    .bready
			data_manager_araddr          => niosvprocessor_data_manager_araddr,                            --                    .araddr
			data_manager_arsize          => niosvprocessor_data_manager_arsize,                            --                    .arsize
			data_manager_arlen           => niosvprocessor_data_manager_arlen,                             --                    .arlen
			data_manager_arprot          => niosvprocessor_data_manager_arprot,                            --                    .arprot
			data_manager_arvalid         => niosvprocessor_data_manager_arvalid,                           --                    .arvalid
			data_manager_arready         => niosvprocessor_data_manager_arready,                           --                    .arready
			data_manager_rdata           => niosvprocessor_data_manager_rdata,                             --                    .rdata
			data_manager_rresp           => niosvprocessor_data_manager_rresp,                             --                    .rresp
			data_manager_rvalid          => niosvprocessor_data_manager_rvalid,                            --                    .rvalid
			data_manager_rlast           => niosvprocessor_data_manager_rlast,                             --                    .rlast
			data_manager_rready          => niosvprocessor_data_manager_rready,                            --                    .rready
			ndm_reset_in_reset           => rst_controller_reset_out_reset,                                --        ndm_reset_in.reset
			timer_sw_agent_write         => mm_interconnect_0_niosvprocessor_timer_sw_agent_write,         --      timer_sw_agent.write
			timer_sw_agent_writedata     => mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata,     --                    .writedata
			timer_sw_agent_byteenable    => mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable,    --                    .byteenable
			timer_sw_agent_address       => mm_interconnect_0_niosvprocessor_timer_sw_agent_address,       --                    .address
			timer_sw_agent_read          => mm_interconnect_0_niosvprocessor_timer_sw_agent_read,          --                    .read
			timer_sw_agent_readdata      => mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata,      --                    .readdata
			timer_sw_agent_readdatavalid => mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid, --                    .readdatavalid
			timer_sw_agent_waitrequest   => mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest,   --                    .waitrequest
			dm_agent_write               => mm_interconnect_0_niosvprocessor_dm_agent_write,               --            dm_agent.write
			dm_agent_writedata           => mm_interconnect_0_niosvprocessor_dm_agent_writedata,           --                    .writedata
			dm_agent_address             => mm_interconnect_0_niosvprocessor_dm_agent_address,             --                    .address
			dm_agent_read                => mm_interconnect_0_niosvprocessor_dm_agent_read,                --                    .read
			dm_agent_readdata            => mm_interconnect_0_niosvprocessor_dm_agent_readdata,            --                    .readdata
			dm_agent_readdatavalid       => mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid,       --                    .readdatavalid
			dm_agent_waitrequest         => mm_interconnect_0_niosvprocessor_dm_agent_waitrequest,         --                    .waitrequest
			dbg_reset_out_reset          => niosvprocessor_dbg_reset_out_reset                             --       dbg_reset_out.reset
		);

	sram : component niosvprocessor_sram
		port map (
			clk        => clk_clk,                              --   clk1.clk
			address    => mm_interconnect_0_sram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_sram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_sram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_sram_s1_write,      --       .write
			readdata   => mm_interconnect_0_sram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_sram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_sram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze     => '0'                                   -- (terminated)
		);

	mm_interconnect_0 : component niosvprocessor_mm_interconnect_0
		port map (
			niosvprocessor_data_manager_awaddr               => niosvprocessor_data_manager_awaddr,                            --                niosvprocessor_data_manager.awaddr
			niosvprocessor_data_manager_awlen                => niosvprocessor_data_manager_awlen,                             --                                           .awlen
			niosvprocessor_data_manager_awsize               => niosvprocessor_data_manager_awsize,                            --                                           .awsize
			niosvprocessor_data_manager_awprot               => niosvprocessor_data_manager_awprot,                            --                                           .awprot
			niosvprocessor_data_manager_awvalid              => niosvprocessor_data_manager_awvalid,                           --                                           .awvalid
			niosvprocessor_data_manager_awready              => niosvprocessor_data_manager_awready,                           --                                           .awready
			niosvprocessor_data_manager_wdata                => niosvprocessor_data_manager_wdata,                             --                                           .wdata
			niosvprocessor_data_manager_wstrb                => niosvprocessor_data_manager_wstrb,                             --                                           .wstrb
			niosvprocessor_data_manager_wlast                => niosvprocessor_data_manager_wlast,                             --                                           .wlast
			niosvprocessor_data_manager_wvalid               => niosvprocessor_data_manager_wvalid,                            --                                           .wvalid
			niosvprocessor_data_manager_wready               => niosvprocessor_data_manager_wready,                            --                                           .wready
			niosvprocessor_data_manager_bresp                => niosvprocessor_data_manager_bresp,                             --                                           .bresp
			niosvprocessor_data_manager_bvalid               => niosvprocessor_data_manager_bvalid,                            --                                           .bvalid
			niosvprocessor_data_manager_bready               => niosvprocessor_data_manager_bready,                            --                                           .bready
			niosvprocessor_data_manager_araddr               => niosvprocessor_data_manager_araddr,                            --                                           .araddr
			niosvprocessor_data_manager_arlen                => niosvprocessor_data_manager_arlen,                             --                                           .arlen
			niosvprocessor_data_manager_arsize               => niosvprocessor_data_manager_arsize,                            --                                           .arsize
			niosvprocessor_data_manager_arprot               => niosvprocessor_data_manager_arprot,                            --                                           .arprot
			niosvprocessor_data_manager_arvalid              => niosvprocessor_data_manager_arvalid,                           --                                           .arvalid
			niosvprocessor_data_manager_arready              => niosvprocessor_data_manager_arready,                           --                                           .arready
			niosvprocessor_data_manager_rdata                => niosvprocessor_data_manager_rdata,                             --                                           .rdata
			niosvprocessor_data_manager_rresp                => niosvprocessor_data_manager_rresp,                             --                                           .rresp
			niosvprocessor_data_manager_rlast                => niosvprocessor_data_manager_rlast,                             --                                           .rlast
			niosvprocessor_data_manager_rvalid               => niosvprocessor_data_manager_rvalid,                            --                                           .rvalid
			niosvprocessor_data_manager_rready               => niosvprocessor_data_manager_rready,                            --                                           .rready
			niosvprocessor_instruction_manager_awaddr        => niosvprocessor_instruction_manager_awaddr,                     --         niosvprocessor_instruction_manager.awaddr
			niosvprocessor_instruction_manager_awlen         => niosvprocessor_instruction_manager_awlen,                      --                                           .awlen
			niosvprocessor_instruction_manager_awsize        => niosvprocessor_instruction_manager_awsize,                     --                                           .awsize
			niosvprocessor_instruction_manager_awburst       => niosvprocessor_instruction_manager_awburst,                    --                                           .awburst
			niosvprocessor_instruction_manager_awprot        => niosvprocessor_instruction_manager_awprot,                     --                                           .awprot
			niosvprocessor_instruction_manager_awvalid       => niosvprocessor_instruction_manager_awvalid,                    --                                           .awvalid
			niosvprocessor_instruction_manager_awready       => niosvprocessor_instruction_manager_awready,                    --                                           .awready
			niosvprocessor_instruction_manager_wdata         => niosvprocessor_instruction_manager_wdata,                      --                                           .wdata
			niosvprocessor_instruction_manager_wstrb         => niosvprocessor_instruction_manager_wstrb,                      --                                           .wstrb
			niosvprocessor_instruction_manager_wlast         => niosvprocessor_instruction_manager_wlast,                      --                                           .wlast
			niosvprocessor_instruction_manager_wvalid        => niosvprocessor_instruction_manager_wvalid,                     --                                           .wvalid
			niosvprocessor_instruction_manager_wready        => niosvprocessor_instruction_manager_wready,                     --                                           .wready
			niosvprocessor_instruction_manager_bresp         => niosvprocessor_instruction_manager_bresp,                      --                                           .bresp
			niosvprocessor_instruction_manager_bvalid        => niosvprocessor_instruction_manager_bvalid,                     --                                           .bvalid
			niosvprocessor_instruction_manager_bready        => niosvprocessor_instruction_manager_bready,                     --                                           .bready
			niosvprocessor_instruction_manager_araddr        => niosvprocessor_instruction_manager_araddr,                     --                                           .araddr
			niosvprocessor_instruction_manager_arlen         => niosvprocessor_instruction_manager_arlen,                      --                                           .arlen
			niosvprocessor_instruction_manager_arsize        => niosvprocessor_instruction_manager_arsize,                     --                                           .arsize
			niosvprocessor_instruction_manager_arburst       => niosvprocessor_instruction_manager_arburst,                    --                                           .arburst
			niosvprocessor_instruction_manager_arprot        => niosvprocessor_instruction_manager_arprot,                     --                                           .arprot
			niosvprocessor_instruction_manager_arvalid       => niosvprocessor_instruction_manager_arvalid,                    --                                           .arvalid
			niosvprocessor_instruction_manager_arready       => niosvprocessor_instruction_manager_arready,                    --                                           .arready
			niosvprocessor_instruction_manager_rdata         => niosvprocessor_instruction_manager_rdata,                      --                                           .rdata
			niosvprocessor_instruction_manager_rresp         => niosvprocessor_instruction_manager_rresp,                      --                                           .rresp
			niosvprocessor_instruction_manager_rlast         => niosvprocessor_instruction_manager_rlast,                      --                                           .rlast
			niosvprocessor_instruction_manager_rvalid        => niosvprocessor_instruction_manager_rvalid,                     --                                           .rvalid
			niosvprocessor_instruction_manager_rready        => niosvprocessor_instruction_manager_rready,                     --                                           .rready
			clk_0_clk_clk                                    => clk_clk,                                                       --                                  clk_0_clk.clk
			niosvprocessor_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                -- niosvprocessor_reset_reset_bridge_in_reset.reset
			jtag_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_avalon_jtag_slave_address,              --                     jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_avalon_jtag_slave_write,                --                                           .write
			jtag_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_avalon_jtag_slave_read,                 --                                           .read
			jtag_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,             --                                           .readdata
			jtag_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,            --                                           .writedata
			jtag_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,          --                                           .waitrequest
			jtag_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,           --                                           .chipselect
			niosvprocessor_dm_agent_address                  => mm_interconnect_0_niosvprocessor_dm_agent_address,             --                    niosvprocessor_dm_agent.address
			niosvprocessor_dm_agent_write                    => mm_interconnect_0_niosvprocessor_dm_agent_write,               --                                           .write
			niosvprocessor_dm_agent_read                     => mm_interconnect_0_niosvprocessor_dm_agent_read,                --                                           .read
			niosvprocessor_dm_agent_readdata                 => mm_interconnect_0_niosvprocessor_dm_agent_readdata,            --                                           .readdata
			niosvprocessor_dm_agent_writedata                => mm_interconnect_0_niosvprocessor_dm_agent_writedata,           --                                           .writedata
			niosvprocessor_dm_agent_readdatavalid            => mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid,       --                                           .readdatavalid
			niosvprocessor_dm_agent_waitrequest              => mm_interconnect_0_niosvprocessor_dm_agent_waitrequest,         --                                           .waitrequest
			niosvprocessor_timer_sw_agent_address            => mm_interconnect_0_niosvprocessor_timer_sw_agent_address,       --              niosvprocessor_timer_sw_agent.address
			niosvprocessor_timer_sw_agent_write              => mm_interconnect_0_niosvprocessor_timer_sw_agent_write,         --                                           .write
			niosvprocessor_timer_sw_agent_read               => mm_interconnect_0_niosvprocessor_timer_sw_agent_read,          --                                           .read
			niosvprocessor_timer_sw_agent_readdata           => mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata,      --                                           .readdata
			niosvprocessor_timer_sw_agent_writedata          => mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata,     --                                           .writedata
			niosvprocessor_timer_sw_agent_byteenable         => mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable,    --                                           .byteenable
			niosvprocessor_timer_sw_agent_readdatavalid      => mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid, --                                           .readdatavalid
			niosvprocessor_timer_sw_agent_waitrequest        => mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest,   --                                           .waitrequest
			sram_s1_address                                  => mm_interconnect_0_sram_s1_address,                             --                                    sram_s1.address
			sram_s1_write                                    => mm_interconnect_0_sram_s1_write,                               --                                           .write
			sram_s1_readdata                                 => mm_interconnect_0_sram_s1_readdata,                            --                                           .readdata
			sram_s1_writedata                                => mm_interconnect_0_sram_s1_writedata,                           --                                           .writedata
			sram_s1_byteenable                               => mm_interconnect_0_sram_s1_byteenable,                          --                                           .byteenable
			sram_s1_chipselect                               => mm_interconnect_0_sram_s1_chipselect,                          --                                           .chipselect
			sram_s1_clken                                    => mm_interconnect_0_sram_s1_clken                                --                                           .clken
		);

	irq_mapper : component niosvprocessor_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_reset_out_reset,     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			sender_irq    => niosvprocessor_platform_irq_rx_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => niosvprocessor_dbg_reset_out_reset, -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of niosvprocessor
