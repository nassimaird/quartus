// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
e4r3ublGN3YpnEc1UTgL6KO68KiSv6hdbLW/9fmzVn3uWBkC7UYdfyrh3ND4opX4ibE77mF7m0Je
BWXFRD7bQCcokXks/QwRq8QFlI/Ti1MWw+hNkyp/+u6g1WsutBxo9i6OVpmNnfa95ZozdiHWRjRB
Rpsswvvm9BIkMCzxavMrj0nxCutDqxL7k+wEc1M4WFMQQy4WIvul0hjYWay3XGo5wfXQcUxMP+iu
FjWzAazqzId0RqCsFw71pUeaGvaIIdChW73ICRRc7xkOT8WlQ6xX4LgMT3DZ67hAsbYdJsYbbeUV
OvLB3nkfvUf47xgeNi9j0RL9YB8+eqmdwX5ZVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 43696)
zbmMLo8v0AnH+oNid9OdwsiH0I3LGT8TVPcB1m0Qn5wCRzcR9njrBs9FE9nXv/H1zi4+/iCZVqF8
g9WK7XblbFIOy2n/4Yjw23PTzCHuaYXAhsWWPizxRzAgk75KnpqCFjJlLDnZrcF3bfRLjoj/64ay
e1SYT1ESpXNdmbc9HX62bKbFfYCn6iO5IhUuHIfNstyHyiTnk6Xu7FdulZ8SWKurO7bVb0QJ4+QF
xuaaFWdJpi2rspSOOCN7gIl63FcBt2salojDxsuuUFMODi5xB/7RTdYmmlH5bFt5q1Am61j+D7Y+
0jj8/HSQaayy+zDuWRtqug8lhIVLdNwt0HN0DOSiZAxx9wcyHXWP7lMTkLEjiKms0PWMD7q8dN0E
nUw/P5SZTwt7/YBJhaD1hR1990AA4dgGVlKVsNXmHlvSoW2Nb3TXCxybm5XJ8NW24E/MmCbO9p7E
5VfyNbr5TccApdrLaU+D4oju+Wwxyx1BB7ikswiVpsArzqaLn9BD2aZ1t68Vf7y7RW5+1Ak34VDu
5Y3rHT7unPFw8TEOIHT7eUdAeNK2BNB4fLVD/r62Zw/y372lbZ+XJRWJYLpHzt96eImVGBJAeCz7
7r/5E8jTeh1o+sCWPed8Se1fyqvcwG4z43hHA4bSK8TKF/IMTkN/kFbQvPYT10aSJd9EeyL0jkwu
kdnSu17JVmscMwVuZpPQlTOtqOE9xyIJINj9aLKW+4p7XvCn981FY4eGgOpQGleQqA0YTFHtITc/
576tRdXoN/bGPOzPIdIjqgmWcAw2EwkO3/qVeWvwW/qd66lTinkXVhApzYMNH+jAmwDXk8NkzoY0
duYJZWU3v55+4KYdjZsCk49CvSEqJkf2zX/Wuc0OTJ2sksVlMiLgCzypxH6zukGM27EMZoE8JouA
DuDkqcOX5n1umjJFujwITbuaAEWlVxxcfJbKgM3Q2/xws8Fst/y0ONusmlLoXiq2bOl9QOmZjXzM
n9S7+mZQU+I8yc3einW+d8gt1jK38xRnWjnfQA6YXD2sqLa7QxQ1vhBZ8SiCqny1eHjl1cxRfsus
0MNKC9KKiZwb1ypg8gXzcExcmboEFsTW5jzoywKdDkxvug7ZwB7btO4b8cTDlGy5ufhwB33z1lvP
k1ZP0e9V7wmPf703/e5YXvkWs3svqG6zu9Zb/S1Si5zmPhk8md7I65cxQWR2PU+GSm17EVoAqz3w
Z0WNSKfXAi1kfpz9VG7Z2nSL0MGikEBCUNHMPTtAPtB9bPhmuHUlvrleW9vqC9c5s+lUvgrCWwr/
c6VqHG9hq6mRFjRJHfevWRZro+FYTAHI4cO9/fwZgjVJK0xzomXwQl6IzxGFBJJPNY8a4LY0G9cP
cAjByEEIcA+f/adlRL4MlA8rQldGCQvpJRN/DID5rczmgLAmXizl+ytHCMzEtI274mM7U1/TfrBL
JZJD+VJ/qEb/l2/8vnHWNsJGkKqnYKhV+pK/vJ2+RWI/InjquoEyWOrQi+odANHWIsSTMfoVjont
POJyPMK9cgFHkG3R7S0XKF3N4criiSpvbLVhByOb23bHl+bScfS/6fhw+lXALajQxySBOTDTsjsw
PT46AR0VvfVDX01U7PMv6YjZpxA1yq2iinqtD360gSE50TCx5JZyPdnuW8DxVCdPuFZqjcdpN5aA
N1MRKAcrHMsPgUIuGtzYBkqS5DqtPPAp1WjnPwjjSOSqgMCubZduezPJt9hXu8uwcPRfa9IytLbP
lhDYStKno9mkxU4n5NDnXJxxrWBcIRkIv3VmrR5SWDOU1aShNRc2Iw6Pvv/usgPye15JxmV5hU1Z
Psv/tNliWrWhqBASRZRD08lmRnybpXDWP1mVMlkM8vyX2JubcVbXKw+tOUtV+J0Hqn70vNAfeb1H
QGQZytg64UAOgfjkubLgvO/nAJRWoNO353uAK0ennKdl0wv9fKfn38LkIXXz8CScwzYCl591Npqi
Lk/pt2dgCQEE19bzAkcIi6JGq6lSkg+KCen1JCSbGIVcqt//IAe6FD82OebfhIWZi6q1U0UNiccP
MDh+zjcTjOBWiDXOa50aOUu8fDgUd6PkR46l2oQz1A28k3ddxa5X5w/uAmFhWICeIew6Cqw8HXOt
4ACUgh4fcCPj+VoMr2Xis5+0vcoK/8CkzsLa2WvUskXCnkh+U1G0vVMUw7h/C6yQTCpJ4MKcJPuF
ymKPHUtMI6Uys1C4CYV3atGfEUnmeoQWqoI5CiISYY2mtCxwnSHjk2b+NmttFwuGlYIlZ7qEovZg
p/+48l7ZFDPcy4J7iuCFoox9j++3t/nDsgiX9bqlmchzs7v8sKqaV4b2EUnwP99xI7knC2o7H/LW
Tj3zANN4TQaMFCE5aLY+0AIJYISDvE3IzZPEyHsjj7dTrBlEyoTKFtW5FoDv+kmYaf524g5fw/U3
koZECNjiVWPvoxlCVK0aS+3hDuibYVf16YqKoB4H1HIKKbL0Hx3QaUrkPc8bzFxoYbFVqCIWgCDr
8hSTnK718nYuak8QvYlT9C+TpmR9xyfxImi6IR71Fo4j8GdTiKVBJfEaVVOpw8PkLo+rVPsGDEmC
3ujEoMp1nQ2GSuE4KNcyU/MP6psiL7Th6jpkpw58W5mZ3pgbCzcOBium8hSpvkmxRwdeEvqW7o74
bPaU/HqSbjwiIB7+JnDZzCHgis1Pe5S+MMngCDElUJ4UGE/BeZrAf1UgNHeZBIURHlQzVogBA4nh
/CHlYzxZ3AbDdsye7LGS2K+TM76dxGOnpm/ONab1jsEHm6DRhzz93mf1Q7WeiSwWdYNp2Gk4IpLG
8dCYdLcKO/3rjVDTZqXAtsHIJbqjW+XLQ/10VFbYgHrhotCa0h4kCHN+CIM+Mhjqru76H64bXIrx
1VZq8yOUKoVJmTK9fMvAbr0Bpjbndt5TLxORVoSCPcja8ehH5ebwVVckl3pvFUn0drpGxj4TtW24
VxU7WgBB0AqJO9NKZvdqzEkX49mUEjXabNgjzQfyf/ZR7EMzhhLuOFGpHD5NvcRKDCqYOx/oJJiA
h6fgNkQEzDJokIeWlpAg0m+EpxhK88zQ578AEbJJKfHBDAef1v0fMPZ++3vj+ynh43AtVXT3GQ9V
05QoeMM7+/lvm6eo1L0kaMq4mY6M5pz6eVh6TT58JQz9raLa+Mb4hVATqwJP07Jg57TG9whMB+xY
Q3nTuo52+igbcSMTJxsFlN0Y8l+UH8ol41jApZTBAAXJthUYHWNGDXWPuC4POk0nsD23Fr4FBwgE
Ve4Gx6awvPqlhYWm4JJYPzmTUX2VQOdLNkiFPj52kUwZ+xhmb9BMh1GZdHy8JXYy/CZM5xkTdl0S
dYoGIX994LGL0TWrBOlyYGdQtaNQl/XRT7H6UJ5VzAQuVH/YKFFsRNVmim7E5b//9shwU4Jha3IE
srIwkEcIHvFT7v91BNnHwez7BMvYjg1bDAtCc+1hqahkUhyl06kDFIqUqP6n7iQbklp/+MCrQ0Sg
q5t8eE5ndio79CcUNK23M+Nj3tozCu6uDJepNwLGntzCDAgIqEJuuS9v31c+spyUK9EkqNg8N3Ew
OSExilFTt/WiZ0kwQ/nf6DlJPPYPne/0lwbyaFp706VFdd4MZdQzNyXWrP2dl2jx0F0CxLGFn4SD
MbU+LD49S6ODAHmgZ/HZvhFWwWr7ZJ58y1Ms31NbiRYPuaHe/skVrZmKRNrI4msF+eMkfQ8B7TE/
lP0BwT4sjUhtfE1FEpS8CL2uSaxwd3MByidmdWyP9HGC5XVffo7c2oETBFQLX78QB3BDovapXcb5
syONuXnV5IkLjCoEXm5rY/q6PyZgMtNMuWUsOrvbBhgaenxMJ8hBCr3yVZfTBFl2YHSB2II8jdez
kXz2rj1CoPU5PkfmVK0kVafv2IBwMA9PIHtu5QGlEYvOfTeITD/uWfz4LpXx1o2TqqySaLnzTJF3
oZW2u6SAPxCgqqZ4ewC2M4Om0DnuSPhV+7ZBCjg8AGK9VWoTryrmOYfGJ/XB1Sw2HMHhCx3KxHpK
4Jrrtri6uRRV0EftQN8NoMNX2eKUX/zuBp7ky8yNrmSf0Z1QGnW1V8jk96hZT2JQbbozw3soyr1j
VNxQrlPKwt2k4yVg1cA7NLrj6U03z+bIKZLM+fuSH/lYHYPcCqVxZ5zkRrMoDgFTOsiA76rzUxUk
cqXfJcpu34LnKt2LEEtI9/pfL2mDlGkMfh2OMSRArfj674lS6svt5C/YVwppdzggfMJRB7YflxNK
symMUGbXPsGNSdAtA9Zc23jGXElvwKgxb2/uXUO6LZpx1NjOlGC/fqzsVqhEzsHD4ehQZluay5Wj
95kH8SsOisMNt9jQnFmuuC+6xTmszzTzC5HJKTHqwANrfjA1L22bB5Xu9WAh14+FJviZD1Wn3iPo
jfbW8JkdkmX5MMzzohITTGQn1cy+JiTPhTaqpV5SpmzxNM/r5c/AbyXaCCVUrArBd39KC6juSYEj
gLgpPwpACsbvMctH9CyABNsaDbMqsoFscWCv6HfG1evxuhTNeiUgXtggofebxxPw0dXFc1JVUIjt
pxgR5cn4mztXEeK9i9p50aCDD7tSScBfY9BF4mieU69thPivLVpmobOQYAhfGK3hGT37UeO1rPvD
M8CrtG79huHs6tjZQQ3Hupo76o9OK1vWczb54JsjE/mVe2lRJ1JWuzrTXrROvkdJqqHTxDSzo/AZ
JPmkHis6SG3ToLGBE9yCz2tyjsFrc4vJCjyVx2TpOPwaL4mV3u5BE+1rGA93XSlz1MUrjo5sFYD2
0hD7Zm/Mcw89NfgN/fD0ABM3Gs2AB5db4FZGAcyxog+xGUNl9nMf0gs+KJCwrxUUOrQClumOcgLX
K2tGUdIbHMC4alTuEB7j0RknH6C2oKzbVYVuk6SNp7rBlpAoOl1ZmkLKw9op+/dymIN9ZcNVUd3+
pFaCL4XH/0UjdZfOgMYv7UngW/is9NAMHWBz5PSxOiwOaMJJE7hqRZl39bJ/LYDukdW2mTLj1Fk7
15PBZ2Cdmq/V+Zzu6pFos4anigDaj5DwpU1BIUOryPBFjz6CPZkVyVy9ztwDXx4ZQaMgE9C36Tjn
lY/rrrJAK+lTNKfquWSQVMlw5j7qaTc5OXvrQ/FvXC2BUVurySo+j7U2N1sMZNHsrXzNAeag6UlA
Nx80d8CCl0Nh0nA2e8TQaDkohNX04R3rY8Sf5/EcyY7X77Odo1SISxU9V+9m9L3Kn+0XZwkwP821
NY/qezWpRPOLpGVbQHeUZMtXmn3Vf9Og7ga51Q4yamt34oupx0SKpFGXYMqA6Uw8MgeWyBxTL3Wo
04YdEpAOuf5iMo6VPS++nxCeCIP0iESz+LlR/KtiFdgwQ+sKBvH2HmCmyXF1vVBcDJthaSBVxo7B
ZpTXyNs8q+4+zUeFIpIuM3pRZB8GlcUYS+zcWg6yIC7i59jOIKlkY9i4pJzBJi1Y0zSdPeeLaYKs
Xa3TnzwDPpTeIxGTXfzuNw7qU2N7gwK/iy7Bfl/w34aNV3NnvpXdXeLT16SzhAxVJmkEjES4Nz2s
0A1P5J5wTwj2/NSBaeHb77oN6ORLlDZiXI2IEHZ0icgp5pQzr0drE7v8nG3HvrAyYbbWN6LHM51h
ttt5wP+6uaIoEngnW4HtU6RFPlfaEzpvFLFTp5M3CpA3maO3tQQ4YRhxc/VwMZL+ojVpL6bLbWjJ
4+SMpMuqjoAKzx72znNsnQ0uT/E2QEbTp0ED1XKAP17+fUL5OWvyK9ke+npoKPtNfTZz9gFiPilZ
QCNoAuEZLDkcRZDNy+g/ivIUDBgV0HD23DNv8E/2qSc59TkPs2olOu5lj8IK8VzddzLhC65F1TZB
ntz1xZcYQJzFUulqfEs6lqGQkZT5rguZRHxJ0yerkZlVoHJNJI+c6G1uHMQUJxQyjpd2V/xygQo0
SaECa9fj9rEV6PnSy7v0yItjXR5uDE/lBNeGmOiGGiLj9xb/O/Dle459NUOdcAhz+uC0dTrAL52y
IfqRGfpnIJdV2rMxAtD6JplsojRcF7zhzgK/0QkKXwtUNBIecf5s3uTzj2ZkxyRtW9xRMxIcedK/
Q/wLfsLaA9HxoSyXh8xmPaeSFdd9OX3d/SMtN6hwyfxq99uN06qawwtYGueO3BrA+gwVxj+U9OBn
hXADPpa/Stfmmcm7JBWRNgU2WwfPxDhUgI2fJui3Hc4trzFJcsFIuT9hLFMvbLA2U2WccQCpCbKg
VRRQ29N9EX58DUv4VjX1ox7dEEEfrDRQuJrxzd6vgFd7xUulEr06Oahbqr/dspvKe/R/GPwERVxk
uVppp0kXoT2FR6HuwVO2SbC2+/VuV5jInf0QXoylKYDKvhvY1HU5ccmEJvU0iaP/Wm4zU+Ktpcrv
mW3ek7h3xFjLQVD+faFCC/miPKuSvKdPdFNYcequJsxTf/fKjD5lGV0oS5zMaiDodhKIjOg+1Z/s
XFAIptj83t2eYOr9kNctjTJ8GgJh5iPzUSFNJYEYCcGNaPnkLfLQjZiX5dNPMxTIremchHQdOB9s
qSJ4VxDgvGQQWrNB0L+MrmxZUs8qUGHeDo8+oHTsdyf8zlOsh2sFelj7YSVEW7qAwFl3KEz2btME
AbI2LmVoqN+FS76nZ1C55WiCI9seF5bxXfjBAsmKNBn8oUGFLuRrOGm80rgOTIyFSraDzKj1fW5Z
GCK+HVvWucHWUG15/0kFyd1GT1U72nH5KI9GF8V/Efca2o/NCk1wFEwaeFaFu9RXFs6LqJyeE1m2
pokNJRXrBR/YXGV6c3NPDKIqrZqZtB2szj7UwJ6uLpSXRXSzVXnXPrWA8yB0H2L2/y4jbL/wjjw9
SBS2XWTS+kGNSjAnkYIo2FPN1ON99zczxuhczoq4f+Nz54YQ/bGK/H6Og4mShuadh2vielFQWu0G
0ZNQuXMQej6juWo+rxzOad1rpz96JZTmnYqfod6NR/ZfoutTv9mC8KG74CZG0g3G1GkBEcUx+/iz
LUg6QXiIIeg337Ru2pN9oWp6AuqYsfYophlwMUZJmoTwT6AaRRzFMlULPLNjFVX2Lm5q2Zn+uHY4
H9/kcweE+bugC91VW84v3NmxTJTXk1waLZciCVrVcrCCzwHg8JvxEyBnMdl4Fi8GsrgxZ/uTBdjD
e5th+K9xfc6Oyk6FO2BjH3asbwbiPfCAyxUH2USuIrEhwaI7QEk69ns8C4UhREUAEKbZ+4yykEie
uveTvYUG46l/ELblY2wHnREpCJHN30tuYO6hrieKgQJQJhpdNADr9/u+xiWcJR0CgBzylDv7jVro
6Wdbee6mSYF8qTPhIVpWQ2FCykT24US9bMiyfLhdUJnrlHiGzRgtUrRxAIICLMJK3VytR+wFFXfW
G8zO0YleVW5UiKwa2u2s+qdYg3WVz33gytYhXRZV6M+b+nkhvLj1918G9WXx8Thz6tPdVEHNVjHM
BWdsyy8j+DSJqrLCqOI4z1zAwJj4SOVVqFgTM6j7s0WzHI8sdC9mmwaC0PMOSc7nUpv0117q2pDo
waP5TCKkRZ+96ouFCAemKyDDxKlQHL8uRVKybCoCfIZQrBsStmBg27EgDyJHcxnJMSGCOp8bPvqq
Q3xkOo/6pkfNdlLBad/vi4QfOCKJ1vG7ekpnG1ybgL52Ge9RNZJ8X6S67AlPg49MzxMIuFUPcy2g
UjgolnUyazsQEZH1/FWkgV+IHFFOfVYvuzBPLxOciB/mIGGbRUmp35nidGlpEBPhAqLMF9kfrlB1
fbAD378/ZW67w0ruzFM1xDHfQejx89MWkQny9pSQn8UJtWJfQwo9NH/Rl2NdidDIDmLmBESlkNib
L6LxscgDi383B8wp3NvaN6QS8vZc4LmJZkdOr18YdC1CDN/U4P2zmaFRrnubsPzP+NypuWmyQYK2
VhXNs/lNL1n2Q7blRSLh4AU/xERdoIDmldvITWhu9f0RG35pLldYJQEAmQyvsQ1ySCHXjJBHmYpc
MpPaOi7Gn+z4ew2QEqFgn14embIQyyrhd7V6Rbs+9sPAtiWTIq8ckP4b7P7W5aXLcQ6HIOPeTE4s
ot9uXFBxAYVaX09/xRZzshXGI1rZum+cAAIb7+SODQbFmOFbKYLWXqmFtz78obCVfJAdxR/R5ReU
x2Z5gRlXOl8uRuFfKtLMMwZG+aueJhclzN8Ap/mRrw6KzrCDLkC5n4EF8amcw2n9jF8ptp8J2+v0
yP/NgTtAVM9Z/Kfukt6k6tMwuqBDRsDh4AKXZUpLeKbUb5ZEOkH0BZIgwoe6imluBe9SUJQdduNZ
VLbVoOmXsU2ML+FTjpNcCBfhfKZLhlyMjFTx42pRSQqz/rdOPrk3rou9Ff5E2W6wOB2iB+p6W1r2
S0LkqbiVllaLVgaM1h3JuzVOZ5kIDVErP32QvO0GC91ssDK920su2Y7H4rskkQqPU4Ykf413OPm5
fpXo34oLd/m4qnXeTIiZyNCEdYzfXt+BqlKGN8Hqz88yu1j/5QUhISVFO93QX6ga9wRv4zgURUQ2
Ub07jwFL/uz4YmNNQoICbIqDsuMmtzMilMhf9vBWBoYYGbp0tMoQKhXsoN0YNF3hVP/i0ggIRqSf
OlVlAi5avL5N+fjKvtGKi20s3WkoTlIymHSID+elpkly+JO28eKry6UQh2y7Y3nBtzvIfx0Rhhkg
6yJrnRKw8Zzu5Yn/Ic948mAM1ds/O+f6v9UmI8RDp4t0xqyYEaXzznECSdPhii9tQL8JdCwDfJH+
CYDvfLLko5qbwbNpeIFWLX0gjBfnBb68WGoYD675YXEfrVvS8jfHTxzEyF/fwpLE4LXuBKBosixT
KCTDotqZk8X+qHQ32GaH4EeQa2MjNexvXiV00QqaFn1TvINRMpepWfMvhgtfv+zQ2updVVG307L4
YVIhoGpdGd+Ccw/Sn+a3hYE1tQJsjr0vaJVCo4j2/O7NjXVa3q0/zQihNefwUWPEDRm+sDYAg5BZ
8EaMEkCJ6b7aZ/SzN6i/h/YuXYKD7UCuPTqpgK5rEG25IeYG37nZhD6CvmQ+73mzKCInKnq7lZ3t
k6qkXFxsX9NSPQt/nRH3FAu2JVVfFnyu20z2hZxHAJ3ZN5nhNm4fzZMVPtxYCS3JEShKch/lqYmk
CWNCy5Dl7j55ywH1Ukcg4hXfDFjK3wkHXl2gJJ0xZWGVQEUrzrEJPMDRQZCzjQHPhDHyTlu2nAYM
3GB+9POtjetRVEgZ6nqw2RB3amyKqZB/DhvgtlhTGb0JwlcrrkFjzbphkQVQFrF+Bd4Uuy9vqBcX
gKaweBrC8vMu1fGsgQ0O9DdHR44SRPSfWT7PpdCvn1Brwvdd08sv01WZb9uzyTktISOnwn5usTz9
Da++OWlcNM5jyQsC2apMEC5Khcj8g+hQ7ioeFhIdCLWqZ4FZ6ePERIdi0kk2EvhtjW5uiDQaG8RL
JuzzWrxbvkPqegho0K2ejJyvarIYlpun8u3LL1a8K/UGCOoMa0wR/HcukkQvUNHais9tpMoRI/G9
CzYS5phC3KtsL9qnd5OPgiIZ1YYe9IesFBulhnzrbt+xaiR7aaYak/DfMNUWE1/gGDDgH5641q7R
pMW0NxbP+9bqqwz+XClfZgafUGv2pzJtZp8oEqFCtrpK0pqAbvtXPJYkXIWPiCt3cjltX9u/QPwY
AAyS35n7rlcwglG/XmY67Oqb4JS302Fo/M3tJcSYRtUfvTuPU+GL9qGSvL0Nvbg3GFI6BVjxY7RT
WnEJ6dXgqp6vI3kFxtH4vJaNFSzn9Ceu8k/FNGIH/K3BTALBcqBLqTZfXfO5fLojrTWjQTMF3Hg+
U9DDSvMi/I+aycG27gQYwYtTlwibLG9MPLNb48lbcaGP6kk7PvUJmNpQWlxEsZeaLua/42hojvYg
lQoSbjajP6sB+0DPirXxJkhdJgoxxXVXpbahC9HCdo5wRmXJVI6Rft8H/8i8kw0m/tEAYrXDOzHL
ikADDhfmJmx7qyAnzMumrXAAHSflC+wruqGL/mR4L/Mj9Kdp/snsq6X+GK+DkKmVVtWBMZ8mwC1Z
EiEIS74cE8qWFB6WAFffiWrNPA0PU3iYsW9lc7wdUreWLBAmEk2JRd0QVjaHafyD/NDuNEK90g+R
KkLa1mXaaUJYSs/UOfx4pvb97K1l1jdZmCa4AiO/nlIRyeu8xI6jYfaSJ3KY7zlmX96dRx53xVE4
9q0LCsxHDzZ6qEscuz6mKfh8YIno7QnJ1EbCXMsSEdlijrKBkRqa9i98X3Yy36RarJKAMna/sA7d
zQp6IcGsyrPDIPSMCfbtnAX3eOm0XnOUSZTdIUvoWeP1DloinWNhhlSRBFvEynWaN5ludkks86SN
bhNI2Jkw5f24ySnMMrFo8haqXkKy1NZL7AQ17DKLSnqPFukJld/clZaRgkE7dQ6DyXVo7/UxsGut
tO+SC3tf0lCQT8uzFqxtJIKIlsW3ypecMeapKgLpN6CCCcwZowHVeMEqFoPvREIhiVT7S+9AFJmF
cu7KkbMZx29n7rWciDVVJLoydo3XwlSZislw214Smws8JFDXUVychYNbTVANf/8hIOdUI5QSSlJW
5x/r5VEDsp9OWmVr3SPpd6t5rHfJisfF4TcSi9cPTrkAL2Y6YYdA9cJ1BDb8usbseFvt6KJhv+bt
kKjHHD6LGDcjvZtAbRpie4G4KJB5QBsAxICJ8mkaYoQKjETX5jMQsSBBRN2ckzMHeL4bLH/9uRQs
V/huvQH/7brAHuSiseiRQYxXwMRYgwXfSVq5LYi08i0W6DMnpsEdpiZEMfO3jPF+V3amMhk00Zd0
C4O6AIi0WFGkmg3F+EB+HPL6GbuFpRAms0n8Q7BVwOupQHwf4wN8PONe9exY6yEBEFHWXmDgsv6W
pdqeBxRp3G/SMfJ9uWgrAbycRT+zo+LUwQOi6HmS8nu+BHtGZ5rNTc9VhY3Pw7Zbs1capJu/5GdI
FTDMSAZi7ZZpyOVDgScOTOJDf7vCaasY2vJohAZMu8cCM4ughOV1mQ4AaLzEl5zgVa4GhyCK0fGr
EknhjAh9xcSaweQI8da/aTYIDsESim7Mr9HvlHEtie6W1lfJ8dxenOIJxxb62w0mKMTBrDbTTO2Y
JbfG9G2lHZewjyyKFYmXghqlISHuTcbsh6YUvQhM2DWkn7PKoxJ1wLJO516cPcR5NKJ5Q8hv6IHA
LUDM9gGolvi3iLcVb7mav7anW93PMT30sfmZlsTCHxh4aHmp5OYJA2hUj5ZeE1kdg+2w6X/H3x7m
pG4dA16sdOWeb5kD/6ovdbNBsI15EAjLHll4qd5QsnWPNG7GiYQ72+l37UmBQpiBwqcyS9ELZqdK
8AP7z0Ma+wcPT+2NUYcwuVedGnNm6AoIF9PRspq0OlOkSEgzzUji8DYD7/4ah1yGfeTb4fhqPlga
Pc55kzDbkcXt+vzTp07t/2r5h4G6aFoWEJEaHvtiwzq6EmWrd5aHgOpziWcddnREv3Lxvi2ajPFY
GyP45SA/A3cjLpbvUxdu6t84PZumj8w0IGQFabKAG11sqAhSWPN9vwjqxKRxe/EnG5azzNxGdbQF
H3ynmnCxlXKf3YqLzy/qhxsq0IuKkAajrucUBimP18H0cW9QGjL42WAKFatELZdSlusP/u40Rxwj
w/A8hQKDCIrcpHxyffSAL8VEhhXn9CoLodCbJuulaHeFyKkARXB9dTAROgh2cCuFQ3naI4rOJ9D7
zZ3Do29EpX27/I8V6LfAEPRB30vVT1r6+pRzohM30PBAwwdxpsTtmNnvd3fY4ob6QuQCCWPCN6Jq
k1rYG1hcn5BKlxyFl+JPiWmbGW2MLDB5KuKMHsQEbBvg/dWbUz6zLVbg9CyIOXfQlyBTk0AnZLer
hWNlxH+mXlVy5oG0xSvsOerca6HX3FRhviOBnOysr2eMvCx/5fjKphyRNBRY3EEVShRQpR9FwWq7
7asRBVXwHlQUBO99qHkOnhEGz1le1odvZctxM2bKvjqONL4RXz/m5hbLltbPyTuRmaqN1DAdL/rX
MxznBKSeu3YJMxl/C1UGqEPuHYq0Bo8o6V9qiY9W6lMizAmb5blBNWlgDlDgFKVZuGkzYZgDkm2Q
7vbyCwdxA0xRGVfYDFGf0H1tXf77eROxemEUCmVG6db1mFcSFnq9iCekpGE45OY+NtLQMyNKOjkn
CONrp2nE28+Ue7ld9lFnIHG9wdB1ETTdr90aV5SEuHrO5/hhVUAGC6Op6lTapiHOfAtj8XywXbul
qDZgU5m6toOpiQ+SOMvUs2T8+a+ln8WEzlj4b0vQaedizO4bCfLHuFTRAAqu/qwP3T0ZP719IEnz
BoBZfKpcEXE2bu+i28aZ0VXI55wd8haAm1B5st8myKOTvOEIQf1zfnCtzBl0T9nvYL2MYlsbjzBB
CAwzTtwWQgeYO5fQ03GRT/bEpfdiyx4quXBEoxCaBWmf+HO/r6mTf54IWU7idIaleEDfW0OB+HZU
ujvRNp4HjfISjop0vihxhPVouQYcXWlSouVpfBSFxmudKjMnBIgzKg5He020vVEdOXo9FbDyTGB5
mSUbdVmVJPMkCGJMqPHR7Rq5LjpzYDek6BQQN+vR0N1ywiSKikCtErC+x8AZVQi43SR2H3DJzih3
PfLQmkdDudvHUFH7fwn0hGBz58do0pcwBTVrLs5JjRkWWXzXI7VWc319MtiDK2E3XCUv22aCNrlO
K0gswKO9CXvPlY1TDzPQqQ7X1tJeZHc/ix1SHsbYvrFg+QB3VdUpTM07VgqtoG5ZF3mmhYAiAGqZ
bJAL/I5Kx+2E98ywYClRPqqQ+RNITXiJAZB1Lp320jfLYRwXH7W0RT8siCP2bk7VpyO/pF+eDJ/R
0ZI3IxIoFJZWSkN4NYPOsS1t+Aznj6ikTe3bA8aiQPyGnDZYug/9rO6TN+kwQoBeVuO55oRC1xTY
9uDUWpyaN9H9HWJGZhHxMBjyZ9b8DoqwpQL2LZaaxJgIccE7oUIyS2yP4Vr4FRrk5rGRQdzK5fQy
jW6lHuIgPoUwdyVpONAl0u+S930eGPsRhe2Klvi2zX9NUMoUh9UvSnA3CRaCpoBqeIhIv4KATRE/
lZK8IYIlsObUZLupf7fcmCE0W0+5U4tunWRZBmjKtuU9MnChySIaxkhIkJZRbyAJFd9F5L2NdyIe
1h+Gfo9GsoDoMbUHdj336j7qDjUjrbepSWfqDY0k2v7grwlONekkQ2o5pVr+y6cDVYbwFgsmDc9F
E5jXu64006C42kdg+cM1PCvll48QP5/BH8P26MehxLoupD/WHSHoY3KoPGwvRvqKHdPgi3974WHW
4OhvTdKUw7pSlJg+PC6/nwWPMy/WamTxpPRpwbiwQKGFbZqdVe2F68fmChXDtaylybn9x7r5kXNt
KQRK6ZxTgHrUhRd57vpF2ZOJbmyLYOvC5xAa01fv9+1uOZVoAoiGThato7HPqxStrE8Q7LR2DD4j
O+0HwwW+q+SJBGnkCUUw7INEaQh/lHeaRo644QaO5SNcbJrv7pZmr9xewcL8XIs1p7CCEneFN6JI
qYrNxh2VBU4rVsbktgA/DYpTDBZtq1UkcjtZ9mghWpw8+fWLmSFjtvGZ6VnkGSY5W8gS9ZEcpgs/
BTG62oN+oeXC4/ZCJ98LIWoECXWLqumThU76zU2LSM/FZCQqLplQcK21FKZvx7zQew51Fi1yQtvV
Ju3kBTPsZ+xYyPgf7k/4ONd9bBu7NJuTqN9JWfvvXdbTKZ4pFpSo/KkHQK0S7toFXeeTFUTl0Oi8
mbw9Ea627auRoAquqHLW3EJAIBNvS9TCyGDe8mCsvOm+/apDdKEyM2JJ4BA31P4JEHDPbg5RQa0Z
/RpciTrglK6twEW06/l7pVeDBZdZJrVHPEVaT+a/xSNSltwdUduF22HTYdKKshQ/kQXxIkPA0u7m
0NK78B96qr40+OWK4eUIy6JHwrSfxKggPvJ57DgORyvOrjpVLzDXgQjS1HGuLDaw8G0PgUe156dr
PfCDUjo81HT0Pz5v6BiwNs/YEA38HIq6MGiaszqQDsRAp9asJQtskwbqTUBi8EvvzG/FxNA/eXNX
f+WOfuQo45A9YKod6sX+geq/FtNR943qFYIxKErWhqINHU2aoVLJVPitZ6/h5amzU7GgdOaHUU8f
8WwH0Hxk6ZYYiQ6pGodIuQ7fRjqAyUfGxtBmdVGmL7uyQkJXt2O6bahS1SxO8l/zcFTl5V6LSXuk
pSWHGKB2S5DHkK0sUryM53Vhn5LzJ0L47znYUKq+VSFFZEkrpHvxCSdUGW2z4hobjn31enz6cHbU
YZkfR8c/o9Fefv1rUMQICa92aj0m0QZPuoz0kQoTuQTwGvec66eZ8rvis0FsnuYbqpn8LNQbhEi3
EUMvAIqAiqP7Fw6vWUGYXkoF9wc6DumjL8k/0j5rK/m51+/UChcolt5pVEslKFkg/df93dGF6mbD
cnS9n/tef5he3ePdgu4OCUdb9SQofaLiw+NFzj2gfwVCAICgzVzEKfUvIrFgMFO7TfvaGojFRgtZ
aSqpWjuXOgrKrZ4hyCLWrihgOlpm2vr+c0Rx/HznCoDUyZvTPgdzWGfQVABJHAcZF4yiMDdAT3Gh
Lwj1lH4tZpGfCssNZzDRDFiTcngogE/42WPtHNsFhcVfcwGCqhXw/NxKbLv8Oy0ft9oAe5LBaP0Y
38QD7JA5fBtWc3kmFd0c4OtlVqMexamKOMuw7vIS3VtjzMOADSspvqpKwdZ/q/NLaq6Ja9NNI7eE
82UXsnrWRFiHqtI8mtpf69TNDxlALyh7x0XY9BlxST7WYti2fhqFOPFrQiDZ10FrNc0k0+XFchi2
jBD+9Kca/CuOL1yL8ibHQN5BZVhfTTl8x/LZAw58l/QFeZ5SsJmpJDbMg3r40Zxj23MOlVHPM1hl
V4LNh4WhUpvGKOX9Cm0wMAuEQwXX3sn8OKpp5P/kzcKECXAe3lPpWN1q6ETfSHEFuJbqxoyvrNxG
NyiQMhmmPa4ghIGDtB2+KiQ2MZ/8jWq4aUlCy8+uGS8w8KrHjZ8ROiaSpHGieRa/D2aIbl36Q9Kc
Y0P2+9QIs7Q93IHqAD3dz+t+EiRPRZN1ooR1Ac031MckOQq6kfQ0xYAK5qRKv7wTU+ufLDs8+KWp
wSEzWLzEk3NkBOcy8cFHOmTtBoAC1+2jQ0W1GsePNcvBbyerDR8SWpJSqSY/PRRZ2F90agOXOUaK
2VZkSDobV6t6iefhdk9h9PnrRv7V+qxcJSVYx1BpW3tF7TBXZQTaqRNv3p/3sVWsU7+BOgZobj/J
yyk+yzNGwBAzcFjiDm7TFEuZeLeKmyanCSh1zM/St52iPTWT5bEvTIR+AyuuWPx/d8RrB3eRCYAA
x9+a/Th3QqKDd2K3P/yeu8Neup/Ics63+cZr2hMJbqlJX1HV596y7lvmyIx2kGdVclm8+GTkHcP6
2aPa0maWsnW7iQGa2jh5aTCFSO2RWeUhLGae8R/YEHyhwhyPcIxsUTVlZXPSE2EDIHvVaSAxX6aJ
1VjwV7ceksvOXEgw/xjcOifdQmG74M7YUhlNx18xWX4thNKJ5ykpsgKT0c/Ay+j7//JBlhyq4T9S
E8jayWYbyl+2XKHp3/cxH/pTDqcTCW3pgFGYueDQp8OeUgJ49ZdfUCaXvwmFba2uhoNS034NHMys
kp/oXiW3yGSMwYpVY3Bp+iOzFXVg7aFKWJWIt6reRxqIMuD0Kun7puQVCE0IFo52b2Qd3Yalw7CW
t0BqBD3XNFSOuqL7XuJbMbF2Sd4Fzosj5pcZaYswk3EN23Gyc3IR5J7hlVt7iovVfWCoLxgZsTAl
J4alUaVKxPbndvKofSVJwd9J8hRnRIC5xjL7ozi0IhIsDGlKaZ6NdwCAzkgxIZWeGuV2RR1sgaJg
iM9AhoQGMih8p90sGNvhggIUMRooeivI5NSAPqHXEqpu8M1+aecJgvRsh1nlVNj0K4mPvQznJuht
Ujk//JiKpL05qBb51esqsH3nHVfWv3dlHYzqJ8BEV3TWpDr8kdohl7ZJRKq497qH/mNV+/cn3p3E
36HCmLL1nUo9Gf6nYb67OtA+mrnflUZpYTUbQy+bakdW/RRhiWT+9DgR4pjbANgYyjCsI1mN3gOx
2Weq4wDBQyTWBH8N56aOypm1WUqtuJzt90gJBgm+muo39HMszxh6Tr//KyhV9i+E5XG3cOg0uaFY
uf914Mr8vhncbk4mA0Qgb6yKf7DdGV+L/B1Uwm8VsU9dABOchzplSP7P8BEeap3sGo4KgCgSUwgB
rR/p/iLSTYe3DsOoiK1WpSNZ35LVdBGdcZlNJaNRCNmoelEeSBG2QYTWVmo6LA+uAdFQT72KBNqC
J2GnI51pi6PMN9G2O/gdtv/0SnUqk5K/VrCoUEcMpkTyxlx21nmXKiHZadl9BNuzrHDIqaDbM/7+
MLiX0yKac1cSJVB1+mbJ2D6khta0akUeKWKMWQ0JRQnykONO1p5LVuFn7IoO2Fu0FJSxJC89MTRr
EAplHu0g3xfYxbtS/9yLzzjeVrMc2TYmxt5nfLDsPmewzqQQOR15Stv2MSCeDoRJqsi//Rp/v/Ok
uFrC7QbIbOYDMYZJAxSu9J09GHcn3bY03MitH5tj/4646p0a3bjXxWcwqLtXFmOaXaqzAASl2LRc
AoD+yCAD8QECB5JdUuBKnLoDuX+Wcsfa/fqx3BcimSwK0Qy3nLNikLXnYJSGigSOrWgXMr4pZEpD
dlBehYb2x2Iu9a/o8RXNuLnNmfLao55J7MMqnrDlY52uVhZePm8tOWfQhfKiJ1nEWj5z0FbbseMQ
Us10lo0T9y5KfN/LynOkT9OSq1LgY1kP9Gsx4vW37iyHqOZCPY+izrahHvzWH5x8p8CsFpRSEGVv
QUbg9K6f0Z5GyHY+ogDAJ7QAAinKCtEpv4fzd5K0IoMujN3U8y2/FYb23CWa8uA61lYWxffVWnCE
9UTGbSCTI4Nuj+A5LS9xglra5PLxVAL1n+3eYi1Eg0nrrLuHrgwxxpr/+58iVxa+OVj7juwJZ6Cf
3XCIslSgARXxDexxZk262NeVudLiB7Fwdb9Bx/mJPYiYe4Ag4HK2VDXYmFc2Spc61yEL8GVo4l6f
NG6TAI+VKt1ypKDZm1pjx/lC/bJ9q9Khww5a63dymsP0vh267CXGHCMy91M1qErHW89+EngIcpPF
bZtvO2yHzpkjjYjWtg7w+KG840MqjNjHeoLqR8SsHrwaZTxMe47u01Ze7SvczXC1xsasFkFV59of
5omU9QmAUUPn8syQhq+Z7Z100FDRvudxRB5u/PbjTNVlra18ivxFBwy5fOP9j9iNRE0+2Dp8qB+2
/1DHOXuACQ/Qkk6iqxWibTtLROVjo1SxELalwcmXetShqRuaaKpUVlCgMCS91jC6H/zYrF+4dRvB
ZC0EZsB5jUhvXx7SHu974XUDqEixodfJBXMbvl8qFGz51ZpRM2lOvN/LMRlYvfxGTl/Zogcrijxy
AN9GxIRkaeD1ZEvoaLBtc5peZaiPPjmN5urgwW8F9G3gAjvPQa/2BR6ngxkLVz7jdI9RqzbHZ75E
gymdFbZf/zqnDuOMRCd4EbvHF8l00cXtFYuzApFpqLEySuNVn2WqQrPCF3T9iHx/D5hCvfZ7hO+U
uReckqscHOJ06Exu0fasgEqgl+fbyPH0zj0LhHr5tlZ0XMFnXsWqaPdShro5Ym47M7A6kbMeNtNx
0EIv2FuSSUfcJdixtuq1zDoEgQ08vIa9D7LRxtCq3/lVbuaiojO+ozjf8HB+GotmWUaDIFL5evvN
6GGNuX/pec5HSQZ0N33LcSViXaxRnVAOyXXkPer9LSmGfcrsHb7yTFl97qDVi9TQ14YavIqR8ZxE
r50PLgm/nAbY0WMNTT3bat2eqPmPCwIwAnWnl9OBJyDuszL2qLQmfFd4UAJSpT+pZBECHHYsu4aB
OtEl10Z9VaJvcE/K5LaNet8XBXuo4QKBlu/9DZtNCWBGVFzhNiTY7yOdc9JNBSyPES/w11KRaw2r
TnveXlsJhwgHJWn0cYyFUKd81HZiEywIDGtHE+5Ez1qsFy01ivOQ1PWbcJodnsyUyABcfDG4pCIC
l3k9FTocg9XoEcpmYitQsJxhkA7Gha8GYN98sRQp88Wvr8RIRyw2P7WvROQkIKwqUyB/84VBiN2O
RsImQQTMCuYnedqsbF2BmHOs0gVlyZVZj7TwH8nBOgw4TUX5udGX0VP37ucK+fQcxtHcCVRrNQWo
iqKwerVW+Lr/7w6Oat0sR5RpUzfpawJ8JphPBkaheQ+oZZrMcgK+khOHB+xsZxF1JlTGWDzvEi7T
T3u2RTliuFczizFn5uKtcTB9/COy98inQ9ahykETJ6crCRkkLQuIS3pApB7NpfYiy0GyJI3JgryL
O9zV4KEmBkvnUyCNVSZzIoL99hvpKtaSQfJEb2+lfWMSr39OdRIo99Js1JBw1fR6S/O2O+UnJV14
S6jZ5lr4zM2s+YUr8kvsFZBCP47ChRHQDrimgCkytiMS+oS+VNLSk0rIHbW5A98NkvWOsFQdpRbP
U4N6AjrtNe5bZ06TMeq5dRGs+i21fH3nnBk2UeJ7e4iNhs457zzXiT7vzlstjez/dxpttQpi1FzH
mM8dd5uZkDfwCCueq9X3o61UoBxWHd2Z7iZ+sOdcJ5Zzutyo1igQKA6k0cOYCANkIeZ2zNrzMesT
kguZ8fg1M2YbrK/AtogREOlJJOZxEellshsHcpbbY1CzaCePmM2MqJX3NwDb5+WqBPCiJm4y02wk
kU7MKIQe+OMHnOnJBvN4kbpGVUFT1BNpfGkSVX7ds7zpvCQoRoMZNhkzsdls4xDoeOHoVRmjsV8/
qMFCZB4TKQ5V0uJNNtGVz+i/3GpIkJTWNCgzuQJWFPn3lgzUcpep4Ga/8+8m4P7rQB0B5zeKsVoh
S+ykfpTxD7JYaoSv88dmFbntsZK/DAEj5zJl0Q3QJqd8Iorm9hR8RL1NLf+jd0JFiB/D9WpBSr9H
a22UpXj/40Ivw/LyNLdfx9qyL63eiDHz8ljHwXYvJ6E2KJBeZ1WSrYwbVaNwNtK8TP8Ts/JIbvMW
xk1OKXFKZcgV9d2T6mWZBrxnMlYrruo5Iq9qcCX9KTIjqZPNZJZZpJAXmagjDhZwW3SivSKMPbfB
rI+CYXfYTcFACt5K0HRMGAXEM1CIekxv4QPudlmQRZNrC9I2qZe+B60nXoJ2GxCG3bR2Zt0YB6vh
+57Dgecicm54KVreMeWYzonhSd3FGft39MyyFl4qdLnykr1NGLaGQTmXbBQVla7dDb+oDH/2DVX5
rl1s6jRbcAsVmnqzXTvvCofiXVJZGHM52kqJda1hsUeq5A6Je5ZPm7p2t7ZI0AInqoFB7FSB8DTk
6HuF6Z4K0n40wvYrDXb4sEECk6DKoe986oWJBl9+mXsLVA+AfBHnNnA+nRz2PmGDkGmkPuCly3hT
ujotJO2dIdzXAwBcHGqK2Hydpf5DITs4QSbKNkS4bEDW3hGEb8cFnhmsw4MnGzNJi0mB5mM0jXh1
YLVYwYXcM77A7hsu6i7b2UjURUHJrBTAcnxnbJx0pjKkDRPadjfsqvRrcu8GnMu8K298RXnqigKW
BH/Tu9qQ/wsAnCjQaQwaUI4UBTWi79fdB0usiT3PeVVLzs28XDJb6kK3Non5e7W2Q0pTgge41PnT
gGD8BnRTrCWGK14HcN+KvHKVEzNiMDzAPlNcDrh3maSK3Mlp7HhaZ8fqrWli7hhh8lZMisQny4I9
Goq8dCjp9ZgiwxisEET4M5tlsqW8SgWmMUDtvdC5oUp9doamgFsYMFbMx6IlFBdjDWSlFZtDg545
Yd1cuF5duljgHRkXJ1C3tru2V99EJHePWQe/xEAQYYaJqb9my8FbXzPrTjIn4hYxRIqY49vWe7h6
DdezFygetUNr1B1ZompANdmmNmazhQ7vemXo/foJyNiTgPWQc700deMR+DkqIwSXucGgJGzBbfAQ
hj9k+VmEQCuDL/rZUyvde+gy3PJRALKpC64suG4qSeEOAKnrslXSmPMuml/2R5XU9yY6rYrOmPc4
XwEEkWiwHKQ9SW8gXu4kLlPKLtTPaLmrODJ3Cl3Ywsc4WKbQK/xnSswMdowxN1ZIkgnMMo+5OPH9
MwjHF5vtlyxQSv/4ZiGd29jN0No/+eIleTCS51pr+psgoyZXXtt0ReJibHsf9HLZhb9EJhw7+P88
34qbOsmNjp0b29U7cKwDLqUu6ay1ifpQQzu5FnYAZjSAa2trlJ8s1gI9mlCrusXvlwFRxMnm2+Xo
SYuI1kgySmTJ0HPS/dMmU1ezH8AIsvtZ/gb6D6zdo4D2KHKPorNGnk00BOxZSiJZT/MlCjb0Oi7u
jyRGN4WpCDlKIGCdBJmxIwIx/Qsot7O2dfzC5bs60aunp8hnE/KtiQFA6qHj3o1Boe9m9zVA1Bgh
/to57VopAJeWHL3BGrZxZNNEDUBY/POVG9JwGsv2YXXYIF0xi1/JO6FRKTKfu/kBgWNq6FqArCDs
RHOpiM/DfN/6LPyFi8A1EJIMpF6tpCGxA2XpG0ovNmuPKWqWdapaJyZThWAj0JFg9c2hRkUcuPRn
c2Umdj4ubW3Nex8ylY8IoH7Kh4cgJ8ww8RbjK/EVBrVAe9PnAIDNLt8zqtPt0BI0GBo5XAblv/mQ
ULA2NbJzSQkP9NQBGIHgahcnwVmYOseNK+qqvAJSRNSmS+oR32eXC/4FWgib1+nLsf0AC3WSlWPf
QeoYUdj90n/DKrDy2TKs9hNPQdJYPBA+bYxdr+Eo8rTcPuiCHRs0mR5X3VVsdkiiVuPc4f54Wow7
BNKat8oJtXEJKAQPPnAPYfeKHH4Z3rgHHzOhJ4HdExNDXUyDAHadVBuTb/z3wdxl1Cqf3GMXmu5P
NsgMyrXvAvI42+SouwDRWpWBmjit+gfhZHcMmgO5gAtgtNABtCHfJfa0qG8ppAI+962xvsEMib1z
vxqcmcWe/kr67ltcN0flMpQmQjRV+hYUVota9PVaGeixBKLUfJWdVHxwR+OPI7IIU2dRXUna6zNt
NP9+Bj6HfQRGHsa2/k0g82u/99hJwKz8QZbVzpQOqVSgvGAXPKdDrKlQIZBos2XDE2QIAoioTFg0
W2OvXRydkz0n10MaHtU7swgbnXi41CN/goCvhyKwyPvSwcHOSg4I8VC4K948khUtOTizjcBhAt/8
nvuZzDcEScz71UyIKEk+cK4yniSmOdiK/Rv840HNd8Gr/JQIkq0qOU9HtQwZ3h4Ol7e2VLjGRbHE
4UM876LzvD3Z6zWAF6/gNywjWi75/xnene8fB4KJhP+tDc3MRH/1W/7woUQBxFc/0bgv3q6Ppj4p
1b3MXPlUHW2YqDb5NiuQRnKU0a9PRB7wiz18G3ZuJ78sdkLGC0YuZTXkLFIOoG3/jPEyjAXhHG4Z
f8qKu9bJkLlmvwNsjEpDn3aorMGrbL4AjPieEAyZgiOs7rVadeFlskwQAZuHJfBAm4X+oS+zwVOP
jDTrGGZS+pU6Csf773nLTayhtGz7LXjM9zYmtQPAhBK4Y2ET4LYj0okzOYvdav6KAHcAMvMKebPQ
+zW3+n7E3hId0g+8opa1NO4hY/CTlwyxT+UWhTlYjuZXG91SUY4eSYkFkcb+kXKackx1tAx8wQZc
DnDB9rH6pQ2rjchUEDo8BeJIu9vYHsABSbwIesA/kAOVYA8d1rU76c44Fsw+BWLGZ/ZH9YwGi5w4
nyjoHPjAuMlDfjodP0NGDp3rBpN+lOUFUSAp5Liy6KlUWjnbc9zz1FAcpyNCTHPi5rSqCW4KKLxY
IcJ853avY62qL/WaSoM9ttqVlAJ4iMV5CTgAjyFRuoXk2MC/UnyAsFKqhpdZlIA03rTpnigXyWqT
aXv0nMPqo9PqlSMHyA4LabqbxNP9NZnPvhUzEx9wjgCb636wIpHhX8Jo01vMNKxjUssxWZ8Z6Anu
5CjMtxjTyzPBnSPFTqnZBx1xXdh1V5jbBcKd6wPJuJZgxaV/s/LlO6CCx2A4ActzYAhLKIeh7K4u
LBtudAJfaH1vDnrBIrTPFIUUK6vaplIPpFsK9pp6f0M30GCCulIjlEPVZmf41hZBfkXqYTvPwJzP
N2RUZ26UL2TzGDhY5vdoogbzMCBw3qffqIVu9CVwl+1c6Lgpp1ESiOA6WJbCVuO7/nF6jPwaayQO
tu6njou7Kf+N7+fZp+ut7OPqAnSyCX4sVlC7PX5wbMQ7jdsM8yjwsOgotGa96MX8uG7Eeqeoj+XF
6lwQzJYVtnqlNGIvk/McwOuq+XatL20GnJ8JeKX3n0P2dUEl626ryFL46rfeQN4UX8B3LGLslTnl
IzhwLZh7/8VVUXQSsCaYQs7pjDd+PWMqzFRZEZo4YIEei8ViFH8rsz1FdKJeDWMOLHW8Z1kcraxk
r+CQUJTu4WcWvZk52O2ZHuNORvwCnA5b3lyKeI1YhSMASAdvnavHAigKu5fi+tuxeYaFKbf2Ixjo
gjVSRG+ZShzNDNXeym9xa+tFyzEv8QgniDUJyhISYakhvjAREjl9oWhk7gF5WgehpVfUttIok+r9
LkwD4mkKfL8+3wspx8ytz/rTMmPJQoFLjEynhBJ4ex03s5ix3B0v1p3VVoaOpk0G9lkTv+qp+s5d
OHMZwWTQVCB/xhKqvm9twSaAwdJjs8t2GNePdaJlPbBf96UmO6M5WW2yR7MhvpYic9sx90FpQagl
7fv0wprSjQZu4RmvU8/uaw3XrWi2XL2Cp8O90mPSlt7Vxb1d0wu9bLXYsw/D1Sd2es/u6basZUDF
wniqyLc4OXUMNkEF68vta3FxZ/2Z4m9t5zDINkKPo3TW/rOA89NNiHo6iizISwh3rJp6zpoVzgjw
rt4/940gt/FMH7lJOUESjJK4VgB7VLg9hdVxz5ly/KAWPY9II26rORstjzUSPSkYXPiqU94TmgEI
/ot2JsvrdHXmjub01Et1n0CVR5c06nj4yJxO2je6u9m+M/Mgnnc831f6MOy1wU6qMn789dm3qL3y
YLmcG3m4TOQzaGleFwn9+8tTC9PIRt8q6BGNY+oYSUVFpuYQ67zjE0sw1xxtcI7MU9cjM5RYzbT4
gKe3bGONJwO6ykjvFWwNTOwypIxJZ62VBm4pdnG55NfZZRGvrw/d3y3+vj3vexiZrIep3J2eIkmG
MZyq1w/bt0ZMmDbrW3C415OCI4mcRvEu3TgWadimHQKsv2nrZFOZrKB2nLxZl9AVPlPjWJSW7X2Y
edO/KyHdwIa/h1R5UjmYG5lQgDCnNyMDbjLVlaXX79+MI1GGQufeC7kgVaZ7BvrxZ/DVrNgZtUBK
0g7AM9K7WpiLNnvaFToRK8aHWPDoNbNSLImlnX+xXTKyG/RbhPghlZ4mncil/IkSgLNJJZmmUSRz
1fyfhMCrP0gAmVhHxf5JnMmWHTrmPb3BNkw5c+MBAHPRTfp3i1cKPCh90FktclU2WacNwhpx0J1n
BGK36n0k0Gyj+y3xhdNllAbQtiIuVWzagwtRMWspOLngZ6bQY0UnjYcCe3yWQJJ150sbr3gCWJbx
1ShFnJ7rdanp4R7XoktrSNeINPp4VWCgqzpW3Wm+uZvi0TTAXQKCZIKb1J3nNtmQzTMGJYRS9zR4
/svOHUudvrZAYfoNt1Hm2ouaniURhAqyIy+er6c1E4EZeUG/v3GFzyMgNT7pyfw6WJn08oELvIpx
BDu1pEyWa/JVmQ/BKJerku1O7wXLkISCJIbRdbFvI/F1D8r/ytKtp24faut9SZghYQlmUKiiGKX0
VC09l7ZXeV/iUVhiD+h0PhBS/qj2xpnS2AQWKSp2xSxz/4U7b5svd3JOrDm582dlxRLQo2XRSf5g
IyD7i+Ep4RgOd2qPZhZtHxHVLkmFQ+x2PHvRQlDIVkB8PYpZo9gyx9tbwHWet2tXYwjDJLroe/vj
EZyTd37Wg5gHCrUA2V3oFykaZSdDqdQjZEyMqFF42rvisqq5Iy3ZGM+y4ezDdwlTcRZIsyMYQavv
q2TNfKPbdzwDtfQlylW2fT3rECWq4FZ84ON60gAjJCgvxQ/Stkrtw4kFDTyXq53WOv0P0Ozp5G0R
/qSkxm1iBvGQY4pbCdEWoIL1dkEg5lAY6/izTSCq4jhUMEpQokoM//3YSLGEkAVggyiu6yoZjfUN
O2q4WoevN1pxEGNB7NBbpyoyFD2yc/D/dR89BOdjnpCjp/2Zm3yCjabockNDF4z9zRX+rVrjjQXS
osH8o6DP1dIVNaXvdmBeTB+Z95+nXFbJCq3qSlXAtTARixGYg4rMMKWGNPOc91Z5n0eInOqdT3ak
Nh9D/215WxT8Rrfif2kJt7KQrUVFAtfLUQvZfQU6187mEknABcJfuoi1eLZPR8n21DsTrAl8SqF8
6j7rAPb3gWjX9V+hBNxG/wggOU0zQTPb4DX2MQ4KHfCqCC/PPf+32UFK8jkdEOfHYwcJREAGQOdn
lvWFkyvu6dBJE5DjrbMIVueYrl7KgG+4a/eVi3U90VA0M/GZq1hiS3oH+qOx9lsxq6i1PK6uxuHv
GVhzcVleidenC4jePGkHfBQDj4k2pDTkda2oyJyKY2mm77g+jKumeUiifdL+t016JzqvArUd/hhz
vQ6t7x4G2AVEgqC3owklxLfw/ZcKWDLcM8JhuIOcLWDVH9D203PzhZghNOvsHMPw+rBWBCd2FNhK
sKwwGYOp1P4+s/NynKDNgaCSevXgvK0C2jQvWDxoEPf4u0zoPPE282nVWayVsHv2bmlOSZaURhQ1
/+sI3p84CuBGrpr/tJjWatDcuUCerb7LOdAvSV3huHyadAIq7wASnMYId1qb93O3PuFkaCvfqvYR
jHHU/tRk0KLNrMbkBNHUbrTMIZZMBSrvnEXo0pwz9z9gBHELOmED7vyeeHciud+DgiIaTspxDRRS
2ttixtJaMyXQv9aJ98cOadI2vSkI1bwacE6hSATCsXFCBxtXfA7jt3QIheP85rSAiuo1/7jz4rZm
UaGCmaljlbqvPVoQLRqAa1by67KtLQ7PHaCG2kUzEZ14lXLnvp4m/uH1TAyuSaDjXSTYGVpqINeP
9eOwUm0FDL4zVlHTQFv1KpuC4T5DP/4Lsay2P+/MbgRgayqo43ISZzTpV+GXsVWaVUdWgvURnIQm
R9FDjTXNEj92XFrlwqybi6p3rdea5Zq+JArDj70vr2BGDUiz97mkOyq9FHbWlf6QSHtKvGFdewiy
Na+tKBDAngsvHvuhWtY9Yrjp0TY2QeLQYSIaSO0zAJ8Te3y8JIFs8e/5EF0oYHH3LnmXb0kPrk+3
efsgK0tm08qJ9iwF6B/sEP5y7L3RLMzb1CiPyoGqKAJ/pZvuEeBvnOFtfnIEhDriNntLCeLWpjqi
WDY+WW9qXBNvrpFpsk88TfcGUCU5wJOs2WbRhk4GW3Oyo41aNxoSg8fwy6heEupxgog0KYvxEIu5
CQLDc7y2wF5ckeQX2syIIUfQPUu+Q3AOysg1CXAGlf9k/qi6+MUqGyt7HZ6IfMmVipNZsyIZbGsd
37nwjCFjcCfuJFAX/WOb+HSW8GaBJ34tPj6AuXR/w1gq/ph7vKXjvvSb8qwkBE/EAw1OK86oc35A
VlPqA2uIK0zLO11uJQfiqKNWCiNBytnNjzCl/PPjpb2YxYzuna3JA7TDQdy+HpCVRCQM0L9w/RW2
eognjddEEr74gvgXQREOI3yhRxj/BoRsv1nPAY9FkB6OT3s3HMvuz+g5VifSpU+VufnAaDKiQOY0
nkw6ar4ag0l5lNQ3R1TzSDzyapsq9eUJCK3K3CvLP8CJQEaGA7httb0wmfw4dJ4zjk8jeBh4UUvD
r1FH95C+H+3RaM03OHp+vqGP9SAxFHa/qWe+2fM6dOF3Npvw6zLt/8PyuG1JGnkH/9Ye1MpWUJgx
DVUKuFCMlif/t1ungUi+W4LZ+TpQrifcceOpNNt1ceZpolzWgU9YCcpOVfRGtNTGRyb64Tgy/izs
k1HUgyM2X1QWBw0zOt7ABhZoz4450L5GOGxfHb+BJmytH5JJwKNvouwjpYDok9gn28ddhbDIfByo
ZEsaLf9fQ4UQodcUh2T7guVRPABtqeO78uouwtSYAoI0GKcha/OkanGLJibqxKV6dwDI77+0EtW1
Md8hgHlpRybVhrz1rmBRNm/YMbku3wd/aaWHDHY6uOPPe69wuNDPOicqD9n0A0Kroj3bCrGjywnE
rE0jYddtl/8lPbA62cdE6ZyniEPwd5TCG3zG8qzWSLC5giphekszc74zFIP0/JR3RhuVS2xZq5wv
ELdP0EN2E7ipBmNgFSLTqLZe11atxKUHuzFvMcHBJXNTOHBNefEVLi4DJsEv+IkAAJYCLZPwM2ly
u1+xPrZs4G990Mq55uQfa+LPnjKtv0QZj7EjiJ7MUAKNBjye23CWeUKAspSkIJ3QSUmcYTlex53+
Qpvhlscwn8s6dCVpTsrSVA9wDaGgm4QgMeNHS8WBwP+V/pqy2MXruSo8IOj/FJG/y/AVkL6C2STU
ry2hiMZGb5UmEQSbaZCx+LhDCTB+T2/sQgiufNntd5vgyNOvj3YLP2WQB99g2Ym2Zlr6c9j6Z/mo
Om3Sy9nasFnRWeyId+HJ5JFahL3EvjNwT8kxGpoJTB+LIdIl9TExV0ux3ZjQ98ZGEUOT0BTs1wMi
Knt7o7+J+PwW1jYtl/hcrb5LaJxa708mThHFWLTQMfePh6ZNtnnJC2Fj5abM4ZZxEKNji8K3FbaS
JqXFX/gVUX28afmZsZ6dw3A0W6jXQd+gVgSO9XJu+yC5GqpSaLw+FUhIxCCrE8QP1S4/qFje5Dtk
R9WkvH54ahv74Dp0t6Lev2mu9+dKLveMN/Efiq7KbipCrmmOjymO1YKLdGqt4HSd6DlU6fobUhLA
QTOqRrXmzCNqx8p1QKaV/2lmruB9NaQUflPYyGJwVpE5hkAFzM2hmkAoauPhjtZ5VxzC5MJCPe85
CO3tbx2t9s5jCTTPvI0HiXrPDQGuJDljGSvePmIXWfgrKfonsBpY/xzsMaDotB7IPsFHzhKNcsdL
m+UWBfT5zPCaRCvlCRZVnhNQyFYF8Q3+7iqvmgfYeOwy+47CcBRyat0zaWhn0Iy0U5hhaTNRp0lC
mxiTaTNvbs95jJ3Fl4bOXqXMKQ9HEec9U73sTgnbiuv8SAhBCQZUFceuTNYuYPSQctIyhJKri5RR
oB9zWMClIKo6+/j4khTqqYflKAI8GMC9+1NNMN2+AdHCA0L1BbhZA27JXz3iqKilmtij5486DLva
3zVZvRd0c7Kp5/t7aY3z8pZ3N4TyS0haOvDvhsQI7PT48Bh++dyx2QeXk4/wJsQLh2zqp9DZafq7
3nK7gma7NorUjeT8CHfk29Oj5EWLkvQUawoNkV9tHiO70SV45YykaK0Q7/Rr2WDbNFq4zOx1OSqo
S7ZvoOCjgAlEERCcH9nzt2szQnUjquIrhKNth1Q19+J6OBTKugs278YXFqeBzAlptF+BwlLrSmJg
9y1IeW5GHeXw9YM7yTKUp3ISg4SIfM/NS3UYKVOwveLo/t43NUFHqESpIiVM0AjfbhWWG3RftGjx
snpq7Z9FYT0DRth4AKNGpddQmgX+FmUIgFTyrcpQwmP9xafrsA7b1PVaHOvQxlmHtsUXiLXyYo7X
IwtqQXRN5tycgyrtDITvWb/hYKqEiq6Ebjatv9veSf57jQnQ/Hfqnr84USayV/J1jawts7Yon7p2
2qQebkFjx0Rz4plovvBhvTg+fwklPTjas0etFCKkAmbop+WNsf+N8vJFNX89hXPkEXzr7MGwhE15
k40U2eO+6SZVjTXq0eDYuF/uoXEJbmCUVd+3AeKjqP0t6l/WFKxan/Iu6RF4tonlgQNMMpH5vTr8
Qr9T++SsqjqX6at85XNVfOAOa3UAx5weZ0jkLaXiNnm0lV1QkhLCDZ1D4F+AkMvrbddLXhBMjgZA
olkKBz0eTtHT3EpkYYNA66tuVjtwbFxS7B4udz4towqlRQHL2mrWLAd1jCQvQcWp60NRS9BvmIS9
NVg0ZaZo/otia2g3kqWSGBf/ztruWPOM6dcx8hs+V/Pv+kg1qGlXJ6q5DdgCJz1ZY1G1xbR2STkX
k8LopVRtHP1HoLIe/4Z4hSlGwkD2dcO9jDzjfy1lNlICnu5NR1Ix+tVo2l+BvzKJkxmcmmGwyJnM
iPyn90Ow92jeZTwO+nFD1vEqMOjciHMrpzzoX1CwU6hH1Gq0fjxFmKqzeC5dAM43iOIfTMU/IUtr
ubHacwvyD7zvYeZi5te8jlXh4ykDYW/Sdjr/zupVzQqaI3T5ntXgunc1hpS192gv2I0NrCgEdAaw
SlO+ptQIQ+DXAry44v5ik3tIO5JHwNL9cZ1LB4ML8IlJjmsVvc9gYcrqcyl/c3jw6WIl5lXNMEM9
uec3+7CoFOe9hp8RYEamzpYkrZ5lV+Mx6+6mo5m7UXe3E3gayhbXzDZqAM/xNHaf3BME+qUb/gXT
u53wcN1EyDztCupdhmVA5qJjjzM/AUF4Q5jZfoJ3Yh17LBLqZtsgV7xkyQi8YfJr3IRxTHLFI1uB
PE8JZDoKbF94+cU7OmjtSqAKx8bvAt4pVtjBjAk+s/LO09rBLKiwf6nUO827Qjtt4zw/Q5fMS3F4
pdIOSdPPd96UvvCM3b9i+nUopTnmvMK6PjpOS3G4aEuQjIQ9ts6IYwr6vF+ON34o5y2dBgy+ir3h
NmcG6V9NZIB8eAfw9568ZnZ8dPzXNDUfNkQ/y8/f3ql6gWKN2oY3lmEIp1WGSsp3gll8MK7Hxhd+
H4GLG26JmbHHFNgXVAbB+fZLMH32/C6kDuITEvCYkAeQedBo0YweaoBa4VvbOPcU8vJ7BxM8hKAa
tj2eSXaWVYZ7rPphq2YXrXPlaqfEpkuih+LEJENo6TJeLQamB1GwSrzL1IdvWoYCpXDy06nXT5Uu
4fI9Ngtt7iSH+ivNWtJmhrcEhEKRipc9sWHnI2VLgVnYrDTYXNuYRXNwx0KrkImk6kRBUpxVN6P6
LzFYwgMHRreSJ6+tQaUsIaw3MIYkyTkF8cqQpqHLXSK78wN1QakQ9fRMctZ7S0SQXCHV/YcOAKEP
cSv7aXQHZ7PzQZdeftutEIQPeeawCepXZPSkzLPD/k2hsqSfmUlt/YW35hGcqCdpAqXcHynvDSJ+
iVR2NonrBQr7ttJI7MSVV1TH8V6O6Mh0AyoRX/gfJKU6ZC4boCAWqTzKuNrhOeOuoqSUqxHqca3a
awUPwPex/gdaRgY02zu+FpaQv28I5eamJxG813QGWuoRJHdUGah1+/t7mcP5DNWV1T8+XwWYk87j
gQgFcjxjkweid/MgzIpSdwUbchCIl3B4Yd66QpLKM0/BCRC4XFGTKPBXqcZLxMQB59SkqEtGXkCY
QYqsEHQtygMf4vPDNq2hzV/ZcixtLFqeD8pZ2StLSa0N2lpArVo5NADVLTxDmq24oEgSWe7pVGJT
4PrslVc0gke8wQJf+L4vMwqZhwJcMzYrkynrbowblqN3arBtqx3q5SWTIayk+ogq4jx/Bz5vai4T
fplqk3ljagLsINn4bPnmEji8q5/iOBlNcH3jkDiea+ERspvDpm5NJba8xKVGeleNPMTLGAlwFoLf
G+Fvp+zNTkgYEgvFGPHoSJI99K3Ficp/HxIrkZFDOoq14q2A+h1LujrIcrBRq0RaCV8TemYKtq7J
FfLlIGcEbX0L2rtv5bn3s4wsYPD4x26AOH2ur5NYFnkSW2isk6UTPm77Z7WktXjyFFFQt2TpsMuq
hpT/yo7RsimdVqe06Wi3YK4xi7w3zF6vUXhAYB5LRMdr9EN9n+iKN4/WMP2Zkfe31b+NFJV2ezD+
4ti/aJWYWqFhMHT2rXJAnCdZZyLEsqjioxufBbVHCIoF+aCLyVS3Cp/tzWHmWufFJSyCa+K01M9D
iyomYsozl/bNeV+2LEbafkRMCLZ6hw2FCynNm/FS6p3ZKpJPHZnjhtxJT/p36GejWT331TCFFGR4
d1Kr7PkfzNPKPDIjdyQx1aKS2R5WCRsotbb5L+pkod7sO+BdDgPyOKv7mOW9Jp1PrVuqZ5FPRCUE
PBhMKVJ+CcudzIfKznnxc1kQF4HkElPxNGGyHira+UB6VR4R6C/7oMhZhfvxLIScbDAgAln9kzgn
VoGTouGNyPbb+igNhe5brK1A/nHLJlkWUKB0ZKn2BIph19AW5sv9EWVVZ+2Y4itAKsL/cRmGV8uH
DG1avyGyplvcuxMpnSrT5MLUeT9svJeY8V0JuSij/YlZWpvC2f2HThDX7jMblRLtUmRzcddJECcF
KUwDCzQ/JOjMmgCc2TWQJ/yvHXciWfCJLrqZsoMLxs6jpLmaIZvYiByeCWovcs/ddOas7e9eHHYf
bASufkV7QwW+ZJTk3s2Tg/mnGtS62sATpF64dadQs8XuEVEEvJ8s1Qy+V6eotN/kvSTW3ygzRZ0h
bKciGNES/oBX5agWig1Mb7jympMxwNinn7OgjaYLv+D4LtUX0blodK9AHSMrKdZdqDzGnKwmF3W8
hvFJpRqml9llAoYQJ9z/8tB9GpfC8SiTAigc8ac41Qs7ET6Lt84n3jVvLVYigfTqL+G1pGkdtTAM
eVs53NYdXaefyxSd4gGQi5AUqRWyy7NUPlCgotLdkJlZePB8/SPhgGtN19SrVyiLoY6I1pJnG+xM
iJktE6K2RqJWlueaLdr4wwVX5WUxPfte+f/G3Ax/LVrCsiR0249Hk6Kj/AlM5r9bSu4pvydpHwmY
msz+gbRVRYXEVJW49GDrWiHXcpfkpKsw0CfKVZqA6aTZIrD61b4hO2S54T0/kFomh/4Dm7g+QGpD
enBvRLkDZOoHV7pdz8zC5vdCCl78kZ07/ipPo1pz6MzlXmCDzok0JV6Ei/3g6p40urYp3Fufs6Wb
UXoAY0RN56WgG504PK8eiyC6nn6kT0IwomYiZhTxfrxOfVD1GvNWNeD4Q5JBhfXJJd+9VYGo9PKI
kAh0NHr/Flimb1msQQBqYWtSxsnu78vUd/vnzEQfFdEUFz+MQHSLlgekjt4X7tIHIRPv1F5HpBTx
iwKcxvZLriZJB1QDOY6auGi7PmvCjOTxN+ibbvj6Ho6fn5BPzxvQMTkCpzG8k9oydmwWQsnCIS7q
za11/mlRTPfX97mQ4sBlZgl+NNIlK0XCmb1POTYf7hGttmZsK5TkTQ0NaKDUb9EgWOxf/l6VQpks
QKNCF1zbFwUE6pb+TQA1Ja98k1dbLZX6vw8yjD27h+a/pGk7oC6pUIMVyphsZEKQWNI8AzX+/kud
Q8Ac2JJDx/7iZ37Gz85WVwhincP6AaUQnCmCETyxIlhNNFXDJ8iPjds4ta9ergkQx8mDJccqcNv9
zuVyTIIwDfz2gyB1UO2deXudvD+XWCruvIgUmPFL/mD+I959Ub6j2xFAKd2CoIYQCLHJBKWQNjL2
cyXSCrdldEf8345VVsPHVv+t2JHuKX39zimfSsEccS12JzvT3GlZt95x9XESwqIXcBSam6/BQRk2
BE9+tRE1VXOzyICrMrEj0QaXVZrL1RQfepk43eqHpcoPgsbtA4wm4AvFVMnvNsEhCXwvbolN1nKJ
lVLHiTKCm7xHV48iC3ivtRj+LTwEpTHMpzC/8P4lBNwz9VIanDnNmwP7Ii0Zok9DJCN1Jmnj7Zqw
BeW4B7oVXx/IzNvjQQL0n/+YeBhztVwMB9+CdQ6pxgqPxJJb2jwAoVrXkijjAhdKC7qeMJUpqc0G
7gycDNbwQ9lByyS2rxAhYdbmn+4mvWBALOzVOWCH18XUxow7XmFBtUoi98hwm/tpJiWJMfDt/4ni
gaXHFM+Mu/K6VXFIfZWIJ9+/rZ+Fyp8DR1TjXD2IFsJwQgV+2kb4D4v83EonV9PVw9ABQW79HiLw
3kIJVvetofFmgsx/SRxdL15XgvC3y8/ZHOl2HQaa0HYjIJk0vg75b1JjHesHu93TpQoQHU+NC6of
8ZVesOvS/67L/lR3DrOU8uSmh9+ocu15HEJVkQigzLtPatqg6KJ2ukwdilU8ZDJ6LYGaHkoUqeKs
W7xsX9wHDeAYSeE7B+rLkkBRNJE/y9pEh1JrvrAKuLacxtmxomiTnCHkNLY1ycqS6+Iln8FmIHFb
hbonTbmZ+2ZIdqUUnRmvyGA9IDcJ441m6+HLVapmr/GIeC7Rc67AVPTAxYjPerQAdgBlyhX2MtQ3
y4LelOPn1ddR9+AwbXvtUyGNyoC6yUmBqnXESWmYnn/foDpiJWtC7RAA8gXtd28xwXSVEJ9RMJ72
dPe03xMa+iMxCsJVUbcXGMLyJLFUrRbW/JN816uwZ/Sbubz+kXf6b+b8pN4s0DmoMP1QMEkZ9/G6
XPHgQsd1XT7w/QQKZWhsktUhn1agbHd45itkIQ8SWnsdW8AO6yQUHxmtW7tY4iWha6uNiQH/KVPm
8BM87mW4GZRBU/D+haBvGir3y97g7CFWLFxM3vj69Juf49oiBXjaDtrhG6q2h7rK5XnTTBNsxRpW
t9eyv81+n4wk75fNsCGg8JQJSntGaWA5UJeB1P1CruHZl3G26HLdyHBAVjcrfMks/uDLiK2Jf7/t
wcgr45+UXV3sY+1m3ReVY1Kac3mv4/g7fr1Slgn+2lOA1Y9SVixcjpBWLPgcDVgMXSDYJ3qUbdg0
2C7OWQtRXLsvRmVfgi2iNYD04PM/elRdVFiMfwG6OpmKSUVH+YqHQHpAaR0YlrpaqISnwoKQj4bN
4MXj2NgobsB6TlCthnlWjorRn6QmeafvF/Hq6wM9Sx8IQlH/hIcCQKY1XaaotK1gWi0vziuTh67w
ebr/ZcFrk//kzL8j48/WYmX8nqpOZ0onS+JOREpb+aWloQBguxJz4pDpDrZP20fTViVi+2PIIx0S
W2lMfd9GHaTyQ5HfnSTx0KgssjE31GqNJgnABaWoGMNFr4g+DhZTIunfnu/SpB23nf1tpXhvLymQ
DM8B3v0bzcmjF3BVrn4DmjB7ITvouSJBUvIwJePXAfB5fYgw6U3e6Xn1ycM0vcLkFzXup0GzJ7O+
2TtKtbAgPZFdxYmH0RyrZy4kjyRCc8NssfZLcKreSPrn9Bg2u7Gn5M/6HZvVpBnpSBA0pQ018OEv
6D2y2VaY4lB3acY7Z5gKzhMbrXyC+slrd8EocBgSmXiMCG7ZRBvvUf0LdGDWOGvs//FGRkRjZFz2
C/NlqJ/MyA8G1itKMVeGsAGIA9tLIUBt6bftAuhk679FRu7PRes7gS8c8H5MgU6N58WdhZsAHOta
EmwWQ9wnUQeJRFrVrHQQvmDw8L9bNGzHh/AgiEDDTBPPF2HE3r8m4kJLY85jR0naQBvEHttsI6Dp
4cEEo4xFptBq38RhyuLqcM8uw0OTU0szOBWfCaJdhUyVPPz+q7WKmNyvZ25S5PtIr9LyzEWOiXuF
+1iuP4lxyfXDjTWfKv8FrNEFiD3JEh/1PWvslpOPMn/rq2fKF6FCJR8ZjH33UnZ6+6hqV6mCSRsj
7XBV/lh1WUsu4MTcHl0Jy0suH661q/Li2ULMqHq52K4fYo6gZecfw4FbyAlQ5AA6C4OB/zqpjEzz
lykY2Sg8FrlE0+teY6bJ6URMbNBdd7W2ZfxYKKdkKFSyqA1OPwr1mgXzAYNEKI8nveFe+9lIu+hH
m9IDGWHKLzw5POy6gUJpeBnb0B0RTRPoDtMfsvRcilmEkCMCD4Y578jL/f0p4DbaTTPQhgKK6lDl
oTDS9u7klrvU92AuDP5fUg6W2CtbKX75lq58IGZv9ktrRKNxSrV9OHV1vLjHx6eFjfjqbBpTi8ni
t14ZFfyca4mVmD8QVIAjOr6FPx7fj4el9e/DZESPM4kzbuAD/m2bjjmRsjKDyWS2rP0a7q5xXbHn
SVu0dxSuYRVHoziGSJ++m+lv77WvjXFR6oJdRn1dO72kNmvxYEBF7MdzHy963msKZ35BCV/hoYmC
jYKvilbopDZKnN/nNiE+JKfLrxCUFRbVn/XdA4FuTlUcMlV/xP8yk9Qolv6asKhNsR06yeEfJ1BX
6qlNiSg4jbLGVwLWP2J4uxa5nE3XTpCZEKTvCj+2yRImdF1g+PjO7b/zNpYBx4M4v/6+io7gu6Yf
l+siQDMWy0g7vLqLlsBQPbzzVqqjjRRS7SDxplF5gekWhiDKKhEec9c7Wq2h1cx8zppjuxI3FAVa
bsP5EFidHG7wdnbO4FMLye588F3XMNJUghXMEwBFxgxRotA6v7aJ4u5wchk0NERe3m1lML9zO2lT
HVr18peHrbL1E9/wr288Q1Yh3//gFCpAfhqKTpoyJzCeDGS09onWxdzldQFwFiceCC9VI+ysc/hd
v1E0SaDGJlOVTeqCF/XJM6OEAqPjvIEcqaeCRR1k4Z8dE+zu9yTJOt45V5En2rmKPyaA4DLg0BaL
x5DXQJi5cL8dur3ZLWDNwJaLCiVVe1kZ+e6LWuR1FeN9DVi0Tj2EfGK9bwkJhQMvgw8DeDQndpJ/
wluSyRHL47Ytb/kaaQI2LooVoUS3oa3b3WKEpl7J7+CbER/cir6VABx7GMPFISvSmq1N5hf8EXmB
GrWXZKGmyxoX3cUk4bknSNu+6T24aoBJ92uWjfbUN7FJ4z+YV17wd5CpxnQ4axzWinqDMQfvqqK0
Eb++V0JO/gO/b+yjD6k8UarFadgXXBtFZE92tLwBdef9qpMkdVR/IPe5nuMwGkddIKVGr8+3eDqZ
vlR4+cWLfAEM3VbsdUCqtmdYg/+IM4i73oo26rU8Inq+8SwFvVNRWc2pVfKjOg36T4JqDSkFV786
DLY9Sw5Ft/chv3RTcMZ8sb/5xA87iZYfYNvcXRFFZbOM7S7a87kKtBk5zeKVn6/9b7ES+yoGq2vP
tQs5LoCtAJablKwI0fUEGs+DIVQoSmmJW9os2qCRQpsNNgTD1qkuS6ayJ66o7lMJ81gJyDrRKQZk
Qg/SQelZgOQIQBemAcaK1JW6QRvo8bcgEm55jtvNtF75n5tWZiFGMZx9BMc+jbU3McHAkpIvTpWB
jSYDQnznW+JqRuJKrAWnYZQikbJjeoZ5UVMY8F94ppCN/Bo8Ah2eZtRGsxIs6BMHFtK8+z/GCV59
Ncc7a2e17DhgyW7WKucIvqVnSGKO464bH9JtSKoUOD0YTTo4fPhRS5JdXYK3s5XxeNvjIoWNjL1M
NLgSkZ/0TXZV6AznqcDpORY3HFxzLSOmOH4AAzkOP+0dbzVKQsNrPDyI6RZPqzzo/hS2X4LMR4Af
Y8BVJuUIzia/6O9sLer9FDTJpc4LgBnhtROMn0If8EnI7JtbBaCa25B4r5IK/o7ahbS3/KjRURAu
Ta3PQxoKcH9CcxWhyVSFjNZHu6GZWPc1v+igxMpTKE8Jp3fDN0XXH21LRAC8vdA68zw5YDO2fM20
q9qVppKiXk5BI8t2OgO9hXPencIYCrUTNoq3iU+/FbNwBtW8LSvsJ3dHm4bjWVTJDL8H0z6hJdR9
uY/Wc8QKf+sKJOv6cZua+pyd7UbVi9fK2EYENiCQOt/8sfVa+4NvQ8B+l654rj37XSYw1gfyzm31
msCotYvwlnNdlORHIfDOODNxZ3ee6iHFUeT6AasRhuUaIDaLcM/fJvpbHGsUhwvTrZzYpLhTrale
1GCotNWATIePuAtcj/CMAYiBmViNJT5zYOch6CoUwJzZOQBH+SE2XisjzT7h3vH4P0IgaT9trEIZ
Y9Df5Kowx7aorqljhG/dLdV6Xoa/YNR4TrAtceTvSOMTFKgXhpojELhAdFwB0Twsx2COn81rY5n3
pO36dePPSbK/Y5cBNlzbh4BK8ITGAD2ZzQ31gcGxENo8LfIU2/T2b1eWUsHkFyGzG2MYsfeAJY1l
GoCTwwC+Jx4w17FOZ2JR/pufkWJLwebudueUEyfqNTUuUZsjvVP+oar//GDq8lM8HvnmMI3XSdtv
L1NXNzmCdkWk/56By4wfi5ib2tzxwYJS0vtTWhz/BK0/Se1tSsfnNcg9dEFe4fIoPqh5JQFfWin+
Jz84DD0yX8Ck5S5T7PnQofYoiQpLZL0nsb8H36r2OJjWxztVYMolb+5JdPZF4EhRoB/1RhXEhnCG
FxR/3NzRb0rnw6kytYyij//WcMwNdQ52Qpb6NKuwvzZqLNFGz0Anaydd6SI9ztj+3wyWEIpGod2B
1aNcF/z3X72jSl0q71GPL+N3f/v8o83ZByVns8U9CZSP0yIiRn/67sO6dlI9Pzds1ejI1qFecYJz
Pwkb2XphZU0VK4w8QBo8Cc2SA9DkOXv4ddSamW3db7YuBzbWlTZPJHI1FFOU+zUNQxUTLaZNj3bm
t2zRUgMCe8OEWt40L4pw5fs8dN6mdVmqLjI7nyP6frvMbxq6jMmP6z+5OSZ2t6QXUPabaWe7PTlN
EE8Ozi4khC2NdFbMs1oxcRTxIuArTQtfjgytp7QnP4wUsCvEDvdfaMFiS3uwxQWAvBqm/30cHzfh
ev9LWK8dIFtGjwgBnGipoHfxSm06vtAYuujRovy0SYLlO0Mh3UOOaQcOUKxAEfS4z7iPF958vPBs
LbY8OuLVka2R3yLf/Nw73F6pQcd8A4eoz2znYBNGihcB0hUkQNEzj4r/gyBYlj4wpB+UggVXEV+L
vNHPnctFz/iX8ptFREh0/11v19AmoRcyduXuWjgnxauhHwDGag4HukpLWMv61sxl0Ot1ZbGAvSY5
zFzReAMYkv8mgrebIbBuhSXp/z3c15ov4+SZzQoZqQ/M8HAwAGUNGc9wUko66CwncIVfpwNTrBvM
MI0VGOvy4cVKX/g8Li16ab+q2l5CD3bIGryaHQRg3MQt/bhFQpFMV6IZvEw8SFtA0XZRpez22Lnt
3pbEQk9JRUCDDe6aPB/cnItG477WMfN9hywi9N0MZUfPk/Uw5PRRVWaUwb+6dhShoypU1p5t8dR/
c1h0IA6+IZN8+NQqL/13g+8uicxUFZh02SB6ZzhKQNhld9h0VZ+tTuug5EMbEaaaWTfj9mu4Tqho
suzqKWOQP11ZAE0joRtCJMhc0KZEXh1NN1Km8OGNk13Pgny8hfO5fx8Pr5dj1LFeUp9xv850jZu4
Q2Dvqrf5MAfGSuMdw1tIp5AybmWEbyHg6eekB5qsvldrf/nV6FhvSxe+FbyOErWlgqjMlISV+CUZ
r4hvI3kZFHrGatqrhiwg+9sXhcvvrvG5wcQHPFar/QXexi4RP0ERCtHjNQ8SDfIIR+sASAludA0m
J5Ze2b5IfYT1mlctqb1y1W0mnIrVg89b3chLNxTnaWXgscMheFgmPQseeo1RQ6MZfKiyNMLRW0jd
Ggk0WrIZlWQRQsfzLNF8i0NsJ5Xuuak4WnpFTdoScR+o1S0Z9jeTMquOQ5bgR99msn/HjTpXzwPW
bJ3dPPsVcgJU7nFUnsNv4aWlOxkH44sb7f/enmcVmus15MLjP0ZdoLS2Yxq2zx9gdZMjjAVBFaUH
v/DIoOU0mn1VPHAEkgGX05qGPyoLcOmzo2wgj2XqFqk955J+E1bkNmXeRuo8/TeAHjU73WyNnAlA
h+tERnzVYlLshNRnRyx3Ov2AcjKLkGbSw/hzOCXQbcDtjkArBHcN1B+Vv1uPZpIpPKooDVUlhtpx
DqNhE5/vZuxEYIgvbOWoaNcFptrINZiabXK/33DwWhWgQ2EuEEVENOCqCmi4WM/OBAUVCUGAmpP4
ZNw9yauUWU0NBatRhkJiTOcedJ2oyjaIJhFeK21eH0AejpigG9xRi3p81B351KZX1R6D9K1Xc+ex
Yy4BLlDkxaYJ9i1UO5Udo3VToMpno9UbmDmsvkp11ZX+MSqbOkG0mFn53cIpW73czI/24Vv2H/2K
6Q/e97u0TwqkKRAqlGwj++HGEtRoQ/oRQnoke5yrajTbls5HFwpGxTW5qF3p4XecFSLJm7DDzDPo
bPBYD+IfYjtsPcOonAz94Jm49FG9wrKqmBqXSQg6MZ03YEdpe13r0B0aihX09i7oyasxHKYLHzUM
TJij3l7olz30B9QbhNdyt/Z9h5su6cozO+p6+6gAya59jKn11Jc+vWW8HEB/gIpWDi1oOJyTh0YM
NwDCr/R/HCmVIXJNmnlBUCm59afrBz6haSRGu26S3iiouKzIA2hP2hAiq/aAt0aG94GAYwieAUn9
cTfHln6VsEew7vqM/cRiwqRPRfeV6rpQ1TOPUqhhfHVHx3TMd+XA5yWSTfz3l4mEYPAZPfbrCL+j
yZ186dh2AeEiWVSIXUnHGMJyHAXtTpw/c6IWEfKyg27rXK2dBsnkCn5lgtFwAD79fWDlBGpYs2dj
dPbzsAfiBIRp/skooq4N0I+qlVjyLq/ZJYokloYBXMViKv/XxWTMk0OJmYanGIq55GccAVn+IYpO
lKDl3T2iFXuqRdhPwH3Eiw4r9HHqEnJESKlLkzbZgVphsFcEWN/jjZr0SBa2lYUyL66PBqR70ah9
3OWbk/x3ivrxTeDtZo43u5L7bbOHW4csmU3MwwlSo87LLhm9054G6uOOlXkwSmV41KAdwIdpdccZ
HrAkEQE8k1CgFeVI15il+3jSs9zy02zyI8Dmo9QvXRwx6Zy88Iipc978HYvJMDwVQWNSIG5i/Jaq
Gto28LQDkOXlFUikisFUYMKWPX5PTFz4kOCO6FduNv4dCtGs+n7X6F6tmwi1+Db+dFF1WIPxD6oF
kP0LyfWI/Y3gkOEJ8G7rF+dc0XiLn+AQpbZrl7RXqaD8chCofqZcCpTsZCpthzX2F5yBRZliyLcd
xWxEw2HW9gtwDKzY4BTNfVSMchEEjn1pCu7U0x3tPF4F2XQnu435rQSOL2/IHMlkq0LKs+dQ/h17
uBQ8L7kkF8cysXhdzsV5+pBhFT9UmPB9Nq7SS0SLnePWDLJX5ii+Oe1qTgKbsxazq2QquYeKzdRa
q8yJUCe5vwchJpVjCYzbXgCiZVC7o9lRnlUteh9IiWi0h6f1D4NzJeO/COSvBA9jpoyo9kfQeF78
7E3W8z97Dfrj1pqsdEjd4p3EEa59+5adIPOw0rSdH0i6XSO9tJD0QhQWbl045a0GVMdqXKtKuTQV
48u+ednqeM5JxOY9AfV+MlUrlg5f4Cq8r87j/pOkXp6K4XcsCRLLicleRAfr5RPZgT0LJmhrbR6U
y5V0g3pPmI+lB6xzyldMn5Y7NZd+SNjSZ4CWkpNK6e9LUU+n3Mf3MoR413eZlxEeFje8+zJo79YG
CQuEkRbeTbvIGd/9+Z1B2R30aKVrZVwU1iTjCYhf8bhzhb/CyFBYbWITI9n1xPRgFB9wB34JLUgy
KyZujYqj5MeaPNatBmz0gTim7fp7wW1zYK2QHNWRVz9IIyZ1Z5323UzILhDO2Urn8inRRyAF9x3c
aYDlG2yweuLYNxrGiGytp3u7uOzywewJxrUu1F0QzZAe7SqVjGra71MlWRejXaPxQ6ttlXXFBIkq
wLAuXDtJWoxX90qruMyhD7sBCqAnOut6vioTUPSfhDQiw2jhMW/Am59TTQWxm7rmf53Gw280sTnE
uABkNeYT2t4o08dwwHSe/6Neu3pw91w2tab/vlvYbtuEEUKCh/OC1WXAG/insOq0qq+GfvtIkvdz
0jQenbxW7ntamDCHnQBNTWilXLPqfmKVRvO/h3yHnNlWoYSnWzgqHaH/841Z1pqH0wSl1HoqYbir
cKJ8dQhcujd6bmenimNLNSSu8tjtAOv12qiJoI0FkAn3GMyX5ZE5XOApoSaoROzwpe95vMFyx+ve
wGY+YtNHtVh9+1P73GBudbI/Mw6LndbCJ8eper/6UGUbZm1FhGuLr77+GEspLQ1iIerAMXTlbUF6
ErYl1ZQJiVGOJIahQhLdpmGNUKBpWTpmvtfDfflhgCTbGM8T4qSnEm0v3H3/joqvCJiCKfJ36UiE
+td9zGuILqioKBNOj1CQ5dWKpSVlEsGjz4EsLgioBRpy1hCx3BEatv8wN3vPyL9r1Im17c3GZ/lQ
kdBlYHg/m+qFwjzWvDz8sy99vgOeCnJA2OTOc1CowW7YN/fWXj0gWSxkBoVef68CdsXTQ+an57A8
N/SnEi6MdFZsB2Gxl6PyiFSkkDtEyBdZukbvkzdph0E9BmPU0L2Fp7kvbeGxdTVaOC61zY3jmF8V
GDtobSRV/ep3yt8lOUBDlFIwE8MMxBiKLRvWccvjJ6Rnxpm6KtZ+YFcuR8cyBbtX++eYmuRqEHqp
EVJesyJXSgRtTA3v2/WTIqQahvj34kuHb5snTCk2X87reCA9+22hqIvJVzvfr2DwjxVyldNQueWk
KL4J9SXR7e1icnmXo2KocCBA6833w2NMHPVR4d5AwkRHg886gOHD+tSclzghpBtlZqQ45KQ9b5WV
C9xwNOTrVMExHwv9RNYVlrj61UsUsBooEjElyf/QMTE4M5mBOgiQNCcRjjqWexdCsgXDsADhdm1w
WKprYqw7kuXJfIeqcrXHS3orp8WME/rn93okyOU5ar+sjzizYNlMsWG5y5uiXytuYEF2rqfWYtfZ
gGi3kBJsSZaJsM19UcYGub8W/kgvaJ5oGAFhG8oHpWxmLtigNMe0lXfyzJmAyxeMwkQgMPizkCgv
oGUzTrlFZvaSGG5ZZINCN5BajAnXRK82Gs4DOdVL7hBoGNkhVjHu7GUE7sApwGivjSyiF2rrMRB9
xPwZAK0YxWQqR5PivsXPfS7Wz881zB3AOMugx2sfY1GWscjGFC57kgAKfJNOqNIFxfhr7Y6uHNRe
3sE+EFN6WhfP43sOKZvqCYC/MUN4VQq37AKnSkrLey2KRLK1NQkChHrf/x2P+t/L1sOoRC5InN+M
WswN561Y8U0xrfiW3NLPCP3n5y1c9S0hLR1Pc9f9Wu3q1uddt9FZxn1GHPBjwC6u5nbVOca554AM
w+/dn0R93kYunV9MqrB94Q2lf2/UtJVcXgVlXur63iOzd4iUqEaY6jP5laBt/EpM4SEsrb8WN8B/
oVpliUan0VTFbO6iyF1DzEwY2XUd0l7z9+ziAwHUMuVgPJqc356NDoDzRkQuDJjISOWt6ohXwlSS
ti9+zuZImQYLC5VETozI5jV62kEpUV8RSdBgF4IRKuEQyxQ0UrkVclteE2/He8uSe1QVBcECQf3M
D7K1CcjnCargdaVDJnY1Gdd7OLj4lfUpsbQ1QG4F+TXv9qzFMjsDEZ6n5o6MyjhaZlg5pprFbDbS
lI71jai9X2fnc2uZaCG9GpBO0Uj5t5M7enMcKUFGgQ0aQc1a06CO2FWnKlUKNb5u5fA+MzQ+bnq9
OuM6JgDNcsLvseqqWzbryMCLvEZvJa44VmswO0AZxtGharPgaXbhiLzOqdFMCmJh/TomEl+ahaQB
yVkWerfHkDEVJFeiKLDASU3WubS/TB3VE7R94qlhsFLM2MitHespuLnVUWrr3sMj20enf+yyx6KO
ileZ+8ZXwVxV1y3puINZ96ZYvoisDJbZdUjqkWhMv+Vo+/ozWti/5fDqBZ6JdmnVjMWtm1fl1D8U
4TUnagxmOCkW8pEQXyozEHGYZd/H16baQDQkKAWE3YKiR8qpXbBSRrjgLVeKpBmPyHIf4UvrQck6
2XhHsSixk+c40lIGCtYfazFZOv0rQCkl6lPLLZhdHbn/HvmRwZtQEse+4xHOCz4Yfew9ztyXnSHw
Efk5rtPb9UZR1OU5nN5xdVCSeixvXoDNRuL76XkDBhyjay0Coo1pXWC264S4yXhH5ivUgkCFIQL2
/jKl6l3c5AXbKA5Y/yYrpsSjTyJuSnsDvBshqQEQzFg6Qx7cx0z48/qXaYWhKSaE8J+jc4JwiRwx
EeOxeb2rtViZIW3UZgt6ufpuQ5Sd5zdjNC5XNkxwwmNPx50uAZxdXqRWMTJchrBawRNQYyd0AdyI
DsykC9xwKekI0qbd4pmlCqbs8cubFzha0sq9ikWTeLoAawegYK2qa4AiiYNLpNODNMOhA2teM4/F
m5+iEQvqmOCwM1K30g4GHMK7LPbVfGJDYtfuQF0x/hz0ezruSNDY+O4wT2UhNmjIKI3EYQg7/lK8
b5Ff9AilSwvDQdI2CZ2CTT5t1Womne4DG4/ncony7VcKnknb/LDTVXl9ihD9T53CbcJy4+f8x+gW
kSBNlZm7qIF/Af3p5V+vvkbA0NJkez7cuYfg7F7JJ2l3myrh52vFzI9cxQS/x+hLHQ8QSNBrPN3+
FXCZOeF4WdnYOU73LA36Ehdd7KIFec+ISUKuN43V9VuEi/HDYqlFv+U3bwjr7kFLKgtux3VfuJ/D
c4KN1ggjJ0BGW+EMywQat9UeZD8xfv6aTwPs9UpI8h2A15W3bGtEWaqcXpLVQYyJwfA+D/tSaZF5
kuXz3rYeNOS2WNJWK1/H5zKnxQsTMCmr7zOzqNBQRy8fZF0OtuWqcGwFfyx03lP26PmsJvZqs/1x
A7r49fQfp/QYGcpouPzNxALdDHvusYrC2IVRR3QjhCL8N/lMScNIAVAdKM5WIzjqPyXHvG7vwz9H
Fhm9NNpjRD+sQQ74s7sYO8Eq7GSbxg1yIAR67QhLVH9YBgmvBH74KJGE+nr0UKX9xNvVZwuih0Jm
BtEJM0bqvt4qhZHn/PuV1yvatl4P+ezc3Aukek1ZpST59hBDjMC7sAP/cAR9E5e9yUG5m08MCqyT
bLroNDKs80USDcz5Mp/8yQpO/9pZFnwhUJIzYQHereA546sWNqJF6LitRHQo/wnH39Q2w3V1zXdy
v7IBciDIfb8EZv7Wn3Qjx8qFr52aWjsCUBg1ChZc1KwG+tw7whLY8RZNIwUEoOt9PEVpMV4/wcso
kfynj7c8hCAdXx4vfGlmo6ZPDF2Q8uNBnx3974C9RFHIcSOtffaPtwRuo1va7VRrh0loLULXR6Jc
BUtsOaTVea7lyirY7g/fRJUuqhCpBQ4otbvBisJ9oag0i5vER5QUmPf6OBcWSTGCZpuJlh1C9cWq
IHq/9syaFD9Xx/EqODSkOyYnaG15y+J7oCdCfLNJdFt9TZljFqSrYMoqFSdQD/xK4kJublAKWpsd
DtlEFX4ioa+M9pAUmQBwQCu4Puaxu5z9htb26L1Zy7BgJUxgWbWqjd96dzNhqfZc9hvze5jhAKse
f64XXExd5OsilZxCeS46wIKP8/flmV4moNfo+0ZesziVuTCr8ya3Lpomq3Hc6HJ1mW6np2UAx+4v
b11Ic67jNAbfRtWqh2XWvXynBH1vt6H1VBJAQZcVxBQkYyaKIjYstFhXvk4zYEKa0yPz0Q/ShzUV
mRGUVTRqNRYp/IBcr2xpNbnCiSCmCarZQswZzssW83WCMvTPFJBlEN1ef5Z+/eDpFePwj28nK0Bj
z3Hn/aUtAQhW9BGEivRO+fXZGCh5vyI5fQRGvHSAb/se7lU7jIuSLeuxTTjxsQGZdo8skDSmlqj9
FUwwQ46x3rEf69NvGUexdc2o414P9rTj8jPcWKIvtkT4OZ34lVc6Szh2qD68uMie78OtybpZIsNs
1zv64kYM984ANwL0GzEtyKT0W1n8yR0ZRQM+k1Y+2e9C4rgp5kqqBvrKXJazMOY0NuSnGkhgV4Oy
x5hlnK3tXo8Y0PPZsrfUZW1A94VT3IxsfOhsczz1ktVewx0poD44gE7li6r/Fkg1UZopTIvkXUda
MAu4AS6deF40P6SuM8OTK3Ssul9h9AePFaJ2jEY0fDDwMofEDT3VjvHcyvS2wW/Bjz6g9qYppeTS
3uMeIeVRFsQUuZH/BZbU8hreUkzriDErYUqDmMMqbCst7nm4iGvkzWf4DMlAvS7ZW+hvYEEiQOJs
SSJN0L3Kyenrpb90R0JpjzNuv4o/HHYNjWgE3S0C+dusw/4kUSC/iTVzHkwOaK5r27qEvg1gIKFV
NnMJO8dguIP2E02pdAqkEIdKFO/4icW7h2xgCIO+kUFLI3WkZnKNCw1e9PPe0r+wWxWPodJuW5g1
Jom8xvhSXTNCLN1ax0cjV+JRF5VrfkuqnFAjdGP4tvcGvS+KdXApaln26eG1c3m1UIDxV1g0V4ao
sB9uB9HJHUMCYWD2j699rfNxN1fhkSIvzCpA8v4ZfM+BH4ngUaJVovuM/y9L4wNTh/6mVMVceUNu
OWa06KxhROFZYMABZf+wOmL0XA86l1+jmNPWJs29msPO6+8jfhKNkmomwvqLweqr/NXaTTBu1Eeg
aQPZdtg+GXL8iet979Ct7/x6RI+gYk95oXTfjMLBq4eGzxJMbvEU8a8NseGkjn8rzv/bilqfrZed
k+xuZvLWN4mus7+yV2uTstso3WO1SfNAfxa99AqXVHzHLVKcsIkLtXw4HqS0jHBPvCnwHIEAEsSX
+k0GSRYseA2NVx5scr5awqHdDh3rQF8QM3htfZtOhC0lDPN19gZvZNTJtMbxZ/ntjg08INhZaMAg
o7qiDiOQuZRbJBAkP9wKx6U52St0Nay7ogovndAgJ7gExsZrqrnpkvABFd1+EROXA4LNwLfxHwlu
u5gYTYfRP9Yfq1AAufhN561F4qgTMSCVxeMl288j6vWCgDFk++WbXWoaKp6/cyf4nvzvUAjzyNvX
VoRgVc90zcm8gpmDsHW6R5TnmnP9IKXLgkWZcL2l7w5JrzV3HjsdVc6r9eOYBu4xtl6huf62J+Ob
jfHlTkDVNjnEE0/MEkxdI+5F/REheGeULwRkCmQRVcs+n/rBa4VDODHTkmkT+xOm/LJ+HFvVry/G
OU22CD64xQVX3IJdWKimcHTlEnLMJF2u99Vj8heYBM5WDLOe3Tk5bxVvQ/OhCbXc750SrIsObetZ
y5O+3/tM/pK4unW0843hhct+MIdBr9m82koLkptH6BnzfTkT0ik7PQFZa1+mfeXyMKJWoDI803l0
O5lMijGxOtZrjPrYAbQBPrhPErki3DcrM6OmkcIOiipaVyY2+ZEFUk1ujx6MkcomlfPhWsJTJz4e
IdeYEYPmhm50Gx9nXtsRWv049dIlYfqJOdj54mdXtndJOH/q5YWVNGls7Tp243DJfRUu5qjgXzDr
yeHghcU1taCUhimz+fdl+xS/GCUH8OtnGEQLPMeSeh2vLwTgm+zlKovf7G/psFTsHcg5hui767NL
eqbB48xU4aQzrQlot9xROxa/o1reIYfEfM+o+DvAMAFYcKzsUmbhJnDT5/mpgDUTQ2EYuWgRcSw2
1IDIHgiXv71HF2n67nGJ1C+zpLjEF3P8utM3wpBnKoPEBBHB1vRT+vtazLhBRu76NsgU47ctg3w0
bUmTxD17aFhqQJGJzsrjUdTQ0Bk5UBwtIRbG8ZFeXDZIMcAgKfnS6IYKAFZmnoCT3b2lFDSKepuX
I637Sj/MwkU2SXYZvejlM9ITbqn5VEiqgFuRCdr25GiwTWOzCqQuCY/sL8UjOZl+peKV8zPj+csd
AcY7eY4PwHdycQuJO/H293t1HGzPGx1f2KJ+CsgBQWLk+OBlj7rx4bg/SVbsFx0avqPHa/KRh43R
FLwb+1rtG93Ns9g0rn9WLnTMN/D5weZM6u20QevJM2T3g56j36VDgbOhMJmHut8X9POEwZdCeo8H
g5ayShxze4XXDM5cA1XX34Q+77XU7bJxzMVLf1p2OQjrOpBkEtbUsVJUjB0x+OJIy3ffNqj4I24D
d5kmsSm/ZlunEn1/dIat7yQj6+TY29EedwM0KTbumD6zpViF794NVXq2TvTFbEpD5T0CWXc/Q7gK
hToVu4x9luGbdtIeRyJ08zUOIkXPX3XCzXZV8+bB09mjggzgsqAgIXFZ1ezm21+j4wlV/CI0cydE
dTJL1kr/mrWBK0fSrzjppy19wL9fOxRO+2qDfWCEj6a3EGFyuoRxmcMUr42kEFETtM05rcMRhvl4
OhF7nn9GL3BtqAYY8FjjFm+eepZswB3/6cwdepY5mWSWDWBT7KMbcIknyCZ6OTYuyCSp1W3x+qch
nTet+7JTJyAIlcJ27lk4XxRxfeuVkcKZGSP10XHyIzkAvYsXscw4j0hHt7P74TAM8fvg7sVIm1kR
nD4wb7jYyioc0NbQppDr9K2+zOdZb2GZYxDtffDIZe8c3s91IjBOropErZfAtcbwWsFipazhyEmX
b687A18+aleoeB22oMuAEO99Dubb3Pz69pW+n0VZv7C1tJuzgbiE1e+ynHkmd1EiUIVIP25/GqYe
6xc6G/AkebAXqWFxhNxFj4aXf+7Jnm6y7ChJfO7Bi7OSVXs8mDo32X0atShka9aS+Y9Vx3YY/XNx
9Q6bK1TmFmEbox2ZXVZTdqg0Zj/Ycb/YJbCuNgSRrR/vFkz7FB7ko+TILUZE/iaDWMtTPUfywzuf
9aXP108R/h/KcYt6qoI2ZSnXETRMsZ+NwCGBx7CWF3KyAtMFFz57nxdzCiElljwqOy4BduvriOu+
6hrMbquDHJCnCBHFMdv2Qf4cOsM/IpHOBEi6oNiVkaclbjhRG9FniQrMo0KiX3cTnT2PY3FYa7Ix
V9SpVMapbVKwW/o1Yac0XISMgmAup2kFFWYqQW1Q5ayscD/AGP27miFx9VhdkmqPPWCrsSdxpRBz
CdBG8Tc3HNpGrUHPjvPLkDKk1v1vV44ivjk2La3CeENH7eSMx8sqxwsojB8VAikcDosgmLuqSem9
88tNI/4cXMQP3E+6BAF+G45A3pSLPqXn+vsXoW8RpA5utJjiRBQr85urdZEE0rNsAkNMbMdLNLxK
+LMaLmlZ+9RjKP4MbiGhwxvCWQ3+fsCmJGMittRsE4kkbJG2B7TvfMMaKEa8PiOaM8T744LRf6y7
tJLUlc7ULXYazJFjDgXdZ6bRm7AJX+9Gzn8iJfLU4snSrYdmvF038BnXCRqgd2XS2y7hIf/hCICR
um5siSxIFDFfR+i/AdshigN1/D3/YTXYL76grTjYEwYIoCOKSZHpdqjKHui47eRVB/PVvYkBeILi
aVml/QjXCyElS5/iIeyAomWA4E9o401y/z7t31I4cze+v2BSRxV3mTUL/IyjPLDJJMF1t25aMtfI
7ve8WlOLVVybyEcpA7oiORdw+WF0tIYocas4uHEjmj7/8Ud48tCkR1E3Q25rj99pfweudp/5TRif
WEcqIwCZCD7KEt0c83lDzBDtKrhIzu5SArdHhSFE3O2rkvibhM0RDniUjvQmQw9GbEtqA86P1VhA
gX1DpPcugAJzf2+Eb3usI3yfnQnm4GsoeYXVHd4EZTvfTwzJGk2dPgrTQmy7AGbiSb+BDTO2oaj8
TjI0K5qBO8CjEby1yQgE8X5b0/VJHKHwrhflOmEBsnUQUdkyt10MehxO27hQ0Iwy+wMHP2oJP5xS
+eJd3kZYi127Wsn2uBq5aVJJwnUofIDHB/cqp6ueqUe8abQ4Rvi5T8rM7Q9IupOxGORgu2V+IbIu
Pxqg6KIbQ+sJ5S3n+iM/6hVIcwuDShobKBnia2lbx1mLWR44MlNTBGa0EYR5F3IfuHiysQkul0K0
2WPMpY5erp1U6y77JLrOQSz5WjXYnJXPfGT0Dhl87WObiOFXHo6c5+3kriAeS9c/qWrXK/2+JW5c
YZIK7XyKANuzF1zWisFkUBcNmAQlEwEbTbIJD6tBg/EDt7SyHxmy6SgwqUjxfT4aNJBERdgzK7RN
R2jbmVqRjKPyGLICsanCn8dX/9XMRmQIJxj+zNrTzxfDXdoZGmw34rMnznyhIVxHUyV65b0BxaX1
uVr5r5O7/zPD6JJxrbB0yk6+DuH7AEA6nxQ9AWroChjnwjtXbgc0FUhc75aj9u1tHG8eFZtfgxhq
LDccI3qZ8XxKlNRHZCecm3Yis0h0/oLZojRze+03zalPO3JQ301ArKs5IENcLaC+7at0LD31hdrx
Vx6LJ10/aIbduOQ1wyIh8NjpAZZCKeAVbvjK9dkGIOuqg0G9ZWSEXnmaVS2QzV+OWmmvOxtBJJk0
p9Jno2WTXN/35E77b40M6iU7LxQpFiSt2XT7dY5mYxoDnDPIhy+IVqlpnWGBFLERVe7T9imrrBRu
H8mmlqqhn1WoDfHAqor3Gi1jKeBrU3aTii8c1lX+u5UJMbpvYLxLqwaWLe6YfrBY2TB0WFtYbhob
weiEb2Uy9MiBBJw20fZxQCXp7BPgROduvfXEgNFhIq8n0ksCxOiTMG/Eh9Tjj6pTBWMNEqDYKDuA
cYWiVtgVjjfVk92H5uX6l2jCWDgw5qzgj/6wnyVF645p/r44sYiiPb9bbc7UXrkH85xyEfrenDf2
LYt9B+qa4n1rDeYc3K0cmt1fZ3zxnh4R0v/KlB+HnV9GTq6QEPPBIqoD2UTGotkW2vYbLv/v+sWf
uRfOJzmK4W6HIMQOSy5w1VOg8k4KBsMB2mttpG+96cwqPfTVyDfKdkqF8exNAKnH5F8tI5ufAeST
Zm54aucjInYF4Ojpp64BG1UdHafT5yCBSwafqSZ/isQVyUYrKyC4frPyehHGIFp0lS8o5Zq0XuIr
LzROvNMfvRMJX6Tr0E7rVGsC/3S8ysfiKBAXCiYsvdTPpsniJGo6V46FandD0gMyVwScuPGOKTQO
QKGzHVbn4psj2d4UdqNzhFlj0uhBReWUkioKY1p2gY8CbsNQao4Fc9oY2U75utUOZUXgdYAji0R7
Zk8ORpWUWVcseV9BwKODAV1Sn4xzKR/xLqfFsYKEOIJ8f6O/ySuPnipjz/bRDPQTikvkV75Beowb
6WXeWlFykdpW8ba0x/io+8H9X1Qykqk9am+9uVoQT2FFzGWc/IB5Z7eFR6E/pZ4wDC2WR7Zn6Sjq
wLlXJKSaSHlxvlLZ5uNngv8Qjkjj2O4ayrJNCCOUPeA2XUqHWyjeEvoe5vXx5+tFN1omtAy6n94g
Fn4nV63ihxutCt66gkt+Nrpt0iUIRKfky3xIhbfSmPUCqLACZ4mRsSEQM9qAWwny9HnZFOhIfS8E
HLvWqRFy1ZtbM4A9xGpLNoNTNJ9ND1P8VCBEvyfZ1+EzAVEzEraLnIPq/cJP3IKiRIUahx7QxOlI
4hTk2iTNk+DmXw30zhWDdvXr2Wr+C/H/8MTh+5tEg+Y2heMMZXsmuSc7nXWvKp6twyJXUUT/I601
I/XIK2NuVRJwMJOKE+KfEU2YmUtaiHmGR8PMClP1bolgqEs/W4i6t+bkNxBQ3PHTIZyeNz5dhcO4
5LUOufrSSE/Kd9MpqxqOc4ZMTYBtVMsrVnlPNFA3uf0ruCOTMQBtbYtgI6XEaqoxmr2tJ7SMxJA9
NPHhbNWjE1oGZupAtgxPGjCzRXnf76f4PEtUOEaDMU3u7DKt2QQ79dUmELUUotublte3txGv9qtT
BVSWSXjXA4tgATKURXmjf/zyKYXJNFyfmLlDhJl62QuP8qHEDjs7OJjTbxUlHhz+Dtm+VywfC8fP
vxRLZEvq92z4U8lqHm5W38uIQvCuHn49lrhW7Mgy9x7N6TSZMdLpUvXorM5mqofIifn2fpJQUDZp
1L9J5TaXajf3iCSph7wB5vmXoIS38psu8kwcBdGE29FWfUTQ793A3+z4UiiJpnwd2K74tkcV1rNH
18GzZxJv29eYu8VcnCNQ+/7Gnfozl1xV34e/8AskAB8dHCjKfjTo9kVNdoLuUSdveEKPBXz7SZp9
mXUZaE55x8K/125CoDeXEgxi2Mld6q13oHhLf4GqjfWbBiQWOkPlUoQLCjiUF0RfjPVjp951iSDO
wPZlY4myoBBUDU3LYsD6m4Wrez9jFjIxkYMGzjPKzP0aFQgFty+Fqa81ZrnjIRDbsQLdLFR5baPp
3XWj4/aDdMPcGG8Ki5/dKu8DK5kvDgKf/gOHuPKSAVf4EqBGZV+9CowuEm36wrW5m/9lvdklBHSb
ya9JoC8r8GEUXvlW2NpC9gVx9Tw5D1SllygstX581mxOTxlLv60O44LL46mxfalaNpJw1B1aseWv
9bnPHN3oynrkid1eoXc5zCz4geuO8txYL89Rieb6DE9CAMDGeQWFApDOry04kYeW/Hx1YhE59Wvx
NJlbblzFKk728QGI00fvRtcVWPEP8JNjnSYRghC5Um/v3TyazMyPE3EUuuNpihmSBubxYHf/XuVP
M6MMTw26Uoga5U8jlrk6Lg85hYzYHKYzT+ISqTagS8kXceD1FMfYSlzviJc0mpSSts8Pkph7cJNh
LaPuz9Oln4iJil3M7PFux57ttu+qT3IHEmWD5LGye6iqbn3J0SBGAfk33CstXW+BDS9osck2Ufa7
j8iCaWwO34vhkNm3mNNl7PmopuuuusBSyxCjYjYjkM2riZ+JYiE8nNINiryX4k8BqqiGEJfblrlL
DEgUekxVFJH14CdFeB/unO18Ea8WQODhJhQthJRdreAWvW70tmAkYPITlJfz6s91q/OFYBaeg9oT
m7egbGIC1KDxBmslgQW3yfXoWikz1c6MKCS5lhqT8MpmETGk+7v+sRtQhQCX+Ha9klcXutioiZZ6
G5Tv2MHnFEVenYGGCwBjl5tvIUiuL0FegcDVSOHfqIpsJDbiQ2ZsiAjLsPmQaSQA9x9TKMkB9CyM
K1pRerNTwNF+NCsFd1AgBE4wpwZK2O+mYVb9+N8IVHa3Wpj8ZeSy9nJCVnbM9dyqh8gA/j004+uw
0pobUOS46V4leimRywicScJ0V1oaTKZWwSCRNQaSYP8ojmTzqr2QvSa5rYM1Zf+YGMDGHpxMwSx7
AOL1DlDD9JdAQ7w7vXNMQryX8APY+C/DNSgCKwrONSOaUxqVKTAZLtBCan6yhOdA9pWOVCoRtAxb
qjtDzmjFcNcNV+/PvCe1RNzk0nAHdLXEBpEDqFjPNVBzTyIdzFW5nxtNfKeNxy+8doYozlyqtcol
77Yg+qjjlVBMR63od6jab3T/tdR+r8vGGvVjZdZJhss32BYp6xuFcYV+9BU0wEXg2+2VGsRaGcGh
xWXUkQjhh1SfR3UOVYGeCS0QuhbC6JMPbs8M6eOJZ2oko7mj4QbKKBmyEbYZir5nx/PbboMB9u2a
FltDLtCo/gaB6SENOmbHxo72oAFs39zUxRM1Hla/bUkkKxUIFRG8nT1uFHZFN6iRnMvsevnTbfsk
OM2JSGqaf/4+cuTBtXCrEnUxi91Poxks0OLODDKLi2a7mY61kGTUXMSbfNOtJuTwf3F7GkjLOge0
aivq6QENrKo0mpUbLeVzNPPCi65Wok6VhYNFnJW+8+PQ+hGjvHB6RrZdPJTgyLilNoCJGXJhBYWg
l/eQ3nqiK5veYuEhDV9X2uCsciyigRQ9zF2p3JabHGtl5q2g5YdOW0V9JcL0i4jtrUbFNFUuy0Qm
MXcRCrwKqsNJjR1CwzCNQAo75aY7D18yTkV0U1xzIU414/BIbfrL1xL5ew/U18GTFlOl8pWbBpbf
UOU0vEzL8jeQYLtbLWW3pvf0UdG/iXIx35irvXznEfIZ/qOQJp1kEllS2So793Njk9QZjqSn85lt
Y4IujTZBfEf8M6JAEjnIYkidZFe71iqsDOQ2ldJhse3EVOmGXYy8JvhaaWCzqykToBrE9D95z5WT
gPUsHPELydP8GXAIoWOoRCUGgjNxwbr8i9KI7jluDcYfZjtNMMamtsqbsOYYPAPqxYQNXuF08xHu
0mHz0Z+zucPONYdM8ozHWGVGCDTB5zVT0e0tZhW7HKuAQbsTt+HZHRT/KkFQ+vp0v8kqwWmESRpr
I53rgExK2KFRKVW8xTLoqAawbRtGsYGe4guRT3G3ThYdjhEKKUaaV05+6onppnjeaQI2LtQNGcH5
IR5cEQH0BouYGQfTzqpsItEUIcNGRVIDWpIvLRJdTaQL0INTtQ08jw5UX22nZa0a+UaRSTrZGNDf
now3/2P+LGt4+CqlQPtuhyejYBZECwqZxkosqZpO/yCCr4F0+v+Z+AuLPcb7wDEgeKGzfXYH8VAP
S+u3TDtS5elYfCOQvS/ZX8hmukzp0bOFSf1jjSG31crubUIOtqFlIKiRMbV98nWRsBUS0xGHCUZC
VSLuMwjUXW4QUiBNX+wv2oJ3rs1bdQ+JGGtX1GELHFHMC+B6uJxqWyZzHJNcrInrpeeWY2SacnH3
pRVd217n4bxk8u4yOGyzgUiZmp0bqMA1Bp9c0hTpXHdLtTrlGlT3IyV+zbY23rvhC7n+/eauANxT
Tw9CQUGctGzjafPZJ3rec3pD+XmwEWAScivTojK91deFevyfgRqZHz2xRvoiHgp4wEfgcyRfL4Nr
PjICtOMoFZX0qdxZXST0bK2DOkNQcFoPvOsgyl/+2qeHzj1BCrng0cVqEYO8POK7q4hTSOcnSidC
m90t3FHuaWk7rpBzEcXtMdau9P+bAZZli5RwZ2moBwAY3+ylvyfS2hJTv+EBfJb5m5NMkCdOZH2G
2Gk3YPdASKtZZ7Gy9TwrJ6WAUvqdPqyqWUYvUeqaNeiIQim/2hs3M0WOAjFkIqp+zywP6LiuVNOp
j1RBumYOJH73kLi9e26W+I1EtruJguh1/07cMVgvrwetbak9eoLjFOw2jynV/5bc5hFTt2QxEl/P
8ImZwPcWISUrnwNaom6ekSdz93F1tFt6P2kTs+DZC9AkpxGot8B1CIXZklYkkFDQkdM6HVNAQLVX
mRdq/BuEX8sI8H7eP0iG5lZHKaXWC6Ol506d2Yn7U+AiEk5SYBwmPaJPKNbynK5htjOYkJ5dQuSD
fXVb/lespEeB4gKaQyhDjAtyJD9ur2Ulj/zVneMSuV06tvg5nMvjucjE6O8VT9c9g9NhEqw+wOZE
bq4bBmVCvnqeiTZjuMtrXPfbm3usynFMLAjZoLHsOxyIKN5ClTrxs2Trm9Y6vpBTteWKZmHgY6fz
ehRGBH3I78I9ZgaCqJUhZvzkkZjL60f0Ah45ATFJIE7XJ3I/+lvzjDPijIzWnaG5jN9ilnkOS+JP
ngJ/r9gj1810qSdAjVjbQ6bBIXVNtnfR47kVTeXDMqmx9R0h5/sC/AbGoSqnk/7xRTwtIn8S0Y3R
NtBZv0+MgGVhg1v82I/yXuUea45QjhM6mOpIhIsRVLlpYq4S7MAsKqcoT2X5oNXGpp66NoKwDdMI
B1C1lfVlb2MQJ9q+J80vWcXo7o/+S3ZcPhI4/hXgY5FRJturubS7J5iq1lBeSbqSCsZrmfUkgjPU
Dd4RtQDZ9bnKGsqJDODjZJw+Rb/TW406siTJXTDuNL+9q5W/KgncQOQMejd6ctx7JaaOJTMN0hNM
n3e+mfCEA482NEwWmALjmH/I4ort7/Qm2A/D59NrUK5UszTCB1ngXs469SJtpmsht5foAo/Chb44
Hlv42RIAyWUIH1NQMbK8qD8dtxHAb4VRaoXpaJj4AAc3Gvb/SCY9yVubj24KcAO5Wvod7rzduQKw
Gn6jp7f4hVVRcDCouKeUBcSLQQAlIC7jEise7osmu46Idx3p+UXSNB1rGuZqdGAojQmnATQZgyPx
DJsCoT90YzH6xdwXqGcjKbsEmjXRATz5IxUwvBX9hfrJXr7dfru1PMljxIER7JDORBmrVqgt+jBH
EZHWR9fxDd+3Hz4wqtVIFEe6RcZFpARtA2VGswWiQhj8faRvO6pxc3G//OX6U243T93oevDH6Gen
VW5ipJLCtHTuW3F5t6PPwec/ZeN4qjw8rhrETbJne8esQMIcj2ZeBExAu8ozpyjZH1bB5QnyMSjS
zFqum4LQXCpIDIcTMrqSLVylFN80n3bACPOQFT3SLHjbXBSd56c424S1VWYDFPmqk/lRC5H+OfL/
klfR9nPAJu19Q36wb6e6zo5B1dSWN45O5fLWPrmBGtOcr7r+7IHYX6qhE1fZDlTKns/Ad/nVIlsU
0oo8C++PTyupXDNhXwKZ+UUmfn1M/PW+1n3iyaMAeHx+hrHYcRwYJDgW+DrDRcV03A8Vc0DQlw7I
yxQTGV3jsDeERv+l3od3p+qNnOPratnWNBepy54hSbjoHTLABaPrl9UMuVTXrdkaHhfl/m9SRygO
CeGFO76mXkENDxw7yWgsoWo4PFx6Z4VICnlDGLE985vi3hFpzwAybo+TbZJ4+uPEn7ZgK1tTwaYo
RwVxeHh3csMCnHHvvaVaj5hGUapeZ7T/DCO/BUBd7pXCZPk1kEoliWN5OOmvcFpgw4KKTMUAbwFf
Aqs4dtHswnlCFbiLfWRrDs50jHMHY9sStjHryxiC1V2D6fMU6orANHJsC2ekKwQpfV4HM1CMvnNI
Is/79pSKJlTWz1q9fnTcNnz8EA1arxFTS+OEwZo+Wiytvm1ZwnjVQgjTGzrdx8qYZHm4iov9c1SM
aBpOG1JhTa4o3Ev49ttnYDqbww/znLAxld+cPniBVo/+MGIpVSxUBQYSIpV9yEo5CvcbgDHdk316
fYSrlJVjQbkb+P7g3y5wDwN/cPzSih1nPPiudEBFQQ5zl0+p5gs4NuntPL6j5xVzxLa9ALB0YUx5
pcrvv9aeiOwi9cFTtQx75SnJHW+gZEivvpM75iTMA6SB3u/+RlH//WQ2e6nExM5yJ9+vPORJO+U3
tl5ylRE81nAty8gkNPzGxlBv0S8kZFIeYqzuHoTRIHXQUWx4s54p+BCurk43+uiNnCiZ1uw4cjW4
VD5LiEQKfjU99V0MEyzvo55KFfsLKRg49MkxCy5Vr7C5mN/qTPe+XH7eKZd+/rdRg7qE4V3Sz5DN
i9kNQFT2K5p+ErDUjCOIryZci93OLsmG3XC6PAVIB1Qt+pzWIHfEyNI+xq4vIl2jdVbiRwEEO6V1
rzkgHqQ8LGy/Ydgy4nYPBMWmi8wEgl/9rcE7gKMxxm/eJO66vx0vk6A+qP4CWoZdsXXCk1EeAq1y
SUHMK3czVO27k/pc5CAqaG4IBG/JrxGf/yr8Guv/WODp7YAwc6PyXLVt6Tu+FLdSixNwC7tq0cvm
ACi3VkLN/KpBdLwqTREjONyxAN9efUEY0XddceI+uMfV0Qp3uwxf51XnY790Ei9KyMGB53Zgwywq
1s/9Abn1EAWW0tgBZvuqJz9GzwniuS7e3NFEUosxY8q/btKxEUJAp1L3A00mrTYRVFJ5CRmxrTB4
Ol0acEWuDzSojlIythRtZ3urrgy9msBZEtHTllbSWQFPvXe+FbovJNSXanMJE9EdkhYdqbYb9LxM
BLeTX8/syZO+ZjuBu4ibcJolhrGSdwKksSubbReO+kq/mmCTuaui3yeClKllz5a8kn1DQlejBztb
/hSZtBKkEgGfwnuoDCiKsE1qB6FDWlyt7kD5yvXQgqz3bYbbYl1thW/2415KuoN63uowJVNcDL1T
XqTgTTRGnxrRJ0rQiIB3y09ZLFfooR1u1NB0MajZ+0ZLaaEg//8cmkFeQZo5xLJ7RN8BvrJ/ntG4
bWo9vb9C4v+TYbOqY33kDHm2dMWE2iYiCPhlqyhucpPQ2dpJyIxpRoX5OUd6fwQHzWE62LtuWnbc
ByBSksz/P8t6vqi42LpFZ6gJrFj8Ig34AzKAkYgXJjSndxPJYvl1xxPX5myQQW9TTaVkdSzm300E
sn4Mq7ev6DzoqqRg4wFwYvIjHw3thZpxJCIvBoFWpA5la0wF6x2QUy6WS4jaj/iOb13ioSmR+/KG
a6hBdH9YMRbWIGlpMwfuNHbhC2oqikwWn+Xnp6r3V26Fi66eO0W6ch2vI1CYtKZelejEiOt5vdhX
2N0WnZirkxVOV979Hq5SvYM79kAxR7Rc3n84zd2LHIp+BHNWArtFUq6J/nth+AqAxrJ4JlL6Fy0a
dQAaAiA00tiKG/BQzy3/2cjhQLxtLzScwtu56/GLvq1v3qVJWRx/EnaPV/Jliqepe+jI/PRMTpgY
+D2Wj39QhkChdPgMHblLJfoKYWYSEIvZBQuByw8eFvPCG4ysDiUK7J3JzIlRD86d/zJLUdiy+wL8
4x0AsTTcTdB7Btr6bOpuC54Frb/0zwld7YHz/ciU5JK4Hokbb/bXLJAY16OfQ70OCCcfhyKFgIms
kWJOJuCdwGBLX4TP5sob7Y+rAfO58/oyB3ab2rP7FvAENG/bLeYyxgTt8MU1/ooPWWTg2ut/fjIz
s3yUPbQoyX9OFocm7db27AM6FX+XNTpvbP5HTwak2iFu+KGEEKE3uV0Yi8Oqo67vTy0InnWRt/Ir
s1C6P0C0Z5uI/1GYqkjtEgJuwkp+B+geZN9mb5y4j8HmOub9IT9kudCN8CU+DhDj57T+UTGofRPK
NfBCAftaOUC9f5LBQa6bmllMw4fmiQxbVRA0kXvlvur/SeT4i/EKUSnHAGxwRf1renTG07Qh/7tU
6MYxY70wSP02/ZevoCEgxSxs0BLyRx2lmkM8aQGwe6EIxd+64nuMWbk19HI5PKa0vpHaYvA/IhWF
gS8Jx3dBTubWxcB2bNvLk01ikuMEk0au7eAcQWFPj+ESYnsu6aWv0TDwsQLYF4mMAluPP1no26rP
psbWXJECmapqEPVmszSoMuTjXmYuG02gIyY4NsVpzQbjVQ+EIUYjueX4BxaMlP8S1ktl9Z6BSAdH
EuPT1bAKXHkdDTDKO9OoItI49EHKJ3lEbG+mXTC4Kf2rWbJum+oiNQ0BS7DCrbHDho4qj6iz6IAk
Vacs1ujXwMq1nsFshoXqiZAGDGp3pLU+N5kIQeaMhZrIGTrZ5IZ/PJ1y2gyibo5Uxq367HZjSe23
p9wtf0smerCXbjkahzRLz7kgXFmtgH9yP154k92zzapKkj3T1im2FY0RCT0Df0IOlPCIxBj1xm/8
LTS/INmXrJCxf2MNpMAfpw3+CKSKTlujiVJFy4xdYgQVk7U9CqvPYRmA76+5kwc2KAQ/paUk4GcB
aIRO/lclNgIi2a0uXiAW3kadgJGuqGIw1CT6tryUuxz1wdc+hggNZu54fTsFrN7FsiGJ+0Pirpmg
2w6+vW7EkreOZ+fbV+Ug/TntEN28nJP6xaHCKrN7Xki1VoZRo5/0ekaQfZya2bR8ChY0ilkpk7Hm
0Ihg3CS0SXRp7bL9PyMvRCCh6MdiEzIqxozllx+G34cwdo7cawRzVo9GzKzuL3tzVQWghvrRD7X3
9HjQPymXXEiZnRk9gass5RWdcSDXIaeqx9Sf8h/B0qJTui0NKGVTF5BSQGuvSt4z3e9TmCx2sAnm
Xbmm441XWcqFYX3EmBy/7HmvpO0ipQYoP8pwRSrC96FYQKKUeQrF54ifqvOkRpsnVAZAZ39gyVaR
6pjxMGgx4afXvsnz+EJAOP8KHx6LKinQehxC8jB/WXrAky4fgKgnAbYm0Ujwe/ayEGjeAdXJHJng
V/9dqx+YLBesKeEN0W0hdZRg0nxtM68tqPFQrJdWAY8dagbEdA20cHXh11pGyJ7Bb3GfsqPXhvDG
P3ZC7lc12noPmVmymv2dbMwrxa9cYZDz2Ed3nH8xsuy9lS3fd7SvS8UKKJSnXPCGXy+xCuVroVr0
ZmKogbW0NfDwVW/AkcIXs5qH8bh9m8vC9O0yjdEGE8zzZzp8gjPjdPgSeIXRRYRYwgfeKqYmPhJ4
UhwEjUBE3f+yTfDf1lqD2HfoSB2joNEOrVBEonm8ulGQqEA1lIAvdCOLMUPS5rHZWH3dpSplgS+6
RMWj9+C/ft7XytN6NKRwjYG08uVNLdpF3WCoDttR/tpJ/diV4fVA8p/hC1jhPFnkC5SbidG/ruhG
JkOdM3dyyhcpBD4oMonU9lBub5iihB4ERMFmsoLgAf0WQkLIvAoN+uHSOZyVge1l776G3dY+vINa
hUhC8DJTGRHpnptEl1DmeCz1CPL8ELegsSc4l2DmiFWmPW6SlIlFo0XsNhNIh58fA5wNpU3I13/k
E8e4RGP0KoUWqd5eUkgaF/fVHrrp4p8/Otzted7YqJHMq5QLE7rkw5q/xMENNv4RAGRHXyseDEfA
1tVRAzHaQ1iGvbf1cG4irOBlTiRg8A+p2zx0Ov55wXhQZjyWwTEZbjsFV0k8yOOY/YxB6e6qqOmv
QUHss1zI9F9OA8hJbLjcvyyRzYwEq3q2vHFE3VBr4G1kTyi1O8yCi6WjzGhw9rNc9BsvS8AZ0DRu
1/PTSv58knNUpq0GQ4MskXqmI6oRm4fpv+wkxacZXCG3DXVj3LiXjaNLf+gDvc3lf0ogwo9H0aT/
84EZJOTa9GnItzU96ULxLrfk9u5QVGyHMC/0VdiRfGChAsY3EFLjrjtSTpbF5iY+iAEr3eeTKKkL
mSd13/c3JpcnsHeolLTMeYEfz/VCBY1GsdS+47pYrYg1tmYZBJYdgPY5Y7KLvE3rOI1dVtFxPI70
N1dxqkxS0LSieirhHSlkjNTY+YrEa5jbq375/yOzEZAFVfMW1LT796/6pQIP7rw3tHpOPZYlB2vu
Wr/7KEn0XR0Qbdojol3Ww9Oc1+LwkSupMHQLcz9/y3BkEw==
`pragma protect end_protected
