`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dokINK0kjr0Qvcm+U35FMmll7Wc6hRR1mS/xwi/pKdPjJWp7I57Iq8sxR6wQj5M0
AcGZ0W8Dn4FLdrjTiFAfIclyUW/Ex9S1tun6pkovJqEIa6qxyYCHU5S2Q4q1+Z7A
5H1IqIRK390QrpO4UYOX4RqLQ7LYwSaEnb4/6YYzH88=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33216)
8QlXcZ0IUZRQVA3+0oetbWgyaC9ywgH+iW5ZP2rDJHa8IauCnl2VnVAp7RzngM1o
B6DpOU9ZVCp36LmkIdG9JUkO1sWYFlIiRJd3Bqnl2l6JdTUT4K5QkRHrZeXrK5T2
2eEkrhaUo0VZ5510pDNT6dCe2lUtmsRr4qfqL78bgpBZO1tTbjlXVszlveVCo7Ws
5jscmz5dRCVL69MOUHsuj7i2rSZoOnI4UEEMNKeXgwAOUryJAkPXyAk6FL7Sl881
XfybiQggK8v0mEy4QGvfSqWGEbz2nPgKBqpuHAuJjy1UPTDyR+/ZGckI0hhxwFPl
DR7nbo/cdWS4cuIO3T546SrrxhnxgM6P5CHB0B7OhnSc2RwjLjQHVTjaKNR2H1ts
8b20ExPYo7TLpuevSBR6BoM/nXkBhms4FxstC2xuTURN8tpMTOTH/8NmL9H1DFQa
xxEWvqexT4NrAqWESYiNPMYpEtIksnH48NhhB5Q1Bx39ffecWWY9B4ESqHLOvk3B
O9hcyoyR3zphZ2NJo5xhzlJoYmM0GvDPAQcs/BHfRsS/BHDZOiUD6HEuwDzdc97K
bIKlV1nSpxuITXP2qc6JmgzFJFc7sRSl+vzluODeydw/6GVic81P8pvQfVLod7WA
ZLnrD9ThnJljA/R/vHSZsUZNENRiZQ/rCvbetDtUApL48eMlmO0EwPk4w4ybmYvF
2ElPmG2md5uQUmEIwqHNLP0/jhyP12U9fS2X0t3tEWGZQEPfjomz6hWSNEhG2xK4
DHAsCC+eCrD9HNZsXllzAULcAVGNqqKMusw1cNaOn1Uun997qPUzAzSfWqLFcSfZ
dI4RG9qVl10ObErNK4SJ19C1npvkIs/8W5wCq48zXk/cwe1tAP8+NU1q8A+37YOa
jTimAmFPC4B4O/dZUl4NdvHJPYxAscCgl7Wk1npmMgfquTMGAbli/WY61vrIXTyO
x5iwL2Zf+XidoXE+tLdfvbVlRuRFW5k1kf7yo29/h2jD0vmauA6NpRnxhVGcm/1X
J34rKgFe3sbX5Jn1YHlvh2dDMb12qzNkuLFSyPiXIbCT1eZ3jnSZ25nnQynMbcii
Lhef1TFqytSVnbCkWP50FuAZkv5bG5o/2LsRr6mVuNbR01G5GqHAAqGKgFP9glr6
o4IMCLlDHtnk27vFinQ7GKwg8DZNPuIQYm/nIVHFUj44icdAJ30IgZaZgtMXeFpO
H7SRtoHdvHhSg7koO1y8vn3uDzSo1XtIXekGcvFkisFkP83JFk+DFm3cvPbjOyf1
ERTwqGEkVWylQZZol2O9MIGNwIF6jamQNwtopHOLR75GjAyS3Zv50lMjv5AWDDGR
QGywcFtFuHU88rnUfPVdwS2YsxUmf4O9XvKTFUC8QxJ0owwOOeEl7QV7/VBiJu+0
gMY0gDzuBU1kUiHV8N9lLDJj2i5riYuOsgDMI2n0EnPfh8ZvlHWH7eF9dX9g0fz+
1JqK1pfAufOcg7jyGGeNo0oP8iBXxhWRUGj7+ZUlZ3KXnTIalAGEjPE1CRidk6sJ
yfjgupI4QpfiwJ9SPQg+uns1L7w5Vh1jY2rpgNabMBcRAoc/UnSW/0YJjUE902l9
2rss4ZkXBPdSwFmpArU32N0cty0WqmWgZNlJesgQmaAVE3e2Ey+jSUmKxKv3vj6S
TZ5GR7CvRFW+KWPAGebj6UBLKe8iqVlBlcjol0hDmrVFw1HSsmAbiPLe3VAU/+gA
akJkbCOGncy0GcZYc4RqINHzeLhmJBxCq38vD5bhd8OoRc51V0UFfrCalxAIY03Z
BOeDufXW0+RtHv3DcyP5cI0Zai4DyFTlTeTFLtU+epiNUrqisz+L65+hn+6Gk6Nk
hvXlrnkpeJ+suzN6PI0QdtOAMc+AWwDjofDwUmPp6cn8jNT5eqK49VJ33ZB9cmrY
VoWfEdJ/CKEYQay7QlkdmqX96rET3uOW41nwNnaEarcTAVPKMIQ0rXt5PIFqw5xR
1kRodTvogQZJBfReIi7WZu77O0RPzme593qydFWvXB6Zq0f0x6wamW9JSYzxFN4J
KyM2XRpkgRAjhAfY7gTwu3wwVbXJpgqfS+lJlHZzjBZaLSxZEs73lP81Ylq+JYaz
bzl2bl8ajd3ZTb+vVFwASGSf/VywTISu2p93N1cR1++62vCvuFXRXtVCa/IfY9Lp
LwdNdyOAF/Iedxayu0jkI8z1DJfD06iQ6X44EWWs1idF/cGLB26pLNOEHwFyOFUp
bo3rHq2MYw89Frq/OXNI47MUZVpo581Egmz/TH199EI9tYtEEfx0qbGHj6xyMiv6
0J0tkjlIX7vLnPgMrYxUymc3wmCYsf+GaucbxX/QBOiJn8nj5odu/bZqaab2oJwZ
pjqQzUP4UvEJXPtKkFTTdOttSantbuBAbU/jB9of0cuZvrWwQoDE+uQE+S/G806P
PDnPuA9M+n1S/N7fefPo5yv5iLEde5q4VBxhdpK4z56Dqgg7+cz/uVOqZ2uWJUdW
Q2/8yVm7XH7M7EJH5BPt94rMTjB/2V46kthAZkNfb8TpB4XYH4kLBIErcC6CAuq0
5V7CCDcLo/B3e5u1PxbmNvTIOkKI5dt6xNE9bZCyO7BxC3rJCdTPQVv7ysPZd8pt
b8OkyBXjBcpVBU1Mz6geC3BMCegaP6JZDYTfGsndeICsCBeKduTtJCQXLOfo8b1q
EgdD8BgJEymY625+wouEyLGrk+8kfYpP0vC7YlsRzMSs/vLDyLC39noD0Ux3ifdh
zeXLprPZQZ0DjpY48jT6zr0LvSrsRot9E8rsUkAMMPGXa2xzLC0RXaOWeBGt7AFe
CSYQYRyEQM/K7loM6WCEAnGf+kgXtLo6TcKVeUWJE9bZVF8BjcK3cWf9x4bwCwb3
DgflKBzaQrM72+P1eeLfbkWNyOlMjlEnmABN9hOCTe+b3WixspsZsA7v0jKLi190
WhersoDowdmcMK4c/1spg59kJ4UXa7D5e0IXZqpDezwe78D2z4+LpiVqfYeu8+Fi
qZFycKtO3aheep63gVc/CmrlTYVFzPRJDJ1dbtbUCfvbtz1FbVkr0eENmk/f/5a2
meZhd9cP1HFXBrMP0dpjogku7JTVs8pgnbhfeNHHjAXW1VqwtkOPWZUhTgmU7GF4
R6tOGhF3AEz0aXy8CFx+vPot+KbxC6NBBZfpsy7bna6gb8p7I9xgsntBy6xY0I+U
kKslIC8u1F/9B7jqPzvaGnU7H9yigeKvlahKAN3QZtWbtODFfKzsqRJbvW1cyeYY
QE+lpBEkxiJxP22zEvxn6LDrXqpCxPlc2kl1bgRnNp3rTRjfXGMoOg6X1JTm2dVW
UZGeMOBez/wGpJ6cv/2Xp8f6R1J7Cg8V6M5Tpgf+diGOSKV55XLzo32OQw67GFAH
NwXoou8No0SskyJM91m51glx4IL5GEYeX2Pwwo32oXCHNt4pz6aEb+2qIYgHtvNR
33W2ATF1swgDG6qcP+IJ/MEloQfVYwV/Yso1DOo/bSZ/jfXNGa+ZB/2fTN5CG5kN
XQsZBNvR4+4y7C2I1Nvw3v5iY6OgBEmtjwj8zfuQdljamkuNeUOwzizFHmOS88Jq
8U580fBrshNuOqDRJvtqFtW0qdeYSK1I88oWmwrJVVAG+MOqbTw8YSgm8uT7AYWR
tsZ/KQ3dR09jMK8S87/0GjF1YKeL6hyoAWgGYEyz2Bh3VrXPpfwF2C9kk21sceJS
g3z+HF6D6FjyUhE7i9znqN2FgAPkR9y5wLoGXBQ3r8TKTBgmWlWhWU0HrUQsZ1RS
YygaCF2l7IPRf5UM8hY6o3mFvs6xnU03Ztc+6jwS7nS1sJV68QHnhP+YudSUjZup
99x5XRGvNLGqJJZhQw/TvM8A2Us6/ddjew5JjuFsRVMgiJ7/bXKIXN4ipQO8UDQX
NbPAF+P/wxfNK9U21PdgYnO/2UiL2HTQWWgHjWP4q/hZRoWVBExcfbykMA00fOBm
FCWBVbg3Y6kad0ZNR5K1lmLlORa+E6Z0Y8T78IIFY3HoxpGn9B1fOEUChnS4ut8p
oJSvNbbyWEJqldoMWcpBbD2FSva6JTMI7LBF34I8/1qSJfXKDquYLtKpRtAFhwWp
TmNjJn5s7SsIu5LGEHI1rVsCABL9CQFBa83scRyZ1KvNpLcv5ZB79F21C0t1VwTY
iGmbeSB0c7H7rs567XqGpyUjizXcqN3JUy88K0kh+aZpI3jHM1QLzHlxan0n2ypc
J0YzyJPGSfnTwlFJFGerhQgLjTHnSCqs3cf3tN8Vsej9O741z2FbAuN4Hq/m1Piu
xJ9f7r+0wfmO8B0wKsS7CxFORimhPNPmUD0OPIavdsS8o/ifdvVrQKuXWNSYHNeT
MRb5mbcOtsAxcQm4gTr8QbvgixjhzFNWn8HxFfLiWrzTQtMxWM7LYNv/WAQCYvEH
BaM0HUrE9lG+oYMODFJdz25+YYPKy9qDAVMLmrDBk/93p/Lnoxl+VzUcRYtaA7c7
Ok7SjOQDJhOmQzh5ubMphFP6w7fsYJdEb+PkgW+IrHRoCM+8ujrrbx3jg5WYQBjt
NAopok3er7AKU3tZWHBPwFzmiQFtTAfa5Mt427yE1xpg51asTjk3jj+UTpXRPHTc
syzCWQEBY385kfVfCfloiMkyQhEzjEq2eE7kj1qz1ZFPIDTG9t9mxfEtI8HQqZY8
LYD6mineYeB0pWfINDrM3IjWRJ4ng/Ikhw3VzZbH5Llu7mRUeIK0T1pRIn4MR5pI
Mc9Pe6/i24GoQMydAGXrmsaXy/2bZjbmiGVc3Yax1hmwLJ3jIvRSOBGUcJB/lCKj
9K/yu8oyCLXLjeOAwcE6ODztKMMDeQKdT/b+Q0AHKJYwvLGfZpUfEvBZj+16xsCH
u/EEfNaw5QjCqjCOF4DX80MC0An/sIoBxo97Cv7rrSmaPl5v0ZiaqJS5T6ahDReT
Uj6SbbKlhWkP/RZyYCIAAkyMpZdI59T9ZmZcoLhqPPxpV2wzy0wB/6HxF2bi1CGr
Xojkw3cf7N5rR/7Dq+Tb1owcFP0Wol/1zg3+wJEG+MU7u6/HsOlLqmZX9oC3OT9/
uEcGOeiaqLyJjoUBt/eMaNmaN7rxJEBhiYq1pzXBFEoMtc7f2fF5DNNGLJ3wqQ/0
E+3W6nIJUcRw3JGvnuCyGHPY8+rWf/IvV9xzlek735FHq7oiAER5sRB6DZfRdsNW
bQjGKzhV4K2k3psOZzGZJiudnsw4S7CbeBhgmkFK539f/gqGE44JhdXTy9YW96BU
8bnLLMdP1mZsuSgr0ZYsQEoeNCzc4YC35+JmMkxdZHKPoH0JakCGYfg4hGgUApiE
tcm7BzltJZByMfjbQJOQnKhQLDJSY+ItzdLDMKYsqmiOD2aCoq1SCNJysDmkaNIT
M2XQl1cmILhSxiuQIdhdGigp+KmAAJtnkpLT5lCaGug6IN1LCtOuDIg/v9ahBCVK
9OXyXQpVLNaJQWGjzMrjLNpASoXxqFrnc2vl5YfDFZ9D/qcFzKSJvl5+h73xwdIP
YtQV9QMccYBNhAzkYkecQ79NIRdJaRTeIcSpju/6mcN9cJ4pZCMGSqnqeHnbndO0
HFCYNRmDAnyV9wPbsloqlUOj+RDvfyLXOZUTJmz2ruY2fzkCk8VSCywki8YYCv2f
MWkhGEL8hK8DXIg9pusEHRpf3DqUzyqoRJUDCUcZcNf6PBmt3eNq/6hfSLkzRAVS
/SdngxPVsv01+YF+DcwhDgY17zPSPfs56748V+sdHjYuiq5jC9XgY8KBiCTIKB0u
eUlrJ6zVitRDntNq45Uwk3G1IuH6WpzVm+HZ5+8I8esFZKKUQ262guSiWAUuzc9K
uxLc2uNxFsZ2o+4v0Pg4GXynjuSzXlCjP+F2YfYABhGnSxaQhHrerGD4JdqDtM8t
oA9v6ZEHK3FEUKuxpS48UYxJxcoa/UgJSK0XWrx7EYcEXtXh5oDqhDvSSQljrAoj
wK86t6FbrfuNrAwnXMZE7Ia+7qDXCG4nresZvfgNN6q1T1rdngMrSpwRbg2VLQcd
uuNA5TiKa3cICwW+ZTmn4Y0XjoH6tfAmGx0FInVVqGvFd+aT0kIhVZwo9BkQvQTT
y383Nj/JaoXaHMPgjGR3Dt/ojO8xE3RqHJsA5iYh1HS5ZRmSQSiI0XBIROwWTz5v
BFrdgXIHWecl13FYAVjFn1KWHhZjZxr0xbIvtcQwVCVmBU26MMdb68NGYJK7Ec5Q
oooEBrbhEbNX44wQVwQvSN76slc0NW0c54pUC0y06bhyesaczYqwxeT3YSeeUqLK
mImQw2anNnctSa2+fJiOw864NwmRkLo7t/aIxmN5RNmv8eSiQUwfuGW90Cgk7hiK
2zafYfTE0EVvpIcmJa7/feGfWwoGNy11iZEn+th7w7GvYEogge2srQXnMc5khJuT
yZ856KXBtYz9id6Fz/PIBPZl6+vuq/yBdtT1s+jO/uhDl85fYx8nokHW7EfAMleW
CIiTNYypodxdlCokZAajaLMGCHiNg9D+FZtbbkb3kod9/aYy0W0CbKMZwY1ASKWp
Z3IT3DiEflg98k9rSiSCnvM37cNgzRnGEOdSIqGTsuNPSX90thDfPma9HI7E418w
ypxaZZTTlp57ECd/ueUHmooheMTSx5QYaTavfatCj+NRNisG8vxInAXDpbl5FIQn
2b0KSTnkj02MVdamFqXFOUQRIjjivjlWZv1wQQ7fbo+ocDON0XDhp/4JvyQiXo4e
+GdoajGLj/STIDMvzKxPFLn+kP+J3oEUWnqtYjjI6qu2iMnUb8MJQRrZNZHJRkNV
IHCrqwkqguqJOu6d5pX/RL9LEerBohHtkM6GwfILK/0Ka+xjbm7zWcCqcOiKabqF
YOztZm+ShXpwcP695xLqL2ONY/8ckVYXAsiyo87mB351jiFnxf8l4PHEPPyXyAZq
X6gFChcrskTNP5FRkACJ3c3NA8OBIeK1yZRa43Qe+zCy/w0Q4HgMbZpTzZto9JyT
xn7u3kXskkFCE20VyLwOhTHMuu6LsWG+qvePSW3eh3gZ1ZMmgmNoJQibmWx5kMWd
qZKSJWFL531ygo1gZyF7UEECIvzG1l5SkZOf23WIn2Fj8QOMy/w3gpgmOVWGlJFt
k6bBWmyrw0X4FhODQyXX/nf4OUQg3xYfuBSiTWR/FTUtxzr9CPdeqC24mCYNGxKE
AadXet4qlUuDEG9Ki1PCpm1Sq1x0LqKsATTPoyBnUB0Tkjnd+RhLBuTT5Ta1Z3Ax
H2bPrJtSy/QtdmNefnIEFAQMKTiZAEaPvtoAoJe6Kdthe/cFlTQ4eycXJGmqVHTb
qlumydSIQQYLBUjA7ewlWg9fJwRVNk8/8jbgOk6X1x2kdz3A36njfo3+241AxIwK
cQx5Z6XwUipTeBaVsNYNbMRwynt0antROoM6FxTuU9Sy2yvqXBBUgmaGXgZWvzMM
QOAtXqtjJmmsxD6psV+4fqJCjEpO1UdaCFk6Kh+07zjPaKtpedgpACv42GJF9txN
etZAq9AGwzaxm47NcCXeGPKqd3NbkyI/yWTQIvhQmiO81S+h7uejOSTw9C6p2PTk
kj7MrvRszTfuk5ie/M6GcFt2BwQ9Yh/JRypDRX+TcSMJOb88QjSYew5RVUM2FVDu
VnKfQdswfP9dn4UdLOePT1sZrBfMXPU0j0XzDro67DwA6220b7WbWdxILYKDbHi5
bXOPneVu5US4dGS6KscpsmVNfODXSUMie5HMfgmcUzwJvJPLpHB5ttNY4NRXddD5
SOry/jAqaw/X4aTsNjnq6B4H5EqOQXNbFbAHXe2KQ0+0jkkgYFnyo6XnvjdQSTHE
15ts2xV3VQ6FVcnwjhDi6le3hnh6VK5nmPqLhj8mDz44XX3N7z5P1GOXTXCX4N1t
oLErchOp1HXgqfLuXi7LhlfFDPD/FuTWmNiKw3J5L17iBoYpYuek6umTqk6381Nt
LPWKRWMYSpUSuJsBl2F5kiTgqe97U3h2xJp8lUDyzFD6hIPdvbMtyfS1nn6Eet1A
NIANBWj3t4bZAvXswBctwQrt4KetT+b+bLViI+vznfjBT5skiLvuSc+rd1W3udu7
XDNmgbG16SJAB97EghjuL+Y5vofB1tY3R7knLYdNdOKYkEajxMD/+pB/nJF069zm
taGag3xz0vUPOpTIAu6Yt4gfOm+PJZTpyOQsQboqzStQIr0CZiPRg5XPK+O4v25G
hwwF6T+GRvMbkfboY5Fgzmhznd/OErorjcnzzFsvV59Nmjfm3/xbkZCx22306Nkt
DXOQ8AxwdFgM46uxJE/Se+N7+K7FX6XzsZhuHAdFRPXOs3z/NbrIwCiEP8WMvWlM
6LIxIlo1tgL55Fk5KT8TSqsQvXXIVLsm88JdV5/oinIAMifCND3sNW6D74zn07lL
SfBldD6UFGXzU1tAIMiBmLOFfUy4DiXVnMMIVs3COmA235VT250oesln8dhXKVam
CmhyjWn1MOXgv0bw8iqqG9v2WIimFKrNU7owC8Ty6tgEznbxTdtwyShVMr53EG6h
rDHHZK0vZALfD61eL+90+Pjks9Jnv+8X+c6yZHBIpsePXiX1NfcmuevVnE4QhWsl
J2h+BQqysc9ptO2Fnnj57ffwKFzS9M4aEq/TfLJvevIrgq25zLZVtPJH91jJgLE5
3HPWVX/WZVm04MF/fKiFH6M/HPdepSd4iY0VA9K2pvrvVpUDIEPxwtZKJSjzmHKG
XpyJzevQCA4gjJF4q26ghZj/5myX2QaEMk8VBDvZzY9YUQ4NpasWdiCEJfGEstvJ
oV52bayW8EwK1RUgTv/iUyOzRt7IWuNcIoVRtyx6PPqQXwtwJvmXGuR8dMREsX6y
QXWrQItYV7N77M5z7Gla/4qEA19vGR1OOT5MiA+S6LrrbT9uj+s9GQe3274oBhnp
BAlwsTkizvB2b2CHC5j8Kax1ZDQJ5Go63LaQRO8oGuut8Hpa3baf4RBCX5akbPpY
hTwldejAdp9OYLIPgU4rO6HTmknGDPlqUlghE+jFmLZUkWrcnJsSa7OvFXLNqFIT
xYnxGmdhrjLJZfJU2pKg1vjA9CDEzVrdtKT964lIm4CwhyO03BNUJ3ZQSlPABQ7I
9afwnCVAZIUj6awJnYxP87qY+CQlk5KGmq6Nxtf3q1nxLNViHJ5pKv3ha23GN07g
M8Wsk9HvRc5HBvhqE/tibzXYCWi4gM595YHOFbe2TkOdz/5oRZJhSLaJZlEzpbXI
44PpGiNYEs+EGv6tAON/dY5i7z8pWw/9FniX9taMp0M7Cw60yZXiPn27oCYPJj4D
jMahyQhdN9tFJ0bo2vXL2+JlorudUKeadSK5hM/+kR+MmKtv2JnGz/G7RU+db3BE
vjFcgIzjxgyHxqm1kTTalPKZPaFpiTjo+dT+9J3IICYI8jcgTq5J8kCKvdE9MG+s
FZHr86MNZ0BCv3ANJWyUlMZJ/CgaL2/eIbktF3n1E4mIXiQITxZfdCFKpSXkJlot
6ydUk5mOooaXh/PO0mVpghP6VLnkbnUj/z4dzfvdfvAoYJ6wlkDDqEY/DcX0YjfG
0oQ1CorfANKK4i8YkSlfJWZYY0546r9wdkkofYvQ53MBt+loOCSQs3cSVQ++Kujw
r+EvPhF+3aZfWmN3h0TjM0Pr/H9uDewsgxNtUGqaCg8wQyVjtRaya8OPfgd3pzGN
ZvqLgJCOYdpo6x+m6upGiW1UnX6ixVFw5FqN9TxjBt98xXxkjF6iZqunG+Sqx7FV
tGD2GvZQdkyd+7fQZ4OAuKdcgoJunok+kOBgA8E4hX+2kOMtN6UicD6Ke9cQp7Qk
GwgLlJUnqROl7PAiaIzJnto8q9PhhlNMqsw2RDF6KvIYM3Jm5I/3GSq6CfsEI/LS
XTA0E2viB5E8uDS8Xdhe5cJ+SKjzUNqiqIa+X3basgvCESfNbRuLDZaNSo8Fl/MP
1M9huMiceDAyChf/Ic3KqfladvV3IJTC8pjbrJAekSseGGCcNIWl/2LkH2LbCYEj
AF/FIweginNxCAKzaJ4SJlaosLMgUM2dlCl4ilRSbF3aexYOXh6JSMOsBo1OOnQG
85m7nxHCapELt0No+rNEkJYHPDic90C3fD7x7TXABn1Cu3pU2sQRvmDNXtJbCkaX
zZw9FIYDc4lwz90+mIGVsX699Cf1VC7e5ONtULjJHBy2CleYlhvq+Jl9L787Q4kd
/xEUce9Xa2xiKPTNMOu7PA2q07GWLZa9pcNYaMh46vWxPK2jFzKa7KYLIK59x2Py
HLhOebOPEGhHpzEBPgx5+ih6q4GMRZZ7bgDac9EVOlm9uJ7i0nQFBuUR8uA/769X
+D6dZZhoKNm69coWfIyImFduCQNMK6gTbSpl6ae1x+wKkEqeb6XNnv4P7nSrxHzX
NQpW5dtFKRhFERGek1y+DWfetfAdSAjbEPdtFmODSVpswwRMBNfXR5xi36cic8e8
g7Ny+bRMNXQOlg5G5ObJ5jUVVM0cgTwo7p5RioFAp6Fr8J1shxeQb0zcxmV/ag+E
/cB5raR/CcEOHClZD+nOD4EVooXSXX83y5dodzZJAAAKfTYgX85UuwNQYEBORVXw
H66cANLbyXSKDWMdTFeObIv+IgTTfvbsESAG6Nw34ANkodAsh7Bv0G6E8VjKk7Zy
JxArBAIX8C6z72h7uxO9m6lfQ5m2KAXHmxbpfONH3oML0dnih7oHVlKZDfw1/lID
cwYXoKC2M8BriMD5bkFbjBZ+2KqHcAmcLbMfue4NN/hSo+saa3D1lFtW2R25x4DA
g9ISyHbL/EkWtfPFYWDr9lqroDvRpuOXHQuqfW3IhfLKh+hy8un3EKl3Wl8Q+D+y
5mBKaiBrvFxC5zazZvK7sO72/vnRvk1up/W9LO6hPCtiRk1XV4qflyDu4L85FT64
oxuGoysiS7iRc+HhUzS+Qg0DF6VmQ4erzilrHaiJUmsoM+avY8EXQZfIUwM24h5d
0wfeYi8Zq1s/3GsiiFFsX+Dq58lVaL/6AjSeztFIWVnnvvd2RYO0aIWpGws5t7cK
LsT/GUXtPAXI8m7kZm/sE5mzG59Vp83uC0fRXa1ZeOvQ0WhPh/IbQLhQBIxIrnlm
NcUAZ0ZfmwWnkg/CnhxOMUGGb0Pt58T9235+xPvDc2mRuSYUkYuRDNXlyAjtgfQ2
zL6vu1IgxoMJ1zL7ijDt203X9NaWcj/heo6yaBveTNt6pw8aX3qkTxprSKRxYeZS
ieTkoNxAlP23LgaF9rENqu1E+PqXQg4Bi5+PA+03URCbXFcPYmkgd2VtE0NXkrLM
L5F+MKe7v3CUG9CEX1vXIQyrwXj2TIwNBwrmePJ71BSZiE/CJeN8x3j0CHuQRInA
vjhUaRbJDmUFmFmEoUfJCuZ7LzdrFmDzJMu41f0fEJ37RYW+yKnsIIOBTeZvchZ1
i7w5YQTtR761nsExBvYcsbAEXsbGmeLuepEISFAKBa3l/Chjd9tNtS7EVAht5O1N
nM7MDq56wbRTlc1c0ZNOI0z7PwBMhTikxFKyeV78412wBJAlNAYfwEy3Rzjcpdi6
ud/5K5gMt4G8l9MOf2E6OSRTHr0DC4+FlAkQ3E3vFSkwH+g9x/90tQ4o0CyUj7gu
i2+0Ts6EMry/+GZp6jsuaMEYE/SPHMITeN0oOS00qXFEKNlIOOKyjeuLsRGGtrvt
jtS2GN/ZSqilf6NZN3zuohMm8mZKertrRlfXTnoI8nxNv2k3Oojlol20TMKNI9oY
LKaptU4qPOZDQtoDKU7a81IezDzGTcUxTeV4+Q15j5MRFHmi1UT4xscwAo3vLWRP
7VOMU9Uyk7B/TFgx3v2CQgIQLHls6vGN151ax2gIuK0iq7a1hpZjjxySrBX0Egdo
atHzDzMMxNV5+3vQsDyPpUQH39teyF2ZOQy3YsfkCsG6FGrs+SRSHdph8mfPV44z
/OwWIOe4Qj0Li3qLMSA9YpvELx+LuS4S7RwSyqKMGV8nFacC1h7XK/DdzdILjmqD
T8kguMvpyBUzbwcZZrcmQe/3NTBNDK6NvlCTfFibdXjR6Bq4xHhMgQKNd4wqPdn0
fkcJorjoPTXYpe8ZGKPxHJlNUNOavN022ILl0q803HPNM/V9ftt7edW60Y7MUfUW
eazyuDpUyFlJOB+gBPKqBDHE/CbQXI/z5jHb/MCxxezdd71wx5VFOxQETZVg4d5H
0pLys1583C385+6vLiJUT0Qlz+v3RNavX5U7cV2TXADm5BDbe+Q8uwl8L/9UCrOd
JBb9tLwnW7W3R9OLYcmlXYe5fU/lbJd8gOHG+u8fxdHD+9CW93eSBQUEx3nQ7aUz
J91P9OGYOs9Dz2YclkOkLXYGPb/Wjx7KB7js019+qQH/7mbwvE3E8JrG9JPvzBoI
9oV9y7lUTBP9FCL0k1Bejsn+ELBiuLCPMWZ/z9mvv1TCrtUAvdCNtEBPA151prDD
bzv6nu2fW74xFmTq1DI1Ms/eaEwQPHC5RCHtQN6WeKxQuFsOD4DsuJ8SK9WIGRI/
moxOgeaShQ0qGVu6n+1wjomtp/gxNxu81uqQDfrATrabgaLe9H3ynO1NVLwocgY0
GD8mylji0p6CqUKaAE71mu6AqQkiWaDO571QcQYfzOQFAZsLCzcfdy4gyhHksRfG
bR1uD1PiblhitEvV+TwCUTl01xyDK3ZqyP0RHUD3b5Z1YWinHsWOUn37dQELZ13z
T0y4BRV87iq+nJgVq+hanmpcTBjUFvzW0OPZZg8E4m6j96xe2QtSiwrI2CCs2tim
QddZHjIu2xF2HWl3pKhkxNEqFx3hbuQ6I73aHVBO0h45Wa5wVg65ObNaoqjlLoR/
bPFqfjvQBtKiY5S4TUuxafYD2jK0k1jeWp1ktBZMboDogVgoDIojyZXjk0CCwNdy
ygJP3cCmOkxB/dXUXl0C/dprw7WmaVgyY/PtYppjDXjppn897gZyRUCcJ6qMDKTs
SoZlFzrZbNNzeZHrXeSRSktwNZEm9rhEc5R5kkYFpFKNeO/sW/WG7hjVkPzyAQPb
uj7s3ZHDkYOXokhRoeZuvN2CNVwjNW1fp9neoTc2DlWChHs8z1g1L7NHnFVdAldI
1ZuuR4oM7FsTp3wCOObMS8uhLnf061NVgTpZsBGwX/9BUlyj3fQ65rvIMh4OLVyM
HekkLbCMU/mzCPBEEZouXsS9CoWMcBYhiqCfKiPFJ1+lv/s26UxabfThDev5FpNp
1J0IyQxiRv4suh0JsO5Uy+/GhMyvZfx99Heq2VuFdwl9+WsthncCzPJwqy1QlIWQ
PTd8ClxHUbPQe+djVntc7SzURN74iKiixwBbtR/MpHsiQCvEDzCOAWoYraaniAGi
D+9a1206mSTqZ5q+wp34J7Z0GX5pOxQlNJxYqH8+RAIkRoauAI5zgLFPmejCxUnM
hCe7npsCj5mx3hyG2bvltw8wYrQOFIWL2th7MJnDK3qBfdyf2NgCnto2C85gpQ0M
O7wVw/FUCo3l8t451cHU3hn2PrD4o8Qudkr0Mnu62QIgzo25dx4BvIwqKwarG4nf
xpuC0LFL8ANC8VNo2v6MNMwFnhQtI6mTK0y15B1PBsYAzRRdOJGG6OiDHX08zsbA
HkXYd5FGmbIA+m1kIezefsTUFhe4Vm0pWQ3s2YpyTvLGyck7S0AGHJzPcHOnaLWy
y16MvFPbEYIlAnSSSqgYg7TMZcv7foukvQi3751S/XeVbQCvAO87RiIqtraA8EJo
QZK1X3INRXhViImPxd5EsXpV7DRB1NGUy+gJ7KAn0xNwiJ9Pxo3oR0D/gk8hXJMC
MuurmKJumV06hRR0huxN6EP0ujPLsUwcZKiuNl3JTbjTnLF84C76k+pTesyjWLiw
YMyYgmBwGgBU5BH4/DFssq7GRR2Br0cup8Qf90+0S4TqIT66cEgfNvAxKhNGowiO
OHm3Cu9I4YysHuDR9983TY6TJL87oqsoeBCritpG4dn7ZMWp6w1RNy2I9kXamsML
nZiCevatfF7n4Ows74L5SfIoL4vjGNoShrkML+dwgMlwmy65BqzeOSs+piPIgNCw
N9YqgLxQtCyuSvgLv2GXuQrCOlGvVGH1YbG/2vEHiACtu8eyEuxtkqu0klj5cj95
O0ef6/AP6ubeRoT5QzarapWgWHh+ByMb7GQ+VKlknzlMwiPenUGiYshU9P0SjLJ2
gBNyyc3qMrUyjNW1tKjFun7qaTIqoM/0USAQfcX00uzukSZXowfdvLYdaD0GkO2V
Yg4lCGtsJeSx6vAPOzrl7ALSN8ACugMIKRbxlf615cZmu0AX9H9Rj3CVKuQNgZvG
yiSVYpgpk1QnIcIDDpRRK/Mhnu2uu5vfaEQ33z6r09Rr6F4wqbGynNPPypshDxoX
Ml9ZVaxeryxhLz+aUse0eFLdYCyNUYeNz8PEsPR6HDmnSERridivCbrRdRveFENC
3QhOXfBnBpQ+kTj5P+UL8Bsj64pto74z/IIwxeA7ns8ZJ0xCUSOpNJRLcD0TDiIY
Al2fi5J5/DYgpWKKeY2NU+XR9dAb2f2H5DDN7v3ELxP2UCZJV6ZU/UusJd2YMrYR
9LsHJN/EzQCOFbeLiumRnQaHzEBl5Efjkimd4x+RCaFU/49+T3AyluRQj0PUHo9+
t3OapPbcBAbm17bqJPh6TyzsHx+JIivZexlFEKQKZ+MWknOBN1utvdW4Xb+s3xLT
6FbGxaGBhmUbk0wYexIjbj30P6abgCcDuOerL7uxk3AtQ29e43Vg+BemnStiiVSF
jcZHYQnnuaps0iBVRmW7+/mxwIZhjYE67zVYgMS5ZAGylaExYImwzRDcq5cG/guc
z/glTGrMX9+OnzAhm1zgb5G1vb7+SN+PRX7caOHUa0HcNLVY4OMO2Btip2h2ToiP
u69MkDdqWfqlBUuSfgPcHQofzBn8BPtLNhCYSg0mjNeqNtEEE4ttaHekbOucKHGL
Ov8g3BCWpOdy1DONDdsumsxNi7prT8hvnNI/LSSJs84Npdaaf3cClRwWq9wwBZ2Q
k5lNP9jyggkcbv/x69IYj1Pkq1kbIGgrN2fu6eDrgpDhVKkBgPm9AUmaafJG+ikw
VSZ51xAM5Uiml3rXJ+orTj833FDLEAXIzYF2YAp/QQkSCXflbSCqmXcmjtNO7+ae
qgfLS+uBaQ9j5vNE3wDsbDozYjhPRVV/A3fYaurLx33kNm+8ThTzqbYLIaT4MMVJ
INIhPfk11hvV6UFkWl1i6unF4wjKacMICouWt233/ii3woQmPtlmdXM31Na/3T2O
wniE6XtZfXXcWYCih90BqI8wLo6XMexo9kCZyb3stfgLBypHO9OEfyxrT55vvAMb
9TVVqLSiXeYGQafRjYRf4ExgEdnLfrUtbGoa+8DTnmFeJ0zNvfMcWiLh2Y45pdhu
MJC8upAqNUTIbm6/krA8F1fOFzf7Fq0WatQwcEb9SVoRFT3leiTD1lrooMKdU6Zj
RoN+fuLP6+Z7Mlius+zBSdmaXiRWePfWQUiNd/m4BYtElzeykQUmG+Ztp64MSZht
YybEW7+t2HLMKWX3ZV7bPrXm6/vJcncaWZJQ+ktMcyQzLYAqZPSFjcu6Dc4Pngwl
cyLJXd6ExK2wfOXEjtoiiT7SHzKkMpYlFFJwwXPj9hOa+qc82jch2i8BBdkJaJZJ
+oudsQHEOJQBwbKJsx+2c0sKqRwBbVoQrCbG9DKL/f3Vn0UOBTLY/cg2QPUYaR9v
kB6qD8Rbp5gZ1HNb/WO8Cr66gBD2Xj1fxiHtPjY5yfaWc0VRpVlIdO4nq7bok+co
oeHYxJuz0M1XQnlXsxfyE56YrgXl1DgskOo0bvsC3+LKDEP0l7vWr+vGU5dvhX85
szurgg5UhBntumwnmwdnNEk63Pz2CS5RK4Z3G8c2kQDg6O6tY+ZSyB0UkOIjQwvd
AzUTTt6f20VtlZMxvfMkOeaKs9d2+Kd24904xaBlqlVbnaL7+OVNxcQVHB9XP4ab
a7NP/LzgUJgjAb3Sjt88o3Qx8BfjpyGkm6j2R6bFgRiPwR+Ug5YXuZppw8kSdRyK
JB1FC82fCXH2XhlTIb3VIJw/G+Qqflpw/tSNMBhLXen26ex3EswG5n5DzmvGtu9G
p0D1kE6mGzrPNmhPGq54GdR1ExGtUVqBKIKDOvg2I4cqoSTiJBi42ou9y3QmeybB
Z4esJnIm2KRMCWeZlCitcpsCmW0Q575KZtuw+TYejkAj+CacumwpjaAFQZNI+BHJ
GNoR67hDqIfJmmY4QW/KKHuVkPJ8Pb7XJLRskqHAPZG+nHWXLB2ktk8LAGO23x8E
uuYey8jaRzXDD6zHvvWbrGi6wTnrEXyZAT0nw+wCCXqnkm10YUw+5lrtBB4fRx2A
lpmCeRYmDxO2pa9YJmK29da3TwOpiLonkLmunTtZeHMvdVaxNJsm+oD3/ozjoSrq
+94qh9vgG2QQLu/syO5pnSiPIUxoA8CL5DTQv2EDmbxFJWsVj2B0kFNqORxG+A6w
LBUBQJ6kQ2CG9f67KAsdMZYjzzar6jSaroCNPb8hbjQr6OWqU6eiZHdBIMSwi9BT
IyInNH+0jAYvHGSFt2vC2B3hwfFeq1SqYvhIVMLakec2HR/VcHJ9zE2wctx30skR
Zcpx6ZZViCpbEPcGCnxJFHeJ1VCVQPzIlvOaKrAMwEnceYD05loIvw6SNje8yrnD
osDAD5d9nLQqKvM7KXTnCSmr15XGLWOZMg8kdNqhRO6Mw7RYjsV57jxuNhxwPlXr
wb2piKSZK/cxhJKLV+vHzJ3nBvB7CgynR3Pwj7qzpT3rFCixEVluC4JE0Vavevw/
9l5uy223dWJiZNcHAaygVjgyX/lhXILnetwi4SEh/V4j9kVl0bYhiONcLI5eZc/X
dvOkbYIZWfYTL3EBwSy6KIrxrqaihb8Z4rZSAlBK6d06r60AN5RjM+FAeq/cB+o2
h0bI0TCaZi8Tu3VzqZqyi/15f7jsrQacXrRf3W71T/ql7Im0xyfrXL2UfcN5+psC
oHKI9IDu/KUayFduk2IDzn8oH8Xms00KEwVUR9wuSsJklclFGHj5ilWB/ojjalkC
m3UdySR+LHdVplxw/QW9CmuTZGpE6k6uEqaf3rW+JMISrStlqDNqmCUdDnpH5LW6
IY3QNlq+emqWa/V3L6ekob3/w8CGmI3Ew78qJENBtoj4DAUUbMOVCLehUCwPBpyc
tFSqDOScHHId+YILpgv0reH9uewQdymlCaamvfJfSxktXpm8kyj+QfZBj1LB4izK
Q//uX/Y0szFdUMeXOTz7Ii+lzYOQycNWoKKwlx2IdFwxcda0JbdS5HHPmOY+s73O
EGuScI4+Ex3hawy4cMoQCWoF47YECeK1jo+C3kxVM+DnHzuFr1TVnmFeBQschkSv
Rde0V6SCBJM5ROYbSlcDjjrVrs6AwytnCqzoNa8AJ0EL1Nvjrw+XC59JxqGAIs/E
30tQi5Wx9pQH6hmCxs0aWeMFgQe6kRTRDliofj8zv2lbE3CVFgTfF+T/Am88i/Tt
gepUiC1qBLafKY7gINl81CI/auZulVSww2xo96DPCkW2QjXEpBcv0QHc8iKulM01
Mx4X9sVj+bi7qeKRP5Y55nezUg7oQy00+zVaSpt0fmHqXaFY6UW8ZpgCp1hOm7Kx
TUQJaYuyiZPomDdokiDDkIHWQ3EXNjKxSZrQorhxH4Sby1xyBjEFAjE4Yd5IFlJp
7iYKEi+SZ4YKfO7x8j5MTG+ML0O9vyXAEHwXv182XzDUE0N7PWpss3z/fhTZ08Ud
XQPf7G6RKTwKi/T3en4R9uhETbPfgeeKqwECmw4ORbkf6W9fAX94zR5vtA8oMOXg
vAvCA0AoViBNWcN9Oe6p4jLtCI7K1vL++0ghD6MLgub7/J6c46EBadP4nai9mO9M
df5eBQhzIGTkFzMBVDbGdwHFF4HnC/61fh3VTenCiQxmkbuUHwdQ7xzq7hqXz3Uf
tw6X9CJ+CbXLPnxPa9QCiYqlcTBBiA0WcV0bVv1iS+5lGWSsk6ywlWHinxfrpupu
qQUod35E2FyXFb7q8lgcb1tg3FQa+BPOlGe2bqm/nVbUuvmQQK1qYeov9hEoBq6k
6yzYYOem1t9rebOsWapj2JmczxLq1lTTQvbMWXQo882muzfQfTmPP+gu8B8YbBPu
XZ9VS5xb9ibUV6WjW6PMwTzo8SlcZazpAy3SgBtLiPAtW44enw9gDwz31yTQl8JI
2kGBr52eIiDf9X1gVCw7/tZ14xLTLCyny6y+VW6XTbSTvmfn7Vb869MzNb7F3Ul5
DcB1Q5Vs2LKsZWfui9OicoykvSy5mv3i05Uaziy2kNlF/Rx9piN6vB27GWkaOnx/
CJ1jCV3bHvlTe7pWkpIBDf9Samfb3uWN5xvi0KYlnDUhbqLoTdWPwgy3fyzDkJKj
+qE9h6HJym/RMQHrtbZY0F+lk6nMzW5SYTHq6Rft2NfofOx8NK3t3mg4kaROPjGh
U4PgzFHFW4AGvT+r7cNz3wSfGuKM6LjJHLgtxEOFAxgj31iWPkWGs+SYfRlKlATY
IsWpCrPMUcS1vUNNHyaUObhi2VnSFYSllOR35pKLMpUj4yOC9LUyrFIQ8Y1T0fGa
vXGEOKjed49X8SrUZvqQEk3++1Jp/bT+WuOB9H53L/sT08N69VKfvqgb72fvNrsY
iwNV0tegDecD8JYDAn3DuhlYMLF2mLzpw3ytcc6vKKgvd8d2rYXusE0aukJpQbZK
ov16dQdd9UqLDz240Bat6EIg0OeD8lUtos5dRbqu0f7wtqizR9nQmrr4/raUAgNs
zWwbn0snT963m4Nso9a7wqFn4AwiapIEmHzaQbwDGozeStUPFARMnZxDG0Pe4xvy
aZxCsXlSoo2l4j2ePbmT40JuS5yqUyCvRhMBe32OQhiQvritYUnOwvyqSoxSOkqZ
PNszznHViJ0nOxT7Wyrk4/o0FrC6xQ8w67cDQgZ3Bb72WO3ppiI+wy503tS4roIh
9+8Ac+c9MjVU0O3PtrwuNbpTpfwlhbEu0BR4UIJUy3zXoIu9+Kd+znQO63XSJMxT
TYe+mnxA4hXj73lmXr7kFK12mtI6p5/NzhrGGVFt/of/PWJbAYzHENfbgkGFSuAS
wESFCMbOw2A7th5xrQWUabn4yOEudtV6c8P3N+8BYaO+TsQ0ZZXxI0EXLyXM0WwI
MX8LcRe9gl9ZKOuC4ecEvbqwnwEoeZkSQzmGmCudd7m65mITB42ptGK3fGzWGiiX
kBqbWKBDUs1N/MSZuBFOTRyhj+tNNGI5Y3svZpCcQ8O6NOU2QgUJ0Mj+F7PQYOWs
VL4y/lsyJFcb4oFN5lmEne8kWVjSIkyNcwu/Oepc6up8IaDdvcWRe38p5ky6YBa0
jSxAJLsKa7X49SodGBnxXKSXEs7QEsd1FwbQCTkKf+Nd73JfGkPXyw+RRsGeKS4S
mJRyK+9fmk1PDPYlpkFVGT7r87KMXfb8BCXd4oFTaapy/PhSkJ/u3q+LrneRkxcT
xHuOnGeGf5dN65ap7HKBxgyRzZk8x9LZ5PsZf2l3C6ZLaBlc8rOd4h2x5YuSTWEF
AEXgZ/M5YglCa8u+zzm5qtbcqZvAC35Ps+Y/Aa/560d0cKXcW/epkzJ5Li/2Q9G3
LM+zhrj8ZCGcHICYk7D6SgecJenSvmOPfSOclDpn4cUHTklb6EZHEa2OZQvhmJtm
ABKB0bYUeBQNcpjzSJQZFshHlDnPfXaQqcIEolNW3k2q/4/37MLTVQMy1DON1iGO
uaYu03GtHAOz5dLtrD5dM19JSVFxXo/Dej8ipYA3zWuisgL0zZpvaBaTibR6asXv
nPoRoF2sWC/v+dqGyYUnK8/EJQXs1LeIgvEUsIvhfmBPaC8vDwAOa1ZNLBIsj6y4
mkUKjhdx0ULu4EkVF0ezOMxpJ5ZQGrgZOMgDQj8tohOD3uX4NXw+IQYgJCxwGWIp
LdEyTNl8Y6o06q+/1FgOu78Z3fQZkzJCpfUCqXwV/7r9+lkTiS62iFk3G7AzHCI0
EZ6v9AB4zQiEvZ0657xOs6/jhUDonWpIRdKavVCBHsnFyhy+Cj0+CvFJ1p0M6EL9
b2ti1dsru8TW1m4smPqI6NB+RYLSxrVxAbuC7r9Md8e9ynbGLRNiIzRDa40U9fR+
Yul/MyGgUoNlWpPa6Pg3U/TYxTWjNQQi4NbRu5XzB/8iUrc10dnw2uMmvD3aHycR
0/EKNixg6C0+PffxymrmPkQEfAfT7ATys/twdrYw31SdC7CsTY9Ab1BQrlyjUMwM
eR+awzXtPVwLPb8Hh1NQTXkctiDHoOXTXd5xt/AZeiKJIW9VPmIp/23iiyqGrakV
Yn7jBcb0HbolfGFs6gPrx5IIeElAohbFf22uobmbCZuNkY84MP+iuAjLBtIGBw5k
hclU9pN156lp+ExWuNAaW2gKBBlSLQBk94zMVejJS3+2Swwe+Gd7jCzymDJPhYq4
4MbEvVWD5Y3dqKuDSAzoiMBVl0SuNQqlvTS6ga+NxXcAKpP1FVfsVNqH03lczqlg
8dmtPEWQjAXIRjMGGrkAiKncGkd9jXCXStIoKKcpF7F3gymErmL5vn39VeOSXsBk
u5aas9Oqu4QAr2rmFSIqjgQGwig54PQ3QNdLvup5HFfexkAecmihtMawCVH5z4hf
AmIXhcWcH9zK9z7BSwI1C2r9ungWM6iq3ZmxRXsY80JGuZ8Fd+4CqaGmG7JhI3ZF
ytrDK12aUWjyMFCeAc9pdl5X1bkQzHUt1R/7n+t6jfuVZWNYkDUgAfTKLkE8xdTC
lMARqzrpkEDB4yHrx0xOQSdJ3NL7qaYHJXAWkeCJuTWUWFbNk2x3FXMD/2FTudiY
WVtTalw/hyZSEMd374fLzE5LeDBMlcAe4aJtu+mGQOotgOJNtSWgWFcBQQ01HT9l
xroS2OW6N3fsGFcki3b/+90OUGbGiar/8TMNgFoCCigf74YURnygVTnCr9Wy95rR
0Lu/pTjku4WTqg0ocnYDQ1xA45WEtT9Zd66jev/mQtclg+73h97SKN4CY8ywgJD/
aQqkmqjQp4yQGAAhJYS4c58pr6SC4D9q6WlVi/C1ivWIwqxgGNd4TDNv//lHXO8Q
bVXwvGxR1x70HQ09buj7T/1+9lE7hLXDiepgR7fk0tN4ZcdQsMFZCTl64+ChXfHs
n3FEFVpXY7boF4vKz8kZeoZjc4cSH4pwf7mckM5B4YHsN3E0OxkRV7r5+dBsCJHM
YQtjz1IEqmLWRq36k+76XRdkIKSbrR4K1tdkNO2OV3nz90BbqqNwBDoj7+b9HmrQ
/2ChKdPhV6dVjHhobWxdYQsen60+c4TTEYNIB1DHvfBXT04Dxh1hthq4s9A0eSKI
BJKDYJHrF6UiT82SrHRTntxSKqRK/plroQ73LTWMI1U6D/WJYuveTesefIaArL+b
MLuj+xmYb1DGAzWFzyaKQsX4qFkxq/mgpFdf6b8RCvzpuHut1DA2LoOxxAJ0QBB7
Qr8YLs8GHgsvnfz09IvnnxBRn8BuzAcqUgq6zmRQGMhMhD5qR8dB2Qc7sIuD2Co9
qWqGXyvkdiA4eq3VDquJ8AqddS647VuIup6dgpGILG+So2CBkMh0DINaKkOXBeFf
4C9jVvb+MbxipmOI3MKHOqa9SrBVVnNZsqpsYXcv0S7SOabHiFZjTiKnwyReBNgz
hMA8Edy02HvMCEDNC4vOa8loKzmhdns4813UYQhuwQnNVdo2yq5VH4oJz3YyKKF4
blMNvNUthoH9FR+0N+9+edZwW3V7yCXyB2h1mI6ICDaNhEtyQNwelJl9nBpJKNc1
ZYOcOk4sjU8pG7Ms+D8c2VUJuFBn3aaXch0pqJPd2hck/U7cT1yZXVZQADXY9ZuC
8Rid6iF0nbs5HG6cCEE+4+wDFBvrHHVhVVg9Td4Iutqe8QoExrvSk5v/x81YhZ4b
VZ3+9ONgnZwHjVPR0ZqhvOO1sKsRvHeVsMyHhPANQNSfY6kMuvrntxQA07OkX0W0
XzzlB6we3mI8YojLb8tky2NrM9ldgVYxxrqdD3MffTKi2O2+1kvTIvPsZyACVexe
dWQ3OGTOV8jf/jbYuW96uycsQC0aG549ajt9wjFa+yrgxxa/4UocfDyx5WkaOBji
RzPQ8go70wPH7OAYijQAV02D7UAR7NNQlrDyQAVbJAiYHVcY4GuiHSnIiQ/R2Ksv
Ekzm2HiYWgVyaU0PAQrZEujWwp0zzVmDIvWtKfKnad80yLZo8O91rWa/g2jGBERt
2vdWEx6DkQ4ThSyAtWsqU7WnDpCkiN7C/UY2KNUGP3TkWihXgw7Xv2zTA9Qr5VpO
/PKP9az8bNpu7jgOgHEXIiAlhpU3XmytiUMoAM2D06McDXID8fWxUObYNHf4OpFG
GNK2TRJSPJfxEi9JWjhlGokbbXh1rO13uH6bChdECYNvXHfe4xWMSEvaZIKAbf8n
cjQ76GJxFhdPdee3MtN80WB4BBnwpQc+iqtXtf8VQv4Uh0C5p6m3vrLC1OcMYqGH
8FH+y7aqKo277yLx+FWtla3rtuo8W7lZLEjQ7pDPTxy2dbgQpevHL051YMV/J2Im
ix65FR+ZRkdos2R1ipBs8UGvKUTH7DXydWkk8y6GDIcaZSxuYqyX7t6pqtIEK7Vj
tv2OrA38ilpbc1fAUAc8BRO5UKbM4mnGMoX4LEpVrIgX4O1zbyxRGw7gb/jATFWe
4srWp/dqCqEl+bIJZLAQpKtUC8XwdJgcozdmppU3YyxHM/AzL4whreL5jNgoQtxE
Si9vcFOK6sor1l3b9f4KtnYoi6TBtzsszd76krVRzwK/X6tSZ1JKQ++zqmVDfM2Y
BdvX/uTypwCpK/RxQBeNytavj0b0dyhvfAaqmXfKZRVwpY0OwzHeof4PcbwqTIVo
FCudGh3Vvg7PRUA/+HHPOxZxph3qzr/7oJEoT90FY6SOd2A5kuTHXCI5wdYRVXed
p2iokDudZTLfcIRFptoQ8qegcB+PpnxNnBRWtx+cw++kUwuLDhWvQrbiVcremR/1
HJvKodHGzHIeiw8jCBWddgRU8xHC5JxWbIP9wJVZ5tmHuB9xZjieunPCsJLim8ZL
AIesOUZoDjzfLH8d0l3NNxUFKn/2E3J+lJuOOK0tJo3qbD0bGuuP0W1TVufeFIHW
+gzHZQD6sYZlugSGDSPnAMh1Ixpsf+k9AuXgqrMHfMBQUhnntv+53f1rEuL1I26R
fyJGw6m6QcZN/YUbGJqh7d8guLNDcyJg0deOchJSXcjqJoa2gku9owlMGmzZq9o6
UG0PowKfm2QeULbFBvvASNkMyainiLxLVKF3gYUB6QRuL72ue8OKGXvHACBswuDb
uYr+2TUPuyOx96FImHGmkwyt2OykT9rZ9mdqMBC88iRXJ/oXVg9e98To9y2RqvKE
YMPae9x0xHBrPzuLV8e4P4lrcC6OmX+C2gsozQo5U+nx31C2W9Qut+AITlQHxCQH
+v2WILJOZYP0UJzVvGG9Ecju5IbD3cBKSyu9rM8/14IOODlyp91Ryq77X6G6m9g4
nSU8X4xvS4JGOfurT2z6KSnweei1fLZ1Pj5LKp+4LUpgTTHGcIqfgYJJMgteI2i5
X1EsEJpRghzRoUs+psQmyI5nUSWRd6cvEwO+H3SvRcLU7Zh6jLi9pokoGBR2cflu
TD3ZKOhXZx+oTAPrugNRkpv6HPjM+Muz5j4vyWG0T8H2LXt/JIXTZeZQSD7PaM0Y
mgvXjPVAJtQaOSGJR9H1pBcRuE5BRo20cfZdZX+iW53wXHtki2aupNvH6ppmGapf
CO681LGTqF18sDpHfDktcgE9AIy4dvdYZjpI34IP3Uvi8Z5FDKIVWPCcNn8wF//p
zVFQeA7LRrTqN/qyG/KWactM44/dU/nCFqks9TXeGKW+Z6w+B5rBGt0ARVU2R5Rt
crvYnbMbSUJ0Gbqa0LZbFYSRBnE7eHNQcf/8noWpAF4e1mx9mnrerrPyAdX84bss
HVveuJPqWbcJL8HeaCJeanpf4PXGsHrDBU18J5SY17KkircVkOFW50cKvvLn5ftN
oFadI5N/JWCLsp3XUPoiwkqL0UrabLykRxcwP9f8MN/sLspDySek/22ZrnqsfQNR
x+oZXdJmlZepVhIaZ7bYn11p6L6K83/OwbtvNbbLlD8HwJUdDf9oElaQzwIou7TW
1BqQMSRi2y3LWB9ScYl4k7TCs4t7CopbPOurO3HmuJRnZ1DDfSKmwMhEKNxZ6tuJ
j25IVgHFQPSRKBPS0e8wIoVZjU8nX02zpp+6nZOPc+wFGXtp0FL2/MkWZHUGtvGU
17oxX4mG8Bp9N5l88eox0Z1S+8gCI49gj+OmawkZy22HdTWXkIZnOXd8rcdElDlK
0f4x2IJNnSDUjjdWYH9OvZXkCuZ9Kf6OnIFkwNEQnIstjkND+tH1wbP71U6FkGF4
9G8wbH2P4kBJoj30Ibso8HEE3qmNVqb+zpUU0L22XjNW4mwg+buGhYcM4nZxO3ia
DzOTl6v39r5WEpj6IQ6KhtPLw5lT6q4SaIQNwXJMid7jPFMAh8nUIyMkx3kmyEvs
oB5ESNhDT1FPjJakvsG5aH2EFH5QsALAre3/ijP+LlLLBhAPI3vHuo68fiIHe1qi
b85zvQKdERjQtJN88hJ6sbfve93e4HA4mTkbmI8i1MSBiLpcwRu7kBLYirPWhHfs
cUIv4wVy+OXTOUbxVE4qvZbzafUObrfSVctBAi120gXKOJ3NtkTCmRTP/fwCHWSY
xarnhLiqCmtL8N5obGTP/t/HbU/lTkeYB/PwUU5g2i052Wlj2oa3w5W1UDT4GRZR
u7XojqnrMJq5ZvutoO6Yrk4EPRxrA0ka/hJJnzAjTU0mCZ+ANTVcQdArSG9VM46Z
RgrjokPs7GISNqTrqX6EN1pCcxrLaJtDazx/4xi50Tuj1iXv4SA4e6jeBi7YssVM
m/Vgy7BwyETBYsm7RfqcLtFD0xzAa992fwq/HWGehWkJ5CQyHjfVss0we7ZX22zT
zKzjcv+hQxfTbjEG+MAu7/l/J1nR+nHrXTPSBL1pmEdXkdUnsQQpa0wUzorOhehe
g5lkr//+GheseOs7atFqP/XMeE9zaPaZNf4SYPya9nmh6RauusDlvU/TQctWHXye
CvfdBrXA2/fl2bhsNCHBeJ5vAvFjJtZw1IMo05BVP+EiXZKDc89upJOU0PZJiihD
LMWGX6vhjJQ2ALWPhq3PhNAsQsCgyqlpR/wlecj+9EmB+p5y4mXZMYO0o+c6Mg5Z
gmhERVHy3RDzA89fh6StejwAGzFK6TM2jBaucd2IvIGFMf46ilI2PMZMuWeBJNkZ
gtfvikc0U/p/IEHS/ucSFFwp5iGGnXJShI4TfySPIMzg/fhMxzrx/uVau/CBD/9s
r+W7H8JrryQhesOEe9W0s2V0B8Q22WT7tp35aQR2QjIuWvavLTYP5k6qY0qLagH9
PJ9Dt8QEdY9alNVtudqYovw72htndzdoqSbPVKTeZKHN/w+qyCVvtkMzSl2MQ5o6
jggXaNe+7sLudIS//uOlCdIvyQZo2nrczYf+l0lrMQxfgtCPJXlAdIrWUhhVkh/p
1KSVmz1f7bu48SOkFoNh5EfZapuU9ZAiD02NQ1pxYrH+SFfKcHBZ1sRiW0sZgngk
jHf8cL7sC+zHFZSdUY3ql1qVtqtsLUYpY7HLsxORVO77rQBmZgGFb/bQqAbtCkNW
3ET1L1ZiIBVmJf9ayxIp6FxuXlgjohlJdBgUmXz/71KgORB+seJ6Wcs+vZ4NC2Vp
KlbebGWYViTTSpeGmi4UZT9xpBOkj+jRp9R+OxtlY46ubwNqkTIb/7KRoNmnP7jR
9SEWjkMjOfN0JCS+QRM6XCTJb/tL26VbYOdL97ngC3REn5gQ59UjXncDW41iS+1O
lJrP3eQ7IkzaLS05Cp3HTE6X3aN0QDQKpTM93U39rw+MShyLgHcJmtUF9r6ntcyz
sTwODKFV1jIhJUWd00DtP/Lfw1dwHnK8Al4RrO1JN3OQ5wVslH9TqLX/bRzlWi8o
2IJlTSgrsdLXTj5eng1+3HNJ/NLDBREN9wD5n9epR8+KluU+cw98/7qjxZAbPSz4
MdRIXy6DzkJKXLV/xYbftmATz/pyh/ROLKsv8J1Gkf+tmgntVqASqFWyKPorvSGW
lifb9oCoc4dyPKEZwZ3Oeg/R3/hNE4JqwFsS3NJI7um9AgyswONQVMj0SZVrksTk
Vef46X2aCYOybeCPob4Z5THcilvTMFPeaxoifX6bWwZjIBQ12ehwAoZmuDLl3Gd6
XtmnQA4J0n8FHHPVCrGSZrGaYPEP3Mk9PHo1cc53OxMvozl4Vwg2GyGC9h8ScwFI
wfhyLRUyTFvf9PeuhkNuD0j5st9IJ9T3jHn4e/0r/M6+imjQfclEYqNktkV2WPOS
szDF2pS327T3vTAisEIpDopoO5yd2s1D8jKvghGXkbPVq8iePdIPtqRgkJnVrn2X
qjaSqq7rECV5ZBHFzEqIgoNvDfA38yVg3BOOmJ2q6B806DGGFzieM/pSHFgSWIlN
S1o3hWmA7Mui680uqQF1Krqds7CRzoJJ9AkHGpd3RFNbKrOxLt45xIyo9R1FowwU
V/Z8e07xyHMW8yMdg/OEMQOjQRhlqIWn/hPR+G7u5lsu/sOM4+znVlH3icZ4+VT+
ucheZP10ydVd0At3xjrP9s/o798muPJxjFCute6lkYy0mQaO1VZwFcHXUbJlazIp
ev9pK2/n6gK4Z289bm736CbPtKmFE9nNh0vZRPu8s0ihyXcPR3hPiSQ4IwJpvjT9
aBz5tTNRTKhFieDsLN+/XzS1U6ObO649/Yp32hNdkWxHtKC0MZHIDAhUAup0cPRl
PMxgGeqaW1NR73sMKUcmCOpcA+6lo0QkrXYnB9kYPnOf529p+JIa5FAx6egfKnBF
Tn9Mpy+hoy4OgG3AU25CRCKZnoryYQDl/W/07B7vgFXkno0xuzFu5TZvh51EQ8ru
l18xTPW6bJPGf46WMTwYoonHt2kp6elCTON2Dd+yhliLTqBcSWW/sQ2EKW3VxZd6
0u0X133la/R4pwFPYQqDcd0W9uf0pES++CAf6SHIuHXJDSNeXyhZSqeJqGVZ0ULW
FCK5xQDNECiYXcVIgTcJ1RuKBz4ZawRyvIzse76aEo6dxa9MQBaj3kdd3TJHTm6C
qJ8YjncjkNSD6D7E/WGlGAbspn0/op8wkYkGqw9COhKUV3mP7wbj/2DtXgGff2dl
GnAfH2X/naYl30q5O+6/WU3ufrU2l8+fPMLe5lL+VBTnlX/K6wUA9QLIKUWDtU7f
+6rpTKlI8IXlOBdTKQVGnKg85wG41l4q757c+loyotKjToSBKTI49kodGc4G/K+h
EELrXrmYFw5jKj1v40z+yKepQ6XZOiEWDzBSgnsoh391WtD0JR3RTYN3/hhkbdRH
QMpV4uJYJowvuYdGgLcEYWVAESV0jVxs49hrpdU29G084giCkaXYuGbuauOGvsfd
cuoLmfuibT+2dpLzbjAPhn3PU8qAUC1ILAC0yETFqaT2rLscg1IkVJ/fARk/PHwE
sT/jiZ1mKWXpucifDXc52oM8LPwvsOHVoLB3rt1N21Aq7IjvKK+2/qleDH6mkqeW
vcrd3WKzDWte6srVwH/XkpROoY1WdOt1lz0/jlaGXaB90u6FvCilrAFY0h3EneRO
S0WsGMUPZXa2NmknJpiTr/jFeaF/x98p/145DZ4Al4withb11Vgpklu19HCyFhlE
jnb2qRsASMV3lrWeI9MPGZx/y6s57zVneC5zMTaaTUpWoaysxr4POKrwa1s4713c
uYrZZ/jViFT+m1EghKjYspmO8b8kmy7bDixiZEcD4OTD+8bHq0fihGnfFmC8NdpK
mVY6MU0t+QwmkheXd8gnpq0anzR8Copxm/JdV4c33/v8wx2GHCSt8OaO/clLM1yi
ch+XXMF3p1lqeJgNAx4egb/gxD9mNiOi+H7Li3nuwPYU6OKrQXsj4Bzqev6+LcmB
INk+oszx3k30RtVxnBE5lXcJwoSL+khZMrMc1KMTXzCx5kdmTqcFmiCwbO7FiWdL
xRXLD9yclmGKS6dA1yp/cwq8pRj4Ql46mErKryCeFfTvP5M4SZ7BpUeEzhnuyTrg
gn+fYC9+BGaSr/H5kOCGGU6V1OiQbIP+e2HFu8bDO8hBATBBV1uwDnXroplwnFU7
+xdr4+qRtpfqkFcNpfjvZQGd137N74mgoNxa/hL2Z1/kcFeddKolDC5c4rhoTrMV
jD1G1ZaHo30gPh/7QeHjPtKTDPlHEZFGEMijF4r4uYk8lYW0QY/YTzy9gxvt3M4B
a473y0Mvo76z9MY/6IYrFfTIWcnsc1lfm35HnLWZrdkRcTEV1TJ3UiP51sVtlxZf
eYL2hRryA76jSQZHkbmsNsChKYzkBRTClqt/asBYGwxPe8vyF6roIXu15SHjHcGm
wAHmC/CyVmGlm+9/Avh1dRkzg5B0Jzeu+DFbuyy9y0X9waQbFd2wq44ElQWgk+D7
ySZEC15Q2jrhLNnLHaKhROFussCH5X6rqoui2+4E/DZGFrUqjuFs/7Ce0woxKPts
XNS9/dwBBHn1wf+GRtlZHDsswsuukNOl6p24xwrSJR468jXgvGVyTUidxLPlicPN
jNYxUADBEQGuGYpd4lmsjEnf5s8eBHMWR+jBKWpbQQsY3cW1FTs33dc0rv8zsv7j
SUsAGEFq5oufscqbz6kltI3M/lcXyX/3Yw3eWOUS+RnGV3UV9jrSmWOXLBR4Qiza
+FULgEwwSAuLUJqSg/u9TRvhemkpF3jBuq4dxT6Fki/FrJO7lHXcAks2oSAh5WJe
K5xi9+msjTiIsTxJDczS234hBKGVBfvGOc0Xg0rEyzAg/8uBOXLCoVLP7d7mITYX
s6zhBzbgLprSP3S/xLBKxXyi5w+aCuAxHESO3bKB74T2GhT6mWIAEQK/HGCfUOAl
qurVMwt8xdCJScQsJX6rb0uU+9aBFhwevoH7H2RgO+1Y/UTuSEvw3jBffwTL1GW1
cVlvFUMMn1/bBTLro77Abbk5rM5t3c+UAFnVjRpDJW6fY+KU+CFrDemva4Xxd6KZ
0PkT5C8LtROtYn7rMCUTXw1fTIz7wnoaK6iAQ1CO79tmWnyYE5Nq/1Vk84VcAWMi
BYags+Yg0l7GbUBPtg0qmlxWp8wm3L65qHCYFhbDL6D84qudvHrhnUDjqEUMBXzX
JIOp/xW3tjeLJn/Nwi7YKhiyss+B6j/2o64nsinypreWYkswMV0gDdOXkyT9kCAR
k77bIyIsQQal66faw5f3kKitkNN0kdlug1bsC4pvGa9r8Sq5Cxhgzcjxnja/13Hl
a8PRMKYWoZMeynQwHnhScq+nPMZbdSiw5tvVvk02qH4mE+SCHqbt95c1x1Jz2YBs
lKeJMuN9QvH50xezeQm31d402ho2mYUqic0PHQQpTqiJOQbPnBo254xg/NJ5ShzM
F6IJhG8QweatUbBq7OhniBHqdD3WS5NwjGLmH6i+/tNdx+2vFiI85SKkwvWdn7u3
DAqnnXRRWG7SEZ5mK0kbWtOTP8K8xcZLO7ggWar8hh2P4JeWTY2QZmefGEXiMGbK
0k4Qek21/EVOE97ao5PcQDb8IyhDLxCh28O0IVY0KAXcFgQAMxbV9z6htb4vLjV9
kd26ZBfuQt4tIfQsJhZ85jLDW/A7p2vRIXfw/YFKi5apnBmk1bzjr+vgkVfDaLq/
/+o9YKknmniESiW98PQA/6Ji5B1bLPcOYv7TsdLiKfwIbH9uVBNQY7vrXMM7T88n
kcAICoQF/sOGL1xKNEKmwFj3/V6D6Q3kBDxxUQAydLdLJv1ayKBErg/XBWXvvz/z
0kdDsAsicqtn8MOncZMFtZFQVbP6vyQYCAxAGYXvQEpDQu+C3PkLcyjDlBHUpVlD
3SNacUhhjQYGb6D1eR40cjaD+UO31DxB0g4SMKh/JmEkaGPnuN2tgrAkG1xnBJWB
lsq371FdBns0whH9WOhysFQA9953j4jH46kVZ9Cp1D9QL5teKidydp9PralSdmgX
cdkJCC+V+mMrA7KGxJ7RE8ourCdFZid+oc63aX8Yu88XNYO4iteT7evPC3hiijei
I1AJH9mknzjIz1wXlSOSpGzP0QDb0GU3/wXmgUoDcTDwiaWWyVC7L+G2ccH9u4K2
jKh3jtR2zEhvBChkzn/TwiWZfnsTZSyN6RObtmo4rWpjr2/EH7Ox4n4MmhmNI8ZE
IqiN56gKmavDPBUFI+3P3qmUIrS2GnMz4I1TlvtZdZvaqTb+1+o1YVtXiPkMYEFt
10C68gcI79qDwWCZxcHgQIW0enWHno8J310cDhOrNVr8oeZX/xUTQSfYpw9fbfsh
yABXzO113y1pSS+Z9V/2pou8hWEl5gQ0L/jV/7zyJ8OqkzznHHxRPMZ2bsAFY81B
lY0DDFgPvHQoxng63WLeM5ROxHO3HUA5tCkJrjUkW6qhezztYYTM85HbVwPPUN3W
o21t357wfgNibJU+nA3Y62rv90FQjDVmoRxVNihNwYPwvsVq3XcJcbNIkq1Xlmok
tBNpJCucVBHRNWfX4HSxgSsOthta7dDabOnWWz/Jlzb1wEQxXx17h0z3QDVXOPDL
akWGjeA4ENMws9VdOEzRlF9En4FO+PEIsFk6PVYsVlf7eqTCkLvkvcaqwtS9pPft
3t77OPgDaQz7Wtkkb/iPNU8POY25oEh2YxtA+CyYkf2uULXENefxh0PYcZ2M1ah7
RABX6jcYXtMCjKFhujukq7Mi6PO+H9GmvDWYwHRXC5+S6GFsbeI/UHCAPYhGJc3W
M56cKEmK0jyCYSOxZyVAHK/0BSTN6ygioiWciWXfz6S9nDe7InoD8ZrYt9uWreYY
VlTo27Zwfo0a1DqTvkMZ1PEKxJaBdBrkifiOepYvZqJhl8P49XUq2RDwjMSBA++7
wh7vTQ4WnVObKSncACs1kzwMmVWGYqw7nnl7dqnuPl53eE5EDzSDaovqD/jBwqog
yTBEoQYaFXYTLu/7CyReSULMxyUGGSc2jKXiV7xaAoCn57kOg3Wb28BmV2Bjeglt
7CgEF4ITHCc045LET7NyeQbN1z1AgtBeIYFESWE7MRmyOtEu1rop79jGCAjCUIWP
ulnlUKMXA67jAf1xqwWuXeAqSWuPeNKno6eJbxc8Wum98zdsxS7X9lkjbqMSVTsz
n6HlZt4JSIWzQ7Ly9j7PSaFuUmcLdMUAACeFqMdyU+63SbDbT2n+otk54qsPOVB0
tuO5JmSjV9R2NKMFwyGGbvsxgomnwNMTdSpd0qGjS2LW+4YjkLpZuLoV559OhgsG
tju8fmjcbHOtzYHhqvokhCA4mQctnzqVZkNKwpO8C4sfkHdpaNs+NZ/jWqErAlM2
irG4W0mc2Jg8LZxRFtr12Pwx/WbeVQsC0ChSJkmPtjtk3s+HVfXCQMaxVm4FzuAK
VLDQEMG7YKRH9fusW0MuCTz3rLl7pMaf3zBsEpqcAEeNyAW63HuyNsx6MiR8ftQc
qzIV0SKd9SJq+TXGrkhkKNmFSvXb3E1+Wydsrdhm+rKFUPHOet1Qtf/YWIKi/EgW
dqMjSFmYCBVB0ad9UhI98q3mgImea5NIFyUxGBbLLdowXnBrtaQvhXvINJlfITpm
qb/4MIN6g/EiP2UAExlnkz/Nf6yzAOWp4fEST5Eg72lr3nDMgoz8qLCCQ9dpT4ij
u4lqhcgviOExcMOzt18Dz3ZIPIPP/HdzT80ge0sshigXTM86FSah58O1GOGtRNr7
a6TokRCSFgjp4ADqW3GkN5d055YGfvjxMWZJCyZG/3zYxY0cYmpPKVAb6oJ2eZKx
337HQW8bBgF1jgwjO2z+Lbiy4lkm1tc7Ramz22hjJDkFs7I4iSoX3neCV3tTYrOA
tUl9O1CGK1XQ+xrHpt6kkn0SlOEw68ZPSTmXChtdJm899VVq+ettcpUEuch5kxQP
Eo+Nny+f9Wfi1CgI+mF5FMVM58c31I0dpiSPhD4i16IGrS8jHquPKdkpook8EUmQ
CMGzr8+o4nr2iUYOS4dHrpKarOx/sZz8o5oNomFxO5PYltJJBeu5n9VNovuxlB5h
zAP+hA/DkuqXG43Q6M4tRTjDW9DMLt2LDN4yas9bIbdanTd2LURh1i7nH+HrNBlh
uTkUrNdHHapg0uMMCx4RT+DnXCtGRsJJ8an5xgirnia1ZdK4LAAdv34NOjhQXmPA
JuDn8A2pJ3s6EDMgFgioxnlMKCa/5SXzC47cvkEuOj8BNhhJr1gqv2TH1aWE+ur3
7+zPhruZJ2ZG5LUyYXIRZX8HpVvqcYGMila1ouyTBUkcDEWrTNgMQerOD9It1mwq
QEMnnXlzeigdM+BrC4hOW8S/Vvb55uuHttvQzLG8D+4k20NPzxDrohwh9JkTtFRP
Hp+p3IgUP9kUDK1sILhYsMntN3tj42qFzXexi8F7zaOh2aXHq37GsCbnJSZ07AED
2tstGTqgniyWFIuzY89xLIECmyiUSz5O0csq60UDS4By+v/z1lQk0JlOpabODKAB
9uTNlUYr4cpMKONQ/FhglZuTTlCZdaWWZ9J48rFuQmcEygL7G5EsPlDZ12e+RR3/
KLZNIywaXitnnRYYFfFwXZUK3MaAxWmVZg7z7xFCEQKSjTx2Nxtq3Uial0/Mz9dP
FuZ/xo7kLDG/A4jb0FTbve56IC05z6jQW+Iy1naW+wlKnD7uSRUt0mNHO79Qdzj5
XnMay88EAVe7klHkqmGRCRv8vQafr7gWqvgfJm8amv/VVpgWOBCs3w8xzsHtHpAX
mh490Sm5JdESILi/kTmPlIEMxJIxjENVjoJiPbsIFfS1jyubEZJTMI7IqHyHxKZD
p7fnTpbZRZNViI+i6vpJB6fkz7MDlEz9o23s8BH5pM86ro3NIfs9NzuJGyyVMWWa
B+a+7Izh/lHq+bXiaxr17ku2XSBIRbb7WB0jxuHYRVkxp9+ntPwj67nLbKb2+1z7
15XstfdyBbBp51ixxup7Q/GnLE7oxImYZJagU6xqz9rViy2Q12PFkE6DBDmpkTCN
x1RFavpYg9JIjz/kRT6MNs34RUp1QKKm4U6dJkCdNaWAVers2MM5e1C/csg4VKo9
6cSN+NNJJKd+l7C7tjt+CnD1M5NHzXBYNyvmADlVBbT/P+Ioiy+G6KHDbYkvlraO
RWAezOcDQ5N3GuwHHvkGdfGRrTWI3ns/9AOPvWDLQyHWut7/733Zk8WSN9qAp8b1
8UrSJndbpLlivs89xIuisNfSogmCTtwYpHDGfJTLqiwmh6zKAiByE2GWU3L4EXXj
EdAo5wnj3bbxAmJuQqRTM+Svlvo7vj8Gv0bvzlbpo/oCKislXAjgYTUhNLph6ude
wgaQOMu0WsdnL0yVR/nNHjDVx4zN4Gqn/3nWxQ+EG51BlTndxqIt2IClKLS86FT1
2RQk2VoM9d3BEmr5a0MWKh8dHRu+5G93x2M+jQniJSaiZKdEuUbASGWC2QXRFckF
IqGFA3ncx83C4yMgE2xZFJrcaU8d6o56lCFI8F2rL+kP6qKiQQ5iijqo0hBrn5w/
zD2fNu/0t2rYDGaMfChJ5cdJ05nAVvm2JjUttqwwhpo1x9lMWmp9teR9H7YIwBk7
GV/fJZBQCGp1jVBZkv8co9dXt3SPuWOJFWi59d6I/atHbEmFQP0lojv3aXwUDAD/
gWJbQlzYh2lc5IeCp2FXJsYrULEBSf8OvUrw5cCdk+VT7OCC7RJKc/2iXvgBpbBb
RvjChkd35dANEOGKsbp9i0ZcnMmgiTX2QrYIwvxr9MSCClMskCNbyyuYpFJb+puO
ZcgTHnIiWCHqtbMWQz5a/palVPwv9ZQV3NbLBOQhpE4txlKVqwZ0n+4XqFJD/0hU
o0GD6vfrfqcxjAB5pU6n71/2cipa38RWK2HQBJhZdkGyWALuHJLlCfpZ6afD/AvE
zZJ8Du/fuvko92jhp03uCelH/wE8yYUTimj82TwnXSlmMbqF9HSn3gyCK7HlP7jj
xvtwQRSxJGZRiLtLtot3P1W2Y3kb3z+XYeMlsthY3nwkvrETDQ2mgWbQ+5jnvNgb
Y6mkSQ84GhCxRISrNsxBQLa9PgTNgjPF1v4fq47hiCI9zpxZc72AD/VrZA54PQlM
kn+Gfj529fDhBoZlMo7I18TzBXwc4c4OsnDjGh9ObNgqsP4tlV5yEdNmniCsQeSe
wEP/weLOsF7F9n/qlozYJmInoAr8wMoFm6d+V01bbhyeCslxChsPKEzKGIYT/8e1
qcW7EgaUHl2jqJ7lqvu5Jkqm/5G3E/h+5DAYe7dXfqnn3YMgmUgL0FqrhQt2uuDD
Mj+IBQDpTgR7Ku4+3sHZtBCDRgV2bU68/y2QVSlOhteCtUGKCMEcb9ehw/9Q1qQ/
IGmncYEeB4SuYg7kXtmutX/Y+zSHGY5iMvVaCQzNfShusLdhssqADiPFMw496o6M
9th1ZOV2pAKEbYNqecQfTD9AGhVTyDgJQE6cz4+UeCpC34ZflklgcSw9O3hZyxu1
MunjriBTtgYxrAs2jacklVNjQMR0+NdHtdx6bAQJ4xE+wPWFETn8xRzitU14tQOE
eKCD10RNeKMNvR1LjDj2enyDeF6IOpJneWFzIXA6hqh7dkyAqlYMEpN4D9ylPGWi
jTTbq81kciaWvJFi3hT8anlrtjXPKCsui1hijtZ8JQrAxVmHeu27+LCPbEhm3B7H
PwBWvuCYDBJmCFww+1CsukJm4nPptT+cIdLT9GjZkwVYBvjKIRXMIqOaqhwyU4T9
Xmdy1DKklqWJBLn2PPfckJlkw6nwmxieA2Vmg8moDBkZzWycz81Osf73c8Hp8iWL
29SL93UXOROTApFqAf7YN4YduOhotDwnv/OUDNIC/BtojyFkecbZi6rUDy6YxQx9
pB+K/NLG7CakcMsvS+L7SQ7bsPVN1Z65rIBzZGbgH7mUretdhjxBAo/9nAf+92Wr
dNhiU13XZP0+K3l3ppnM+UmZT3fCMB8JB33F9ynKcuAvtQ5/bI3faVsX0+LVeNhn
qnmJH7jaROxW7YH0YWSKPxJPuWCz//8p0Svz9MjuBF06ec0TCAU9G/n/OjpSkWqN
38yu1Auk69/2tplWL/0j3lQMarSYW1yL1eLo6YYN5Gjau3EH9Tltd9g3VkdS7BKB
36N8Grij0ZC6AG7Fx3wpfxRGZFXqxJ3mIrqCl3r9SIS20wM3pHDlnrOqTicz3IhP
VQzEZ+gOtki5GMbi0kn6nvIO2ZS9H4B37Id60np9339HMHVT+kdqBc8cJR+Goo8n
n7cZYEgfuzufxda04r67D94z5B/i5RUl7ni/MtPC9OxXHJlcD1sryeMquhqJpGba
jiu4Kvxd1UuefNGRI1xDMZtn39C+ATjG5+g4Mp7CWb+bK8N+rx2/vobHdDQuK1KO
MxmsaMwe3wdUtUWcr3CBg7zoDxmD39JnUf8aXwTUDwnLGXdxv5GYR1DWut+mYlgx
w5eJMeBWVVMeZAdburNMfGrbgPt4V9X6qUpVh5VrKsa6jsiv0fSvtkLM2nDuN0Wk
aR4LVTiAumQlaNVXT/6BogiwAk2mRElvcKGfGDudr367oS+AII95iA5F9tJDgI6/
4SX0iXsUZJyTq1Y5AHnqDzX9VCepk9Qic8UcQG02wzJMIgSwhLZ8FM7t5sLbqFX2
ivtU5Hht5bLe8i5qbV/jLPhKWSLwnmwh2eC8EYZIA8qKme7k/fPF+hm35sWuDaxj
jF9HHGeDrAdsojileEanVUDEnzNKapWpsEDGyUmfBhydAuBT2Uu8NqWTnD8aiEIw
M321bRtbULRwSIeDEynWyfTm0t3n3DpAW6vleDtZ9GvAViticz5iZExwnt6ClYZ6
UK6XoERaGCF+oGTAb+nrx/QrWEdRCi/KxcDAU+acjd30umQ1uvVDiEafFBNyVUj9
zYRx18PFnJ6S9rIy+XG61bpVH7JxkuuK5D/B1ls6Iu4ZlATXq2dGRKFG/z8H4CAz
Q+RZO0tjEmoFy07XI6rSoHqZeH+UERurWIxIliwdibVo3HH3Od1mYc6HdakN76Oj
plvvjE90pY47OHyuttfhyg8RgZGnpZD73Ehk+lGfmi8CZ6ZBdNNMVRvzREy82hI7
k/G1X7Pus59fyYN9/qTXybnuUd0asPE/JzFUclK91ZhRiVJwpbEg4tVfxtpGqmTa
p4ndtPx4jgDOcssXfl+7NCWNoS+hg5SUH52qj9+OrDCY9NBU44nKbVkla5UjjQu1
qGEIFxKzn8rcnXK0sBxGBdygbjcTuAo12eY+wWUdhLvHTAoJr7u/1HzFNpV6K2RU
fS89ekDsPa1YBcSQ7m20SZOasvbV+tnkRAJgSiwM+2/A6YUxb8bzOz2Vl/qUNVZ0
RuBOgpIaamru70slV8nkRxwHDGzPKkwb/44BpFGc6Ihg5r5sjxAs/HLhrTJILu2w
wZEvBhgghMwXUw3zLp+HaZxXhXxeFeGFasF6i6FKr3CfcmFUN83nk3ce8X5QwXM6
a5H/GZYXNy9WcM8eFdC84IVy6KaTzEov0LmpDPxVsi5bbFvwD4CcW0Q2eZzT9+48
m/AoroSVCIf/OtaRO7JDq3zhQKcqW4rIC2gXl2zpiYGell/YK3dDkP8EnsbKtDP5
ofEp0eXkGIY5WuvoxfKtFM6xNEPJlVfnuKDlGjPg7iKqpM32KTvHtftLyRaKH+du
SJcReIkK+kMabLkHNBwDlCGinLiEiz8DX5i37OowIpefOLWo122O6IG9JSH5k1KI
XrwV6EHX+PNWvVZFFRN5Hp0EbR4BiGzNi/QXsKAHO824F1qBEpIf66HNqDYGCtM/
VKwxfvgBlsFECOeA7MjXtR3Hqm0rK2aRmpJfC6eAzmnY6Yl0bua/G1tOiBPach7Z
hiA3O1KHXgQTDBcItaBp3PEAvao6Xf/js2fVSeMQtbmnRKsaVKDcvxKbyFu/7I7W
ChmySZYXjhylXJtcHASkCrta7yUBZJ94grTHsmWHmwEtkHoxmeaAjebbo4ADs1Iv
7ewpsQroazzgwqMj/0gIB4vgO3AHv70SKnlFAoObo14vi3lEkzbYXogCMZ2leCDR
nQLAQTeOPSN/YgIRE+3rqupNlATtEXhqDpUif2PprsET3Myrs8jA4pT2jHQIGhKI
bBNt9KFb5uqUfQikHKQeYN7pz3avbTAAdy5Q4aoy2Ft6R1N0rf6EQB/TWAhiADfx
anvvdPxCa2iUkN4msVo1QyogGjLhJX3jPiKagpP9sFH19pxKC783U67t7ayrB8qs
ojGXDADtaYYjjGpw5J11cvEkrdJ71W5eX/+WLkLBea4+SbGyyPHHeF5tWPsUhWen
gYDsaOHxEFuZIdhtQYNgFFHiSdW1jqzJZEJZPEst0tMwjsWNAL3KRopSZe1hAq1B
ThzcbMZLzSXSbiZ+vOcSedmtYxgF2uiF7uvRVVf2eY/8Iy2aFliVz9cxm+dtw9HA
9Sd5o6Ld+ikwAj3jogtSGnMsmEuSForjzxtHMkRe8RWoOIRdg5fpo19vzWsZJw73
BMYvLwHWzpv4wQEZgqyIxE4ZDcklcGnqfEieeGXUSsEFgfe8ypGI/Kl/HXSOz09L
aBN3gdzgWBR2i6OW7ZGc0jp4Zat4V3FZ1Bqo+rjAe21xWbf8xyc+ZnpCkcHlfxph
ydtsydqRndJNmLjCeG36sX0+9OrEQorEyyW4VClxiNlr7w/tEtQ7g14377MqPo5z
D4h/7O5jaFBTa3SITmQHZd06slV6laULgHaAm0hvko7zwCw3xeeb+1z8PmSSUuix
TmKPu4DledB3xpJAFH3dv8xGXXvUN8CHcG0Dg5B7rn+oZGhIX2NfOO8k8A5618XB
w5h2eL+4yTx1qtbh05azsQLIitryFozlyRtFs3NrV/9q39DL37+MJ9b1MNchXcNI
EaCIMcg1nC/bKzA2oBro7XioLQhoRFRPmA+TVDA8k5kfRhyxJx6m3ys2sLPHAn7Q
XWcEuwKwAr0A0YWUGB+/BqYJwwCVFcoYS3yT6NSbLZKBrckHexqc47aoBpd4towj
ai/6sxOt8ZFZJ+cjQ+hwEAHK5AwHLsjhxOtm53mOHXOfo9lsiwkmxxr2bJFUg9gP
O2ybFdIXUGANevnna90xTEmLCPZv3qBgSKMj/WtKZiY0JaK1EF4QiCnG3ejEB89W
5ITfND28QcN8GLm0QLM5XJAgeb7QJF0Cjp1knOaXpKDVaRsh4wi6G7/0Ge9bFhS1
ErEbCPEVrfwK+npdX7NyxGMZEvBCrmIzPmWzmXxsU1zu4U18L2F4L/xE6AljPUNT
SkMOAOof4YRsoaXx7JulaKmDyNbk29XYrMAjeuFW76D4Tl4Ja6yJMGfkc/vvglCZ
cSXheX8Xryjl42X8jP68GgHVg2pZczpNjqeeh8/Kum2ibLJcWoSqLvBOrl1N9IrU
wRLMfLv+22KO5gIJUM3N/O9uGIkweCCj7wOYgVNHAMrs2PaE0jEFddFgP3Ulqt80
6SJM3wygPN99cdzuao24TuRruV24TaxPeDNlyhw1m+DV9GXIKMuxvP2u+ruhGG9v
50YTD9BCb8wc7e/y9ICpGeHhw7PTBa8yb35KDixQwOBOgirA1Trd7CzFPQKktLNI
wyUoLwFgoMtEtFBQI6ZWMpl0rCazmmXstejfSh13Gxl9kr0Elaz16rYpGFNiBZut
D54ArzOToJqyzN6TTz+xdLNqAzWMU4GcrcLNR4Oo2ipDS1hVM87Mbbgl7C4JzUhT
5rAQ0pw74d2r5U8uhzkX+lnXbUxes9niaxUhaHCAQpulg/Pq/YJeqpebidwm/duf
qdZcZAh90XCQ8gOIJjTo+DDh43zT+IKQXyVYyKIxlGkkDBIgRZx3T21TftNp5vNl
F+pCjb9ql1ocLsOs63d0o22ROVYRNEmQYwLT00P+SC3Fw6LofT3D5AHHKewguIXf
MigkmEeuhC7gZtvCP4wdJ+3zxdp334QmEb5q8aV8Nbt+So0DlkNLjjtN4YbdgZLx
VynqhLdDv68ylzTNfCFwjkSMBSl3l7fVzVzhcS4pTJsf9h0wggJUNGUT4o4c8+L6
pLFfqkDon9UBxBf+5axTjCV0kH18Myj4KFefG+K+bIRCa47hHI8rVD3KPA6sxfDf
gBcKrqg8UZHRxk6o4AsBsXBeRW5+m/t+PVY88J1eh+XVaCQ3OjXAZrdzKbXcs3AW
qmbsrN5FardNi+gys6a59HLkpZDDKuiSvGpMSIvMrPpctZTvUijgGtjpeLwsHlQI
0rPVba+7/UFpIr7MpDp/8DzW8iAfUlGGr5BQE+RvSva0pVFpha/YwoukMeftPzJ3
UcVaVMDdtbFu3ikMVDfSgGvUADjM4EMdDPvEyiHbHIlX1/qLjqe+rv4Zx7IAFpv1
xSbUv3g8+hbX0fsg2HvxveIBN+m/TbF1+npRVgqPAHlTXpsnMo30/+V+Z/xLz4tI
oLN7El+/zbIKtnEVT0BAGFXZbzzrbgSSspuegoTyVcsShuIZVIpAeAxXq2fPLTkl
MZfzs/8XGYq6AzhX41zeNPlH142j7P8St5+Xs811riNSVGbtcz6cbEkF1/ovh6w6
ttB2AT17B3oWchqMQ9e5fkf2NsBf1tNJjCzC0+sR7bA7bbqJjM/CkvBcrUaIbS1/
C9r+knbenQ5LJY0kqIxq8lk14mMYTDhYvHnfylrDouCAXXpXyqvT2LeqKd0Wl8Pg
xsC7823gCGKeukKoHtSZA8YuKyMxIhqjDXpacdOFaIsIr0bfFI8WM8OPHEK5cMOl
zBI7KF+9eESMzQbIHO3AGBs8T3axFKWKYQchekBHmhwXVfd4+IWLbas1VZ1u4bFZ
byZu8CMCo+DUQSbSGcYENiBDy+Zry1H1hh04ZOS0eSiB7M0r2cnfroUf8nLmLGnf
wKr/EM5n/gxOC20CegCVNurq0yGi8JtguGRb/HwmodVMgJrqg0HWk+xhiRZmUddY
LCuMcpEDUvFOhpP5PrBaITM0fmlqWMilE5tilDQqD65AB9GCQV3VVGlrxEhnsH8T
mISeyp0Y4Kr+rAl600HR9ZrnYaj2CaVDrK8iarbxZTHt+Jeo1K9CC5Ejk8Bl9i8g
TTj1vTCmZAeXAAw+xEB7C5XWmit+3cWo/6qixxozP0uW3o5fL4zN5T1snlv/cG8W
i5PmtVi9cSEJjYNgAboCmTKkLZQ6UqYrUVZ9iyj4ctpew+ybS/I7mKo/PJdzK8jQ
R5QUKPbziV3rddfAGNpGG5NPvA//u/W+BG8CjKSQGQq+c+luisr5QBIR7nroTWiN
cQsrWOVM87+fRy/Yh01QzbI7gvmkQ0WxusYNURucqTeP0GxFD1RdIqiBVn/n7mSR
hrd505AqEjbmiGNKM1bUHakUQdQfSqWrQyiNTvfttJpCfnu5oSxETPBzmtd65h0g
JeADw2Nz+ZGqm3yYzgoWTOV97c26e0gB7xG+kfnueE90EKgwaIKThzEDC+r69CVJ
DMJ7Nnhg/RI8yR8i5+wCpmPAkwqjMaYL/X/I8Yd3IkbdK8PeTga+kXJvdEObVCfP
PQyqOUUFJZGh8xsIe88HbOlTace6NJ6Jwev/vIOtZk6txNSbNTqWdqvQep+S9qQ0
8reHdR2ATDB4fmEjSX+UmxbtTtVbuGt7eyqlUcQNhx/eMtnMqgyqqy6UnqUxR8Lu
if63VuXj5yNrdZyOYsP7WWLWRLYJrhNLoBrWfrhuAovv9Za4wMgj+6hNX63R094P
ToA2bYuBHTFyCSGyLybIP91qiOMcFgR6OwS7/aaFc7T5+OcMZDo79kUjkW8otwI/
qzm5gLV/D8u40/o5jtVG5G9786ULnylC5V6qJOR57Qow6VPsxj23RpPlErmADnRN
ttm5ilUnokx4h6ZRZNGjDiN4/uvuXyyHL8WQIIlS/O8d7TKsN8NKrQts7Hg+s3Km
He/lDlGwd4Ao3ftUL3HrsZYqFuKk2UpObMxShVXd7WZJVHU7fTA7kiOwq4BQZ2md
86dYNjb4OvW48F3tu4sDbOfYs1cHA6Z6dtAmqv+JqSkencC3CieUpqkGI8UPiZ2x
pimDzCrUn2U5sf/vw7CulicW44FFxXj82Cf744NRGfQKJnBbOHJ0oPJo+wEm9Rgz
4iCrO9RlVRHOR7MTKr+EagJiwGmVG5EppddkpPIpe7Stvvsn4PPSfCH25A6NmHPw
+YjPeJ2zbmnUC7ObC+FsUr24Gc1IwpxViQXwVsV2JMMMN4JGOZeD1EGEyFT2zSMX
dS7koUDgVZ2Q3sjk3vfRKx74UUvES1CYQxdy1BVibfMWLFcz6H5aQPnjy9jKtrra
+ziMLR8K3VUlZkoynog5AIdSYcqS7Yk/sC+g/XspCLKlO/sfQrQ/EjOxZNrhos5u
pf0ls8QsEgMafn/IViLFaxBi7nPuil4rJ69FByzH0QJHPgzYiaIetTvO1iUuXlfX
5I+ye5mThIXzWg5wwOCoV03/Of9ZfKVgtOauzDs9SnsyeMAJKVzyxBiRqfWKZzaT
6Ff2TDB/FoWk2xRvkLb4fHSM5zcRDeEJR3goGZj4YTPHsFh7BKpNrnruvIIqgxAw
NQZpMw4OdWMkG9WcMFjIkjrvlM2Pv4ngKlynbNPhH9BCMRzXT0Lm+AsBJNgVPj5U
aAjXYIFI7ZIGhBgUWWAu8gXH/Fwyst1jmHARIDe2INUOwV/MbmG3aXu6WmAHvY5T
pQp6yZqdxRI5LWgyU7jI0qppMmBXefucd3axQ5wWdtmY9IzygQSTZK3WP5mJaS2z
cPsZNToS2NEZ2oOShHt+J8cGAueELxsS383WUVfccFSn9RvZHaCtnDTh5glCrXfC
KkbmzbOYVMVVPpgz1EVUsDKaWYPeDa5r6rm2oTzappurgwhRNgf0AMSqvWKeNfUB
DI0qla33XxXWDoGGQTH0POkHUXToQ8XolNrmW22Owte+tClIOd2Xrm7ncJeDu8rI
XkM6PcY/tPJvFlh3ua4ijaj8gwVB5eyNPFq5AwFJvvrQ4Q2MrePofvS8mjfOxYxU
vqMp3+1jAk8gW/CMq3caG3fmUJJVkfceTTw8Nm3OWZeh1hyIQVaV4aSJdVMwAgiE
5bGc57bak1P+2FtVxltmrWS16eoj2rPuh3Tsru07tjkxC7pB4x4wQ/5OVN7YkS6J
XslN9kKY8OhwbHvSKERnM8xhaMGR08ApwEkhPib5g2cVtWun3XPOdNApRn4KScgU
bMpbZhl53OOSGUQdZgOfKTkSCepRCx4Er064UKPjIweFiOWLbopFc8Z22DdQLFVY
7XTqxuF/mCCV4enY4KKGoweBJvsFl2mNPqAsvJoRX6M0ZNYJp1VvJtPsNR5wSRlh
Dw5oyX+nMAQUE48XL25su3tNz4Fy0alN0QD1RtQNMaYxAfi+3/9WD2Q4WNHyK2Fn
uUXc6t8/xeD0QrafSYl63oR7Zutmt0Zakop8GHyPNanPyzL1HAFMw4VCeO3hZJm1
LiPjzyZTKK8DHAuGi/ECOZsRhTVNJRWP/v8yz2Lg949RWz3lAPmq2KypPEzG82yW
NoRSkRLdwBVYvSg6+usGjzJVz4hfio/IZz8gDFgWVts+UJaDMxkMWyt++WjCkwj+
EG4tZaKRCYjz4gDF2OSJ97nTjcBK1VMMH6kVfo9Cm5UM8AivpPnOfORlE+i6uIE4
OjuvuWX99xj4Thnxq8+WY55KjfGpnToc2O0ppeOXy98I5VJqKxHwOmu4FKUtuG/E
6jRka8tWfOOHh8TdQM+AUUwMhogVWRmXfbqYnZEG1kGP6dCFf//T0nTECQe89LDY
Xn0aZ9k0fq8jem4imEC5mcyhlRVkTwcShZEVRDK/NCbCALvuFNzqaywBHJHFrbM0
44EboCuVOclVib1yhcP6EOvNn6/AhEMCc7l0ZuLkf74PckIJ/ZON126+gfZbwQ35
ktq/rndh4zIF6lf+2cLSxqWNF3B2gTGf42Ksba7fr3tlAahHh6pnqTvvkQTmzeDk
V9aGUsgGoHCOyFct2X+xiO6AVMzWbU/89+QnqtG4d9gR6BH08chbKkzeUDXUTzYa
hHK4zdNBGssBzE1nxB+m29bpJIHR/Pvl3KayIzYZ/0dmKh1Ue/pdpjWZ+qmEYjmo
gaHX84bO5rpkQaTYJFe+NyP1Nu1PEPblD/ijv8DvshqKocByI2NXvezt+OBkHDec
NMFxY4uPbozs2wpt3LEaYSxBl5DeyEERUi1NI1LXTJL2OsVR5ImPbYlwoYyO7/Tj
GYWBIgf047bQgi2gpnMjf6HENNwqJzTKpxCUtDWLWnPPYcmXebKBx1zBPTFT046y
tOvuFZkR9yWXYHIn+gF94yLq5jqVucF3KornmoAhjFcOUjYXOKisKbvjhXrctRvD
UyMoO9ZwpL8lA1J1Rp6mq4LyRBn7MxdcdG8zcgXgc9w0X/QNTynUoyd8STCWlw5P
59tYPIgLXvy8sFpkGMDZIVWkhA51eWM3lEFvbYf2DkpU/gkYLYJL0UXpRUpKXLiI
H2qBUVY+OvXCFGCxW4gwuyw4NLND8W9s2AZkJnwSGZfPuTnW7+qaeoqkP0RN2rxS
YxXFN8YLCI0A5Y2YKyqSxoSEuVXP29fKklFfUD0xM7V39SGTSdbGpRFJ6lqWg+e3
H+YX3Tqe9qi2v2+zJ34P4+EaRudE3uQR2jCTr4X9sD+1x50D09hHCwk/WIadt5co
ipEf2wHj2C63+ew6Z2adbNfABrXXSK2x/QxkdPHGDaU5LVjH5hpYRtKC3uIEGisO
5tx85K+ngbgmqaL9Pz+srI6z7DkEBIhxg/Z2UwWLe81ztg+ELqZDwJJT5mFUkhhe
8UbTtkX5Ptkc+CzZdSMbaMBVL+GynxzDzn9aHAH+Oj7cifo2LdZRrrGoMBFRXCbP
8ui4bRec40oKlIM3SZ8V2tt5pCvAiUTspBhJTQkxwdyjxPzLaUXJz89F36W6gvH1
abkVVCMVYjRbUOu53SXwL1O/l6tOi/1/fZ2WssUUvx/lEXTJixaEfcZW5+u6MUWj
Xcr9mpe7kyCJIuHzHJn3Ooelu8o3CJoLmtysSGzuik46Y8uIUW07s64hxV1FcQe+
ogn6dDOVE8tITy7/1xr4VP7cLlCDDyckQtK5bnI1Px93xG1xovutuHYlTUO/MZfU
Qev0jtNzbmvdTHP5RKeoSCAPUwtRr5WdR1dJIAWgsd7d3t/e+ibs9uO5Y7WuC7Fl
ExtNzn2xSFSdoQQQrXMRj7S+jmq+LyflBw/2UkSJk7zA2QhQjyAGni141dKRbkuz
ueaY+LVB4xEiDij6sn5a702EWki2B0PFxZpca0PUlSdJ7mUbL2IheuNHdGI2YNh8
`pragma protect end_protected
