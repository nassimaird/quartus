// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CwyVR4OGCmzC26b5P5IfERVqut1SToQbVG0KTW2ggbMFn0swEUUYJkabK8jPQm9TAv2G9N6MP9b7
GEVLAcS6Ptp7PSNUmGIx7KANpEjk14bz+YXTNO11xeZ+kQJbnrsTtyNVwx72rzpnfGqKvPsHzz/o
YamKx81czF5TKT2cO3sYx5KnJLnEIRG5yPbonBZtA+OVDcpP0w8qnYPkrVJssqFVDpgTQpxK7xwq
rIqOWB9Lw5PYqF6qO5t2dcnKwHEsTOlwyzmswIuUGmAjBFQzbidJEcBQt9h377cptJlpWiPQ3szo
AnLHE3Nh5X0rIn4co/+H+Uizh8DdUFjyaiQsJA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11456)
OZs2dz0ekP2gksJ0o9u1h+Qf3bypx+I5LFsONcaljNWcf8jA/mo7xni1eTwTbOdz/Ib6ghkrR01x
WW2ZRcEjMKuX1v7Z53xurbjjeN5r02HkKFd41IcElTbVbg+GV08+mya2bPzhWgYMW3JiBU6PAY00
MTRcpjo58791q3c8eTQckChNlaxSzXhN1kC82phKBsguD9gzaMyhjyxXG32TKYzt0ab5l5mRABDc
U6DovS0lIUvk4+6hRy1eynbROVVprLPKdxVZKMZksrB4C8/gorm3+Qn7azK7nkuUSH0UcRJViO0z
BJZc+m1T8UJVykarhhjOYVG+lY8Xe2tNw+5iJofNy9x6RtOtTyoRMPME6HgHfTs7l8iR+oyi6eTe
3NLI4efJxGHrmGsB5BBhPFFaayvBlxqsoMlSdqAXvNsCSJ+d/HgoT98IOO5LoqARvqqlS8OSJhXn
zsl/1Mj0h3eQbexnaSTnTnyXtBI+ebNuoprZ2FN061ypUlZarcDA+C4Rl8ZtULDSXzvDrhngZu0v
lNmg4xw+yS/DOBa5UrM/NOoKKVBQPCiCsO0DkTfy6pbrrSa/H57eOAZMQroA9Fze/9+cFKgwXHoj
aASFbghiPWj56OHuklTQv6HyIAv8tvu6IonXhrj77IbVb45+NAbGnt5MJvSZP3fKfN+bhyS9z9La
JZRPSbCTOgigZYZlWfPl+i/LFs+/JIcFDXbuYwAjLnRbOztkojARRsV2P66myMvdP8DvyHgebGS+
C6vMv5JMaBWIruMkyCSsTMMwJpD/fi4XBV9+tpZlbpY+d1Bhb/lttJX/tKMSBAb2uoo7nZgixy0p
MgP5JTWwzuQf7yfF1Yw4HJuPRcztFm02rxa+i461a2WYIpRIwDHeXL2/pXmR8nicDHQJXWQw+4WX
oP3MOvwSfVorfwGaQJ6yLRlBafUyq3wKiHXAdRk7b0/E4RHNKb6zlS6VH1wfxPyilIj9+r9lFkFe
LkJo0qde+oLjeueueGhnK2aQZi2D9+2g4cbkOtC3hZe0fH+CcqUb+wV934wlKvQp9Ezyzspyd+Ko
aHppu5eNMoXPrnaiMAAlvywL8KqMO3nonUzf9FXTTIrVuo1RJPA+1ych3E2mdpJxctc+ZzCpL+0z
Fn6cJFL9Vc4CUmSwqhNjRr9Y4bq6/nisMn5jRZ+FIbUE3NXDv4voc9/jg0ItPU0DG09F2xm/FTjG
rCRqUZE5cMxyxO9EC42r+Bc1Lo2qtsvRrPj7GRV/4x9mFIIqG3uNIU8kC8m+YTeg5dMpte/6oSU6
TtIwNM7K8V+5qMnV5iLxr3Yj/+kU8MUUhb03QnE+n+sM3MuNZ3eoMAyPJw5Lf4YTPwiDhqg+fcj/
Mm7d/vAf344++AbwQ2ya13GEpkBVwTWR63lL6Yx63AzrDhcw3RrM7ik20WDbKSq8ypX55Fk2OrTe
nZkNaHh+NA12dVGven2MXZGxwMa0GushtF06qfQv1JpNW4xfQl0UliFu8yUTGsD3JIhesgGgIBqL
DnlbrYAfCy6rVAUvFTU500ZKUlhbNC75P3YUNUJUYNYQiK8ZBN49Yx41AZfKIv+La64vy/aMG3QT
zEqxuzB9zzYI9x/Vzz17fH65koBt+NIrSITNqiHjektNTSWMBQn8++TRdStHkfcQoJYQd/7HzaiC
Ky+Nxi2vU6azTO567HBVf+OyMlucI+gLPwMG6lUA6hcKi8yQa61BMXsG6urcNUI8wOkeqK095AAW
GZezFTWVQFuz2zned427epvx4vZQF1alAtN5APvHCNo9cn0oCGypjvHkaD1VzRFwKm/g+ob078KE
ePn58cLF0ZYQxB0xqaqPuuXeRoc/v/Trw3pk2zJ51DAk1AsXB2g4aSxVnnTVYy19mYY0eoqKXK/N
RN0ZznUxY12xNT6rXs57XQPUmctq7q43g0YCS43qPUG91xRkcrgM6xeINJ/kZm9RwuCU+yrf1/uR
d2ZxcxxslLWBsEZh/XRdeXN0EOV0MS6ZyHBxFSi5uoPm9z4lRLtg4vbOWjaPw0toPQbnzHsIRkXB
4glGUtULH4BV2ClrHSLJcDWMWneczllizh1ISAZpJ+HJl3iAE0+3N9pfhBvBS4nfvpiBUNxAlAXk
mlQVC+buoSYO0WscYpldUWGIyFAsRywNQM1ag4ZSprpGH9Kj6o7oV9lWlRbRVAAQYwi0KzP320Zo
yfj4QTr8ugX3yT/TJE7CdEr6TBtEt5qpubl5Gu4PGccDVflT4Qt/M0fW0e1KcEtr3OA2OLn1su+9
VQTTybDJcB8byFNDeyOH6xaHYqR26vHZpoJFHqOa3hkfr5igmJbQ3Zcz8HP546zrobRJnFXKEzRD
zEWzmXCHPMhug2KJd+PEHnrQt3csTVDp1n7oymrwHymGrwM/rGrNm2JvOieD8jEuhSIiqDXEGb0b
FmFJew+hCFYfGCIcoWqP9lrsdyvGNseXLnNERlMG1ZNk+7ly+EKCC/9TWEDn/TC7goc7RZlVC8mo
9e9by4rUNPj1SJ+XfGfOOkaVOtCiCS0GxdMHHwqwBV/MmGBT/U3JwRgyVxyaINzbRCsmWNgCXphC
i/Y5sDNiqrbSKlMk6cXFK7JDHtUP4LjPrML/5KwfEseainfyXTb7kWxa3OrDHY9ti7NLEIx+2RjZ
5I1zQrIknzGGXtXz/UQOmuYt1P7dvzq3qIl5W2YE4nI3DJVrmfbJs8ea+uNLulfFXrKXIlqMqKAi
MObvxqLSPsYVHFFTWSn25ymMWgJtF8VYr2uw0mdaUeSzNf0ND9W2rsQmBfKGQI0VKFP7/XdmWODA
i7jsEr0z4g3Q6vPyJmnL2H/d5cEDr+3jpDOtra9WL86ZKmImjNLYtTXrsMqAGaPOr4MlONIljHXF
E7plp0ytf+sf2SISSMU/cJoHCqan2zPHTma0tZYXSjCLTT1+oFE8kqON/wLoZAGE1d+MB9hw+CPu
x5dPmD3VaS2pvzZtM2PlhbviYELMjX1+Wopu54H17Z/jHBvPZ80ZuAnZGu8ah8SExpaZnSlsJLiy
qIg1bOgoKp9kNhnFRHIPnH1D3eSUqBy6xZMFsal8zWVe7ojluVJugpAWO6D0bu9aFuC2hZ1EfWQ1
uRIx6Egwssfcsvj037yF75EKg23lhQB7hDRj7ZD+4XLn4/pRpnlxxkzEfgDAbAxRwsDz2nJSZVyt
o1vdiXWIq8rXrT/dyV2shfvx7XCf+LyNmv8MHIJ342dW0HMrTZGslx41pbhhDDB2zzvimpgbteyX
PmT0UhrvzRsGOcJ5RSr6+dgVtl8+Ru7AKnDn8MRTGeqBuaX6aTILk4sLzoeg553g5QN1faXZFdSW
vUkfhW9npGxEh2VynfZ82G64ur7VFa0z9T9b/dWOfd9ToReU32DXN1mb+e7hzXnYZC3bDcE24TtR
5nbJ0ru1DQOG4wei02fLPT+Rccb29cUKiCR96VKGos/8nQ4jO6vghDk1L3o+2ovEdv/Sjd/4HQsM
euNXoEnGCoiOx3yzH9JOIOn22wU755ddgpkJMq7Pov3y4aTaZisIiVhO4WYCg8BxByJ9K+fT1+SD
ChoFL3GgdtQNqTeJLPM2QEGDBU44wz2M9iHgA6YqQGhUtHeGfMihc+q+TJDA9Mwfz4KYtyXLJdla
uYvYb1Bxio6kBwKXxICrHooHPMYyq0o3hCtl3GpQVel/rxI3GE3mKxbh2VUfn53iOROAmbXsr3A8
bZDytZkJ1RRr1Mgbn0pqTcAa673u140gwYTfBMH+BMhP/Iedp4aMSslFvaBxeGahylAzmkDRNp66
b9ziTdCuj6fX5s18xvAXoygx5k/gXYLgmcTguoj/ZLK7y5N3zLqOYQ/C1Ug2U6IliU3SCEpfaLVK
TVvodhIc7/ezCG1rCqrWZQu3J1qBDyVX0Yti+sZA0D4ZFeM+0fNHImrii0hZkvk5T2V7OoDtkdFY
G/cxp5sKZpZ7wgXltIpcmu+jtk1127Y3mlhSnJF9VbdPQ7vC5HNS/yqtiz/Hxe7afoS0qTM9J8XB
UwV/tfljv/16GNEznNqvFQxghIBgWwJisdLR+fa3P7A8doaDrjBRJr5PUBhijRg2PvQpDv2V8Mzz
PHAtCKL15OpPFvo9/k6iWpoRqlO/fCuhS36nrWp2knoUOCNIb/GP1pAN3PbAxfz67Qz541HAzTmr
+N/wzouIIQBi0TK2lTVzxe2fxLMeh9Sz/KbL2tIi4ZLBJTWvcOYCWepJkwUwFSP8jKbjicjbuEyq
iHq1D7bZgmd3RYASSe3L/VIJ6xSiGXNcg1djiAoQ7SovgzeCRI0sv5QfN+S4pPRzEJPljH7I2mFE
aMeLEV6QjN3nIvWG+ZB2g7PpwdGZMvRrF41iw5bU4foY1t9Ih5gbQDnfrhNFXl+2smnHR7OAulYS
6GL6nxznNfRFAUNwzuWWUYVr6VOmr11yVShtOFhy/YZde4izw/4uC22gochziDJByhN7y41lL6xO
O1GLKz4bXptCXLAS6Ul1O5oq8BVQUvLoM2Kxi6wt8EdilN/FpwTBG8yp0W+JtIdR6VcWFZg2Abq2
dOkxBfHRfZEtUYzDgWQPrmd10HsjyBeDIV+sYYA3xaieRZWTO2wn3PmmnKioI1exL8bzpDVKXJvZ
rQPNCGuSLVs1mwNdL85URPHZiD5GblbB/Vh9xJ6dj+5KN386Z7bvwezIeqHjMPNrppXF9xCb54mX
0ripExDAOfLGYMtgRz/zpjaExCSN3lEXj/Z2uP+bE4xH+1O9tvlYPvgQhfDp1FQ3TTje6xWXbcwY
VOi0AgtyH8+DGmBSiNv/zjpVjWiV/zP12GTidGuSgIXyHn1hRhUGMeXmT54Ez2FyBtXV+uNa6laV
UQnrmlEmEkG/f4ChCJi6yHwPRuOOBHa3l0h9FtxY9uT4DKxraOuX0Xtn0/t3rg9fb8GALlElguea
DX4VXdqnXQpanN3tUJnA7Wtv20O1vIrKSDB33f97mS9oXkdoiHOs8zmBcl4+W7Etf8QO5cypAo32
iriWQw0QT2QAkx4p+DTkDYQV9+gUvidyLu9U9eAOMkDL4bC4nopTpzHvicztxIHg1C8vt0+vnHHv
WU0XT966X1M0Y2616aWfFOEi5BeTCG9ksH3q66WzR942F20NWCzZWpQa6+t2MTyjaQepS3SzExTF
QgIxXpcXyGWhUo31PHP/GBMGLCAPd/1V9aTHVL++aGbjSyNAWgNewrcAD5Jm59NlRWYIbh7Od0u/
W1j+3S+4OIIEm0F1m9x/i2zwudOf7iuYMG1IGQOisBBeeqe7BxsxNn9nHuoE4At3VGi1fouIPY8m
q5rrJ+hTVO9ASZ7Ch4uFf6dVUfN6GIzoaRaYvHrYbCGVrGQz7JcZSXdEpr6VafCkbDPNlIUPmMWb
KjkdeCJCgzxLaKR8mKH/vqMZoASU6ssW+nAVEyixVRsf5IGYDSy63i436L0Yw2GYnNTGN/kR0Hwx
9kl93xoQZFpSwjmPo/0c8gGC0gXu7/C7bljhUXjXu4NR6CNfXqfkGmzQ1IwSWdzdcgYkMx0bl20R
E19yrwtNdg98AyPtsc008AerhvpOtocWFWnkLnmyTKXw9OpuVe0EyCRLvFwsaNXdtJ4cEO0UgwyU
CIw16875f2KEx1dajQo4nQvqRZlsdkZYlCt3oATEQgz1+RvZAVMmOXDL/38eEfqn9wLH6aVPO+2p
uUCejZe72n8JlKukVzEqIupP7zai2l/6m7gkJ7CsFxVY7vqNmWvSiMF7um/AGoGEZSakS2VcYroi
KuQUiGuoyR1GhYf8XG5cca8+wvGpTHdJkbRy4xqoScVc2xNLnrS6URmxGHZbiltRvdOBX1wZfTrT
z4Hw7Fg/qlNTAH/KJIwqu5u1UQuACevy+zQue7Zi+cVSwNlmpj/Vy5JzI0ENUZvDSFbVTJ024cgX
p+K3cwQ1O3O0HhN1S0QPJ8NSkdLXr/8q82IHUPx1Onj/urNh4ezhLWq4Cb3jMZA904FjS9IlN2jE
H0rcgeKOhMjc7QeK8+D0rinU0IDUzYIMC85EPsAZf6TiyWnSFfnAFRBq60cBaCcoXBOvtLDD6jNU
U2Zv5OU7r8lcuG54VULHvyLOtL/TaRYSVEYVnsy5xP3DwB3Yz6Vm/7OuDEVLp2WMIXoOJZ+2S5h4
dqNnd3ka8E0Q0/Wr1FuGt+rgIItzLNYcWDaR/ADtCx3I4m421M59tdV2jAYVrDc9L+wjE8p9J+tf
LZ6TqvOUCsT+dXGY2fyCtlHjt6L/tQ0LonKf9MQQw6M23TEI5E4Ry9O01vwFOXB47Q/sQ3JUDr+2
QN2H2nIxFEKabqj5r810ajUrzfD1XKWrk1sbXEoIuoXWTtMpw61ToSdvcUZ/scQTmEDjuLQMxksh
dW7n/2Uf0C08OXRAlQvdXToiiX9BKulZuMJolZev4+zUYsiRIMQHZUsydlChsFoYnxGgIbL3pkj/
38852AqNLS6OTX3jV7XBhuLfBx+9Dz6Ow8sBVwB5o7m3FZ+LPZrBeeZGkzmEV8kWUA+skexoE2Z+
IcjltYHPwNhgnV5MqlOhFO1OglKH0uxi9611F9zC+jEv9mo13crccp+V/CgtBwLPbtne3IkxRSvi
5Z0HWQ1Xs+aMNddZ61YwxIPuLoeKDwQcLAh3Azy6sa0ddObEXCe0pdTZcg6S7JQabNHYf9e70jPz
plxgqx6+yUOkzEQbSR4M4EbmnEW5E3qA4P8BOxMnROnV9NK7+P6OCk/3o2wHI5SSX0o9D/D768L9
pWtMs2yUmIefkEcFcax7X2A6ZjS9cvhfl3ZthVFwUR3bx7fveH7w9eOgv9ZPMRMlfgu9CWDjEah8
9aeY14nSQ0psmK1yybiKanU8aS3KFMSfNMIowQIZZX0com/g0FeJvNfcFPcjLXugbQZ7SfrIiJvl
OBGsOtHYI9lPAROU2qj3wzffg4IPUUrVmvB+YNAktVFAwbUSkW4Ykreo4IrD3fJMqqoyD1viC233
2ZqJI1YnahZ5KG3CRMVPyXvq+yhTpyQjiTCX9JumMVKMwim77fOOALNS+gbgAW2sZWFgsO2GnnI2
fMv95IE4CiMuJuI5rZVXC5G2luS2wxiSl6xuEUHpvW5AhNMEmfKEJ5EAnrNFzjF2u81ea/4/lCQe
AvUjb2APWyZs/2/KiOTT8MxutmSPHhupXTiRMSp5jI/RTEsG+FqNfedFqjnUENbbrrGgqGFdhRD6
coqdSxzHjSa5kXOzbZBT8mbux8PQku7mN9kQ4pBka/7ReoQWMOnTJ5SVtQ4BpxrdgBn713XPVIof
LEPClaeFy8ScYiIo3Jqm/GbBYUK5uQDe8X+5ZMD8UQLXdTUcUgbSj5MEuv+KAf4/6UMJ2DRhmgJc
hc81nC5O1LtVLdM+p2Q/INwHzFdXcxd2W1Bn70Jxli0v1wCtt8iDf1FICJwxPPHdbz0ba2KSQq5K
pvFtnFcUrd4xcRkrRfAaq+D2idvDy0JFfAguy4xxNcI5ER8KQ2U/IkoZuF7RScJIKOmayPeIg8An
OHSiJdofT6fPhXV4SGS32pxCm/qFsam2aEZ33c5zYzqj4q/IHvLSk5LPTvEJpTxH+BIK1/GBM78F
CFu8qAqwvF44xZdTr/M5r/l7vtQKVPqqjB5trsTJpveY1i89f0+vuZwapLvyrNB3B2WN33+ObGNU
cli/vuZe4S7xwE2LcYL9/pGCALJw3Q/Ql8IgXh7tqhq9aeLF4Nri9zpfG8I9YdZO+/IVe0hOrNab
zaQhI9oAvr2mEmSRWCAwF1ghPa8oDzym7v+BzJsOLSlKjboTOF/Q2d94DcST6E0i6KjYDSu7XqBw
IUFLLvcvMLKAylpp9HKCsqNiHb1soM1nL6xi/mPCoOo/roX8XPVKXZqQ62R43v+Y9uSrQREDhBYx
kqOeZdvVLmqXNT3Ds2RvuXaT3h2AfsYXrvOHqYS+0T1dStaqvTFTy8DY+BNFnPFl7urYv6eegvHT
/wf5MT29KMF8fEt07FzZxUdb3Ez4ED3Dj/Yp5gAcaUXj2Pws+6p11FjfVYyGZSVTVJV72ZqIEULH
ZFBo8nnBFxAzKTNnUMNsVjZGPCq61/kPGPgzrRa0ARH88LL81IBaQ2rBUuJ0q8mThhAvZ1SzF1AI
Njj79sFuhzMHzs1iiV2ZEb1Z6nN2Iv0UqOKkw7nEduF6iLDEwmi05XJuIw7cm3lsUc/S5+95xaPI
FROum8Dh5/wc1rBcHTZWpDj3dT9fPonfqrPdnoM2YhCK3P5UmDZau0fwKD3QNN5aXoTOntSzONrF
JTDiCy7V0Xhrqp1eN3VEm7oHQaoLYvKv17bKKcwxqQlMHCVBFptYh/YeW5piJYJZxnVsFykPWXjh
MUQw90ETr8zOWlkLnPW6M0u4PVjV0Y/leLyyJ8bB4xWO/ay+TNvAFgSHgP658KdkeTvCL0p8tQzH
VpOp/yhevu+aNE1pvtbF5vhHYg5IFT+kYDsGW+XGQdvwio29id3jVMCLrBxQ3b30Ge9GoI3pkUd5
v13QD457LZLYG0KMnoUNXhGk7LJcB5GfY21rGDAQ0jxkVyjIEhj3HmRYk3gUn35mcKWwnTtGcfDu
3DVMwYQA8hbruF7zOUUm36dvCHsKH+OOczd1yj44PnmDBmJZCDpiz0UUMbyRvAELP2/RWlXB16Nh
dFh1nE5Ub2VJXuwigLZkwPY8Lm7vfh8oZIjhTL0/NrNz67/TwNozIH5fvqmVavD+iukqAWBNrC8T
1H8+PhrSQp6El3RgcZE8q97EkiiGkaVpWNjbpN3UuQa+/pouO2E1UCgAy2vdtBRjNjwE+CWnZlpY
jexX+LE5jBTj3cvX4cNgH3HYDX3rccrtcwVcAZsHjGQFu3INj1OtRHpcT5jfUeHlRVESWwr+ZK2a
A1ehTbo4SfTW3nuke7DDQiO/WOEjkAAFvbX6J25MiPI3QyJO/IAVA9d99eXC4cWcX/8W+UZmPKo3
k8q3aPM5McSMgGAa0otbO0+dyPGwEnfzYaafjJJkttUsgkqkNSHs3+vPCpx6E8XIJP0sYaks21uv
sa+vSFwdy61fij9iez4Rs3+8KCbVAePCsnZL84jEhVTKNU3KDTX03OOzvQhqq4n4zxMoHYsaOJcS
XcTuCQY2h2u9MkLWnzjVQ97Eed5nseU1G6Bv3WyeSL2AWkMFLqLR4GSrynZ3b8wVpzx42SY8KGT5
JoKdDkEBuKzvBu8f58NyPRp2YTr1Q1njN9lppyhkdRUwvqg6woe8RDEeyNkOIB/MzHZrwyT57ykV
VC4Ct1PmYEJxrOTLBXw1z6R1wx7JGTZG8jcvO7anArVDV0zKVfZkd3tWWJooUui/8zv13CW9uK39
FC15EczTM9SDkLmtDwZLxbEMTgczNqy/WFueAKlx5T3YiO6Bc5kl01cW9NTX9yshQeDKmNrHNkZm
VOvccL6MjKN1Y0pjW5JKB5ERpZRBgEBVOJ8XUkC4Wq2WRTbYQAZgoYhIyboCUMHjyVZut4O9usTr
R14EZZ9Vunh+CAwpfZNu5jVAyu7/Hgu4iPRHRXIlIx867KiQQ/KaGVcLuS7ueMhikz3UqfFBStDn
GPwYG0GlvimmEir+l6qO4KEJAtJ54J3MVukwDX+C2eb4uufuIcyncv++8y0QKUCwxTHrj5+oQrrr
6liHV7h4G5Cd1JAiX57ROU4cTx88A0gZwnq30304t44HeVQ3Mqe/qx7cASnbVfCny1Q4Zhs5hSBw
ZLdnDfepRkL+EPNEK8lyWKcKwQZRIdFlAL9/29psDRsmI3bnl9xguVGp6aX6wuCqYwOyuPXDCu0+
6YoyB8POC/E751TvuoGlqvYQRhHv8UsuHOrFqdIbskh3Nl+d5NrDg5OrsC5Kt2tqHgz+zF9NXF7l
tyrS8W57X+VHH36W7bJdKh8V0CGavrXZUamx4pf0dMN9Q/4c7aljUEk+UcAdlcy6X86RgtRuun5z
oq4VGUU/+EiSfql129y7Xeid06Ka5A+6d5g+iztNqwhRFN8LxmFP1XLo4buYQb3yOio08GAhsg1m
hn3SkRRuDtmWog+PMMM08Aj4cqQdF9pIHQ9iL0trV3l49c3CtS7mS/miDD6fjHq4/TEKrtOakf+h
YfaSZ9Jxl587Iy/QalY34s4QCtxOoudXmCBP/UhSCAbHLGcIhja0UpJny0wQIUs3Wvm3VExsKmXi
3tHy+88wqyt44crEF+fkKgELiHwSmT8sgzEa/6mqYLPpmV7UYSZT4rCc7NO8wj2lPapsY8XVBwJw
6PCrTHFrjHtWBO6XEBDXZ3T9R+NDNZCpJKRtbnf5g+3bxVGy7BMe8kmXMs6gpxhSCY9qmX/nocq5
/LXfRQLMcZwMu7LJ41c6MpwP+ucW/z4db4gAQIG0u7iDYWfNRFmN0U9GsOoOjYZ9OAaTD/KwhiQk
hCUfXLCbxeMlYqGBMsNliYB3pl81tNL4104y5ckvs23kzzAUnKLo1pkrELbBctV1/bc9Wr7TAU4p
3TYvILFghSFIpYAcymrMSeHgwQstuj4plRTuW4VQxh5o7iSLz347y3s+nmnTt4WvFuwoOAzvkep2
K1kIAJ9kuBWBwAkZ6iMGyB5d3t/demScAcw3KToc6bqIaIoHorqwm+Y8LXn2cSoKqjhVtZA16LEJ
H+67vxiEOAZ1z2rhIvzQ5d+nuPouvJlyxrHE7hSXLebrKvKqyRYKiz3emZ2SwoKDC2YKZYAV4uZF
oVp5rGYIIVY1jInZcik+WLmtWimFFPps5+j67EG46GFyfrebxIm6gNBipoyIOLIMXVHkvwGo/3m2
zlGOK0VmF3DqE9j7W5rGwXOF+j6Pqpbzwt553jSGNyY1UZo/IuQPytIxy0vu8Zqm7owL7Ovl5FQl
4PvX49d7kqDmR7R8bIOzZUio4WTYniYetQ44PcmPon3YqpJqmNMT3sbQDm1baCJkOWfdDoFHfw8g
PNR0i4ejX3sJaEYYAg4sk5Rxd7E5jus/WjgvyKR1A2vu3qnPRMMyVr3cM6UPCKEdF422S/uN6Ne1
ZtXRivPPleFJwUvizdzwN2BWrOSS3mUjeU9tHqb2xkiO/cTt9IVoYTk/aETJMG5VHqjIHAE47sAZ
t07K7uuIz8r+u2tae1GTPffvNQZFQg2ZP6C7LvLidNRRrE0NuR5cxyRenlhFoIL5dcBxOG7xXbRG
tIDOGHXc3x5Lwm/ZRibqa9r/3Gc7/mghiZzasYlEgGWpza0PtxLqkm5gWjtliH8HzpGkqqTZs2KE
e+DxGTwaB2ZDIq/WHdo0W41pDo5MQYDMXBL3OxWzIfuFIT5PL3gbwzgPJzzhGqlyz167PbPZ74Lh
8zTKSCuVANJk0Ex3EU/oSJNp7hyRqOCKcqGAXbiqAg4ayylDbASlpMk2ed06AA+xfcl0ie98aU/9
uuTW6pi+fjl9fs+iHwcZggDp6zClrhzZjBVI1FcBsb7df9iTRVfvlEMTk9Ht4ExoTauQM2HVdyEh
3sxxY4jzEx/4DStZZ/GVINev319Nk2Q0aG9Awq7BLHcjMM/wH+f/qS+j8MnAO3rqdOnlhEdk6x6/
W3MxYRcPW0zBUU5DvhW/T6yHRn1RfynvHaEErLJKkMIXKFmr7MqQjriLuWu70RO+ogV+7EeQ+JYo
iFbY/bu2F5otVoffNH+iFJNF+d1ADpqBEaHb3V3JOhkKnXADaudIoF7T1MDjsJ1KEcrtGur2D7UX
6om+UUWE94++MkbBQBVMednn6d1AzLJE2Nk0B1fsZO1oSRw4Yc+nx2tsa4G0+fjT/vqsdAfMuMan
n3nUKVVdgOS2luxXCL52BrEzftjerNax4kSkhhFptZWq5OpDWOgfl2LCHKdIsJFqBvSezpP61Yfc
joiDo2pa1Qc13x8jLNxWpv2hqzT2/vNuA5OA7E1k434l7Xl9K471CYFsHMkIPLXrnpiK7Po1IWdH
xAq2+Hx0oQVSd54FZXGcRlENdgzg7d0uQR74q7lpw915zJ6KPtFe0LYVG6X6PTcUxxKWgWBWD86E
qUHY7lKqbTuXSDUQlYn/vUBD9BvGWqw9AYyPir4txWr3k1JEU6lrnitRRoXZJkTVXNYfFsgMIw6z
eK6Ln9lawAsdIkSJzmhQ86PbLDFTpXBwQT+n8/JvfYzG4jI/dmajY2Mi3hj6QIbG3aWOASO5uoVe
xkEzp+xphXkncVWTjpq0mBzv1k4uVFfrxtBx91TjDr3owmymZrTHg03X8snldFmxZ4bzPIbFtQep
Nb9wZNcvZhGoVz5rerxVE9rVItVm1R52Hrcgw4nNXAs8REc/KmGUdVcXJUUn/v6RDpZB1leO4gK3
92kpUdZvcJrdbyqatf0wo5qSqJq/cR00PR8xgPSYhj4baGUw4GluFBO8xYoIi1+b7MwhACZkoGWF
AqpArM9xttI5GvcvyAzlVDvQXnAidDVaa1ZClpZqCQgTD60DfSJNuwbf28KjRT+G4VPNH57AU0lG
JCvTpLWBQyKK3HUIBt3er9siDsRE8MYmYMqDofTnBlsC49vSoeRgXCdcoo5t0F5BRIhnoc2nhhXI
5oOXO5EEi4rKtcIqIt4XzrrSygLdkd2zVrC2CDyBLPM0YoFl/6CEZLs0TLyk2MtVRnh00/lCnhvS
TB27npMBK/jyl7OURw/vWuEMnDxQoDCw8GnTC/7HpHZLxkT3aP0SZx5k4CBSqP/yCS5OrubMjKdd
l1guk4lIfGPa+3Qr+gKSnc1L8v7fIEDFQ0GqbrBijR0vibP5VyPWa8bHfGr9GGQTkTgBk8vOiI4N
pouyrGiS6S8hcwlXe4VET7pzyeLo+SXwhMw0YwWT9cZuT0XaQ9pI9+UOoyMgQy0j+jdI47a2ljk8
EBcY+p066+tZEQGGDfxq4KH3KLVcpCNEytwl6pnuJIBWWKPEOQNt5malFWmDRTQghqAxkPLNjG2I
gpO/1iGwewmFQrNJDPsieVyO53yWnwwDdHgsHg9zVLqHTy1Sc/l+W63Z3AXYsGthU29Ke/VNydHJ
0Zxwa+wQPBRkGy/6Ve5hoWOsoQoMIlMgmk+OfqyY1VVCmYkpjvsOMMhMa0PIDK81yJ/LAdQoPg5f
EOV06EjMTHFWEYEBEBxPO7bFaJ7aA9nfp6StEaBKrZ7JZ2l8zRotGgJJklcsp8wR7ACpY2zojZNH
2uU8YZEFMJ9WmRnjTHciY+SwIL/r/xoqBbKliOxttDsMFVyiR7VP/Ncz/6k8I7hJbMfud7H+UYnY
2vJJ0PV9bh5+mkM3On0BF7PhunAMgJiEKjG0WgsYbknZDE9xTU2laj80+raQN4XP1zwmQw7K/5cv
o2nMXkfYT6KMrT53bla3i04eylWdOqNGJxcGiEmm9Mp5Qj7w4WiMVDjh5GLHU53WQgYQXWPfnt8e
KRNmgOI2RGaXVe2lG4J6tq+hwwRPP3qzsv6oUl8hgNn7TdaeI5X16+TdsOU9XEYGE2rq5xdC07qc
FPeNfZM2VcKCPOH20+jTE2cgao1PYq9b33m0uOirJTGCaBPRRRICKWXU7fpoVtFcsW9KY3fBvXvs
nr+2YOnObosIz6Dhcws2k+bqGRu/jHLNJzGVDN9K26if84kaULPS5gp4VtBvf7PSggH9DeLKOauU
6T2qbAb0gJvfRbcRyWFNhl+hquoaj0HSLP+srbLSqcZD1USRjCaWdy9BPv37Klg5gDufIKKC+As1
RPNwYY7zR2NZ7SiKoL+YurCaiRH8OWqPO1cK2ezMqlqnp481oXfKA5KUDSdq2OV4P0fpog0upG1U
SSZJhP/eetsuAnHZ/73h01oo4A4YGPi2JP0ThmjfXjvlV8cYi46jG1lAdZKwtzVD0Hw0KhZE/p7C
queh93WFKLIJzi6S0WJa3cbQpf1balhUhMkQyAv8mkf8qkxQ8ZQ5Ee6w3YCdsjhWTRAFc3ZrM7v8
lDLkvzxksn9gGcJJFZdOGmWfzv+pVL3zaBPNLf/wqtxiGMba3JsnbgfjYriKOBa22jLaarX0jdLE
v4HZh0s6oe2h6jYtpdTSIviuBHQcVgZle+CWOUmM7tw86SS5BSgPFcTwLMrubfSmOTetIkiXxBIB
Zt5A0S2/w3y8+XoEy7pRm/mnltIBS8uSuwjzc2jZ8vsbgTI/T0234mJt81y/Q+/YykOHRAnbcGY2
6oKjXwxqTA5ymZoGR/SI4bUmlQfZGQJI7mKdZCH6YDZtB+7MIg+bnrEiggM6jddc/Lnw1kAv1CNQ
fOEaKJFMOiRoQdg4p6wNzZ36Gvh/QxEEUzSMX+j1hJOOnCeLj+LENKzMXgBFPLtN5yOsWoyLX0Rw
knAJ1K70gUzI69ZNdSE2HzOr7MRy2PFDFrTQO7kjmfG7lCFdcRV9wA60Cx4l3FFBRCq6PVak5yMc
2VbK9JUgX56SlMPWDOinpwOuNV7O6XRC4SCbnr0rHeINC897B5c8btGUuaJgE+8SPSFatiVi8ZSK
dYIsJs0KX4bxymf/6tLfG3s3aADjqWFtUh8QDbMAJzwshaSSIIJym6jSsULA/asttZ3UtKaz5/6G
w7dVi0/Won1TWLQkzM9N/nqOh+E4A+M6HWMMCShKEZxKOihXzczWQ7VEpDdjm5/H1n5Cjy9svWDD
S9zTBgn6yqmouoRfMmx03W4ZH19cDbVyIdN/fJGzH8eJKLesujJf++X4il4ONNfTDiwhykDyBEpQ
UNFF9HIwxjRbuHzx3m1XDTEd494lWbwyyVCA+50IGCfdIrLozlHpm6hNUyyniKFx8IrrOglsV9YM
JsWKh+zDKMtUNG4DKQkIjtTzfQua/kkcmuSYk9GH0kNv+l4aXdMAu2Aj809UWP2hY/wkIxuVNomr
3ag7UKls+h2Mga9+SOhLEklLYdlbvdjhL1MICCOm6uAWpStT5LOaXM7BH/HYpFUzt2bBZi/6x4RG
L1v3N2QcHCGsdvdgz3619Yg/eYoeRhKOTZwojPNwQD4/XFoZi56Bcl+C2kwlCJu+sddPdJfJpmr1
94KQgAFUHk+dYuBhaIJESgxDjQetFYXHeKjh6VbeoeH01cPoXmV80zXt/Z85/VbqYcqd3a0CdNzk
zBF0GHcGsgmwNWut5KwG7EKf7nJ0eUVBXKEzO6izlkC98ZPkBY/58sxGblnfSfH8m/XPU2n0psXh
suomQ3Qhe1tnWKUUapn1cpu5+PAYBAdADhgHfGqOxBX4R/kTSP9Ak706ZjGxBRvsJtUK1CpzP1TV
FqPScPTVv8i52r2xtChkK6sE4nthEhpVC33nZnKH4hwzSgmuc8r2k6dJYWrYMZasIqzRa+x3e9Y=
`pragma protect end_protected
