// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UqGBC65mio5omaAENd1TBDl440mB8DPzBYSuAcAKyYsztoxDMmNfncma2DjbEPA5RiLCdN+GsdF9
SeFxYrmS35cxXPAgQbgFncEh3VE2Qjlas1OZIqu7U4PnC4fzjAh4lugp54rqw1bDfUWmlhQFSskN
gbAYLkIrjNx5Bu13zLuT7MOWXXU6hRRGuM25DBB1CYlpgkpoka/YHv7P2ZzGouIg4z1QTxKk3A3P
aiZqaN3OtbColQ5cJcH0QRI62Q545pC9wbJaYdUWXBVtARc0AgDtQUnB518Q5+L8BeaRyD4hCEfa
dIR6wajPmvV6ZcnOevArw4TF/6sIdMZpLHw/Yw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 50720)
2iAARmh7ppJa0D+jufnuGgIAFC2/zeuxAR+NsVubrieybzlZRCRRv5Cfsx5qpQIU15rpyylHqwXJ
peg6tMavvWyQnxV+7NFCvKLV4qvFS5et0XIfQtEyj4enTsRX30v/efpPtXVI+3j47RQTrieoMl0m
prw5FUUOGB7l2jQ1Wf8fF6OpUzfOE+nzbqjDY/HKnzg3PiEWDvES2a8CfCgCafU9QFgH9ZXBrLRe
8yo5LSgLS4xXLWOfVPJUu/La1dqzS0D5GZBbiirXAIxdADVxrC8CvxL9rOQiRcZ216VM/7mAYEea
jGK7IAfTf38wGnd9fCYLj2rb/Lm2ZTCJY8srMiYgsIbD37i3M41M2EGo2y3GG6mC29NTlFr/5GKY
NXBjySTRjzztNgYVt5gaGhaQo0A2wuCi68j5+UXd1bURHVxcBs0HOf+htsVu0Bnu7HZUXLe1PR0G
yaXWQ3ZcOVZdpjJAoCM6yMg/hkijmmwEFcondf8H34SyUbyUPmQcjV+A/8p9dujOuaG489w0gV4g
Z3p8qfJEOs1GQa2PL4FNnzrglnAIJmSNCrtzM53SUm+4HflN5iGT83us0W9eT9c0ALyDbArBq6UE
rR+O6TwFG/R/mCp/XaQCzfXeqsMXWo40FkCCO1HRDumBV5Qrx8AkZxwJvv0VOHkECLtHlM7zDtxw
//g3m1Kb/Vz2B4+6IDE4CexQqJ5Q8wJGka/zhzuVZ+5oEtmeKuypelKjjDOarzCUqg96u7tY+le+
9ONO+aEO6cIulauj5I29mJheSuBTPNqoYuQpAV6rSDugXHP/XFm96St9q9Fj2qhno3xPg3rxuogS
WmFIlJCD79GgZOoHrVNXgUNBaZkG1s7wI7YJSLwkJ0nNrvxtibXVomDW+1CNDUgkPVzS1jl3nVZa
eQ8/I3Yat6ww3tAmWJIhVm3KoGaAwG32vDkiiMkOXUGI37F2OvYWY13Lov0+pgkeJpsNhtUOfkbz
3Bf7gmRhFm3O9oo+uLTrbDMexjgWoKpEWwDlFtY3PmZSgQ8uSUY/67JuoQg946SiWk9YSTL4RpYY
dd7Jgz96jgvkfTFNw1BIcSaUKrdXDWd/WHll02ulBaaKIuL3ftIy5qvOExKh+17WLPDqrDy3J4HD
gjZhtZCIx8hImAD1ILrfKWMaKBEXwTlYpa2KfzkZIls1PrL/DctbV1FS7Bi+L3C0/J0rpZOhyGgS
T30H8227brslxSkQBAn3rZ3YCaSW4mZYfo1dtzEE66354AEi6ltqNr4dc8FwGwceuZ0nRFwoP3hU
0G+MEpvzqW/7e2KdO/yxVkur/PYL+D3ISLCJgZJSCjyStFZ03LKDaPGTLkDPzAbt9LZj+WcrIVNZ
jHVykjPlDuICucvLLYZSGsEmmNJXBTlUIxakRzTbVWBVMFrzEo+Tz+D49dUY3ayI7+4noWFSA76u
zWTm1Lao+M+qoUnzhgMdn96jwMUCh9/vR2XuzyoE//ssyym65ow8nM23xAQdu7/GAyVbfqEEkkLg
6M4mb8N3jkZxdUw3w3KxohqqIy5e3vV+7bAlwzA62f4eN0uv0kfESYaKIiaOzaY6kTNOcpsUtORr
wRTVcOpkjlyxV9AStfvb8IfMbTYCogycQiMnfXoSrUdKPX5hrk3LPyaqGKFQk9gF2NRho7Ko3MWH
Y50VV+Alm7GNiVs/+efEvXBruwCePsjZU8SZ6H3ZC5c07cMbRMhP36IPpWox731TqN8PLjcUzLWZ
3QOXuXstB75DcQSWceFh44R4jKnWsltvxRTymknYHacdZ0aoAw636NaxjFE9T8DkZkOe6k/c+rx5
8fiiMR1u3xdvBoQO5k1HvJlnxpV0yAqSTRs0W1HCXpgFYYkD4dTJLA3/C4gIot7lWw1Zy8LU07t6
K8pEupF1baoN4NHvt2xPvi8ttRG4g7sDUsg/Fu3bYy45poc/V5hOxSZmqSBsaj4tozbtw8vZ4Y1v
OE6fJjmRw/ixQv74ONk2s6tfrhdTJ0gWUySHKnHnu61bluizuQv9EwLu1UfH0ObdWjmjZTn43I8/
AmLuWS8MFitpApAbgJ9AJH5tXzEA0IElKVYSPtEaYNDEvfcY9MCQLPUOlx5ZsvD3WPYagaCjzFnV
Sra8X5HuWUMC+aIcNYZ4cVc6KNHee0mhIgqbrXZ/KIDb1BjwCtPazQLwwRe3Ye5Kqc2dYkV3BkCE
wqiiB0a6wP14/KKwAvoP2A7gUdi2lKHu6T+NKAOO1MtfgC41iqQkj3h7Yk/LpM3iXw3V+VXp96pv
uTaH6/w+PedZ/Thg/3EPEyPwLzrH6ZXWyxUb9SYhNhkI9MhAleXOSalmVXH7t6FLN4ZUa4G3VLIm
/PxaADO2FwWCpqlidN2SLiLNoklN0f5JydDY/9THiHatpSIolV/S6uMeJT4Sx0VoVTdhWSKCu7xa
VX8MC0Ukd9M8QykQJUbO+l1EFgHqKiRqcws5GqWCTimMNL8M+e50mRHIK+d419qpf1IvPx4SJYgf
Wjn2j6p70UOnJ/Na1y12yImPq28vnQhI0HnmMLgSKDHmRZtNf79FXOYEysOZg0cGJQjvxDDGqpfq
lwSvAxH9qMjomkaTd5HxI5mnocYm0hSMoWv/89DnboJukP3OohLfl3KuCN9lCtSsRcRlJNM6SiTs
BRrRflGyusejPsETX0kCLKzP4i0DMLpeQYROu41DMKZsS6NLR5UL/kxeBAPNfuVAtz0McioNlddG
U+w8/wetKCxYKikH8n4GcBpYg+vu56wvKbl9PCFQWIfiU17PnFASSFVfXGpiJNeJZIX5On+4eM6J
xQ9rH13+yugvC9N7c/RkYBp9Trh333fINWOCrbT3SajwamICcTlbqDw/CakcgRfwSFOTpHYWC46R
mVuORaDkRJ/sV6VRz6VCHwWFjOk3YuUH5PjEtakimfr1N9TuUm264EuPK6eYHeEQMfMef3jPKzoB
5kPETMzlx2Fv/bxZGOkRX11LAqD44sv70MuVT80WzYrvkykgMRLvpZPxaGRpILKCV9ONpqP3XVvN
2SgqI1CTDrRZfACbgoXCW9e+xMPj+h/nq0kFDf6XAYsQeLVBqJfpL4O1B6WVblx8iBpgBE/vQOPc
kUJ5NqshcfHIA5np4PBQ/KPG65XxiFrvOrmRwO21aw+wD4jTkp9IShJsrwyLbbSdG1tkK7KUaM5S
sQpE0NL7Ltbg4tBrOkALkguG81XCfU3JZohHNnVR35yOARuHvBIaad22iFmnn/dkBB75PNMbSXYv
nidcft+VKz7Wi8iy/GGL3+tRnssaGt7AWi6KbFV5OjgHJSswtjTjCNbl1tdEJA1BIabScs2EkBuH
QEF73EUY0osooal+IVgqPfHSpPyxKKCMxDUB/aC4MBgeTRJ3KeLhhKSwj3567bq+JkG/DRee6JYG
dsj1cQwlt14K6A4lCHXVmqOibEy31RYU7nktrCAWyMXtnnje7SKU5os99HhgDRssznxxLJ3/Dnfc
xq4PF3ocwkoUrVlbDVwHz+xBeFDugHWBnqzGo11k+mDYbUYw7iu2l7ONOGFJ2HfK7rRvhaMMwB36
5h6jED7TwwY5F6DrU0NH+B1rWCLNEF/opVSFGJ8QAub6NjI75HFdwYVzaKclLKjk2Cifl7mSr8kX
sYw+X1B2HC4ja9r3GBxAd3BVjyuY/nHfKH8a1QOPoaIlEBtHCMzBmldulxaOBDDmJDHZ1NEIV/4d
0TuaSVVgHuwkZWNMMUTc4RSPgPBeuocrN/J5kq9LH/Us8qBg8FjLnUJxWWrBZCFsX/60smBKiEFz
XdXNFEq0hjRV4krDcKwUE6oaaAym2AGdxrKsuID2hO/yREFSuQj8zhAytnf0c0upPLCdk/FtP+eO
LKgvUF78QjRev9hHVZNR6AwSTE81ksJUfpzS1hfTW3qNXO1jcI+cYTyrT1ZYsmfyQLzAuFK7MAIV
Rv7+/eOAcJvQdRf5+kNnQMo3pjzCdPDsYJ6eu1ZRKETo6WRBYTeeBQxOG04Q6D8ds2tRqcKE+GZB
V4FYAVzTia6r7tUFKI52ut9PQbak2S3JViHOPKJXxGQXkM9KMOzVfEN7jmba95aO1pqTRsj1y1GS
rFJTpvv7dNbowlThk1xat5LTfv/gV0Um7ZjnkAeqwrSX5q+cFT4JlyQX4TzdWDLo0OvEhLsl1TDV
TaOIImJFeOMJcSq2eTvTLqJnbtDX5ROpQvYBGkmCkGDjgWB/0Um40S3euy8mnc951cjuPoK5ImSM
h0NFbkViOge7vsApfgByHR4nFfmFVtfs0cfsADH1LQzo+d0k8Nb4VZXglESEtXFMsQewe433n42h
mUPuwyUmHi/2Kzm23jM/8ahaY/BJFnbFf53JEFvAz6+MKe6rxU79lnXeep6VGnJtCzZi3hi+N7o1
oogBajORlZRdogwtyvbzt7jPO6EAmwfu+IyPGdXCHj6zSg0FExuGkjDbhFB8quftuPhrEocgUXhe
zQz+/JnR4izrOlHt6JqCnM622ZhaVvofuHaFi5iFBjqncK5Px24g7swfeT3zkWeJ3qfHinvLGwoK
qSUjLXAPV85KLCIwRPKDuF4jg2t+ly0pBlD0Thqt9e2uB/xdkcE+Tsy2A51jGs6Gykvkf63Z9vM1
rvXtt8ZKo+sdmvh8n/Gui0X6ooR2hC9xUAFY2obPRafjl25HLF2X3Ym1bxgYACBq0HunL1uk64HB
uvqt1DjdHrCprTNO5MU7jMaokDMItArgi8BzWvrt2gbNvTyNmiKX547MVRcMjaieVYi18/Y09CZn
LKqn8RKBrJr02MlEyYmewHwhVIaS+gnDGHHYpxsB7dmXDTUAagXT9uhCE+Sa5GduyleSNwxtOX6u
iegTXq07R2prPWwlvG2Kvjrpx2NtV2x7aGRTj6SGM+gdZwiQlROO+fWkZ7N05ewzL3W6Bcrz6SQk
1DwkTz6QqOKRGQN/tdBarKzwWZvO62RainthTldyWgL3kacl6ZVBl2n4zhfJGOg2nu2tT179l7sE
3I1ZjSpge9oJtONYhFtT69PEtSdsSFV2kN+173pREfBYsLBkPCRv19LahqOJimGoCL7D8+WSJ09x
+LUSEfsAOUW977MQgEHaXxc+8kiiwvuiLOS2pnNn84TJpB+SbKLPCRwZMnLrFzxoUfIHigw9+zRy
i49jiaW7aBTNfFYr/KnXp+GE5HzbyUi98wwhAzmnNSNG6sAHEgb4C3gnDNuSanGqYSdzZlZgiSw7
vAC/Sc5QcyNhXfnNggGxzIMhVtkkuQ5uyn2yhpU4SBq1Yad0cfc/azq7A+SFeeBlRWLpEdqlBv4+
DIpQ7v4Qo4Xk71cjZ1TD8DsWSxhzqYWg8UhWg/8QTbH+EJk2VQqtx3TO4Ae/C/YYLkdDIVJf2tnZ
MsYRQ4plXwBD11tfBeaFqY9woFBrV56XdX3rYS3Nz9qk2ij8xUcApi1CyWBq3UdJoVyJTzK0eFY+
Lmf+aLBbCJiL2gLHQx2ehza0xi45CFcggh184RldlggjG3B4hJOJL7c675VTI0jFMAvv/O4RX6dd
Jw4umXJmVvIj4oIuaA9oYFuQgIVhhR3OP4xPPKtmpBZzfkaQBCIvbQNtlrkX+U19pWM/gppNN3OW
cDR77qSPvJ5gkybdRWDicurMf6wrw4MHxzTVF0sM7K9jQd1tMUcfIZktzU+4QTFR+nZ1CzhpJBgd
r05aDmJEXT8jOr1kO81yslmd21TTFht8FXfL5rdHp8hIpLQcYbRuNx/PhfiGU2Z3tu56UtpIozlQ
OXHTEmJ/7wKKaOKccJRsvrZ6KEMMh+jnhHig8fGY3By3N24Cgan6cDv46Kwc3HPx0S6LErkRvbK+
F/ZL9P34xuiYBLAy/OP6auXctQ9mA+/nxWV4WTXPBACTyQOrH71wVclZyzwe7Ibv+7AURtPiwsjj
paz2jiqFcthoc6kBCrCrB0AQFECJwuxN3eEVonsJLTUGuy0vX0UnrDpqaptyPNyD1oMlXwgob0zV
Fr7VDy3zAvt9P1pNIQdrxlBuxAHz79bl2RAJfYsFiAl2IwnYR41/+edzERkKjJ3T4qMtEZNd20vB
C2wym0Y2ILNChYvisS6gUzKn3wo3mzSo7oeF524q9NUUtdepbJzmXOJuWy1Nw5Sgb5VcRYY2hD1M
b0UxOjXwgb+W2sdKbRcgtgN0ppx9dWgFFsOYtgPp/rptVjwL6B0WwUUIo44ZbUoEksJKk2LgX7f7
w2Vd2NRBw8FEDdjkrRIrjfcWAXpIBK4iR9ecKBYwhHEDb8N8ICjq4cBhLDstidvBXxvgFc9Hu5Wz
P68Qqrp4odEAVEmuowJMrQVvFGjHWLgx79ebhwvinCK+JfdJEBYj4dNbBTLtXydykDX2iKovscWJ
hbmLVzSorqnrPJr5gzxoAPNMdKTmNSMAY3arBcCCAKpmAYRuy4jbwWz8UzPB1l7D95aJv6GeJ8yy
dfVI6b18Yb6/Iiqt2pWFrFGmjuPSeTrykH++yjem1GPJcrxohO02CDJodqcQD1a9k/4rReibidvz
2ibNPAEYF/VUV5abKYJsAe0witwRLXEvGxzwJAgvNGf+DLoaXWWkncrYbvzepY7yDoUYJSNVgl56
3pwGnNunygHg0j5Z9DeNJ7pJ8Wy3VbqF4/0nkmSvag+6F21jvfTSZww5QB9D9cCEruxTXj/K+WxF
HjT6Fp7gWt/IcR9WVky+ZbsQav87MNYvero/20o7jNIKQeOnRH0rfeyAweg0Gp8zXDO3I27YOx5X
W1po4JcW7p2Wo++4dWEGokpVH3XwEYodCqSuAhUA2fRNqubcpoOXJWZwRw4TKGJ0JMDXca1/4UYt
bJc+H7fZxINRV3dvnQDiQpiRs/eA8qzZ5rK6aGW2GEkTYufsCz1V5ICRyxaV9/PfAn9vAHpbSjgt
OTVooHB0oVl8uOojsE2MXXgi8gaEeNEYDDhXeto2ozAbq5yUDwwQnB9xqxbYGkmZy+Qm1uzOnhcF
Qp+3xZe7XkvjTtrAl8eQLSIMeUzcLBkrcAft3L25KuoAEKiznDURmdGKvGn8kCJbVLd8/wpOHx5Z
T97cxKnFnuwXQhvzJN+m5GDlj4bg0e36A0NpXrp0le/dofDFZ3ZDg/MLQJ5ALTDWrNTMwE7dPK0a
hjnsrqFlU5GvFuTrHrX4XFQy8YNoz+nnQAhbC4I/locZRIlQNxmLaalbKFscUdygEHY7X8Rr3ZOE
mIOM5dG8zs6krhM+3Ue+IDAd8Ojkd+mmRBp6r4zu78vh1WASF9H2+l4YFMvRgjTqr5a0rePCs10c
2M78HGfC7JCkM/JHXwn2u9CatVj51zDQfN6d+ij+pt+luBW6PIXx1Cea7bbeCjgidb4wEzV7OJ+5
k+RBy+12LUWlbj/yv16wR3uOYWF/KwED/0/GdoZa/0J/bTgV8UP4vPjUnCAewecmFtmQWdNyg3fv
GcoFIDyImK3R9JA5YicBk3Wvm1n2bV6gL/GUjSIlhF98opSlGN1gGB8sAQrBSR7/ehFEkcGk56ZF
TIF2CG3jgkDnt2+2KUTTCwUIe+p2vWLrbKCDkj+TuGuWqSZxI9cHOx/KFhQPvTuHkuYIEI/twXSA
8PUUPvRp52AuRHNafQaB9SI1Wde+E6lIjF/MoCkmgVd4u+99T3plGF9Uyxedi8dzh51MiXTfY9SW
W+JkZ2xZLG2HdWVbqCvoRAawoR3AaX11Mnn6jGHcQmk49gh8oWqcOm6kR7MboJw/rKojaSzjkudm
DU23nwNQHcXDbJDfDHWPT/sdwIysPVopO2rIGlxH03cxaF/URuzDYWpixm9uUpJr2UL6yhl4bVUv
uQPAgkg+IdC4uoUMOo8Zpa6GsrugbvRfa0sI1I//7Zp3oDZh2Ih9x9bJl2g8MccYmscjhKgnUGPh
8b7QqldWztsTbLJ9TV4XrVlGYVH4MR4Y+2y37v+y/KUPnMQGsydWgCkIKPkvtc4Jw00qPSlx7KpL
x+3u+EkCmcCSUZl0fDsn8kODJFVGGzmtm48B+4q5kij/fdHVO5nnjZIwA/oAp27i9YoLYFM/uWMy
kfiMIOeDVZv3DVSkYnQTJJXodHeE97ILgJHXe3Sd44Uf7nVbCm+kCcNbdbd1IEPGzGtEMatKLsyG
MzLlafY42gBiudnwohLnHRfaPsh/C8dZY4U9FoyTa9qEcDqOmp2Rq9qsMB2kqV6SfUYdEBznLu1F
t22JaDlBc7D7C4eBmz6KNGXMnwjdTLyJmZAhVfhm/WVu+Gb4KOwJlWIXpNvoz3uzkkfHz8OKor4f
/PJM6gQwoXFawoEUmassECfx0rG7rx2YDZas5GSxfLv2jtFnEIIN0uWSMFDxy8d6ksPz09NO2cIO
+SA+oIWMQXMBK3Hapfnab8W/vfl0Lsdz01C6BJz3QNylvWLCfIvmCpYxFmbEL21evvoBGZHd4q6D
QWLvvqNs/6hu2buKrANLTs/IqJRq0fOzTXzJ8+L06ulWqo8VehMXAYoKvrEQOjDMUJH9GjZ9b1Hb
AtcHoRNbmTlDbdQ1DBvu7GJYI/3yn8Ut+Eel2HbY7mHQtYolSa4nJMqPKPsd+BgHJjZ2jOuM6dtU
7io6FhwZQ0bYbbOHPYmxPV2Mak20OpLpjO+MhsKfhO8vWTkRkn/36xK4l3KN3N+fSNnzfoPc/RCf
VCW1mm3YRINI4Pf8s9MYqp8RAfzxUt9badcqjbCyelN5ri9Sl+XNWhIf1qCvY0CLWqlmFjE9eOAW
beUGzad2dSJHXzoCF49fN3KrIuHVcq6TtLTSGG0YO/zwh8m+EjxCcPR1VTMiTy5uzIsko2rXfVY6
7CYjEkHUBLCl1n8TtvtqohvK7nvJnHkZzSSWNoFsFe54MKiINUgQ2IKJsKgxe0yTL4tZdYa2EHB/
Bg1qJjGgS13zHGnru7FcEOJkwVA/psrKHlr8SDPHB8KFNmTMHCVDpQcIe6SDU/wKm34BtlVjze4t
hjPsFskyqZsR2l3kfP9yqNWQjXlrtVErntkgaqfJgV2j0gVY4SAgBHkgJTH9FLVWnyNzESHmGboY
VpdcwqLk5liAr8QrOt9n577tMW0Mndy5AVbojZb9hf5TZELySEbIW0JzD/kr8k8B8/lu71loybYG
vHBlNyLeNihYklTqEDHBEcJ5sEjIIYe4VvJ2sLovF5EvfnVermXsh1Vt2PdVwwzHefNFz7EZfIss
UNfe1vOqiNWTTMpxHT6xWy3SIXi9yLSNN7shnguyfWTzVYb9ncLP6/r261LQOdpx4vrWi/UwLb19
zCeIYg/I/gv79NNprtszs6mcZvvli+uWB9N3hcZJQwYzU2ycnx7yipbPpfgJ1ouM7j9glUvc8Zcn
iUmhOWkMuhkvkGsSAdfYv9hXSFzWfSNaDC0CHzITn8f+jAuOR6aChKNq9NzmACdxEE7qL/FpKQGX
osUJM7r85nJ5+mQWeXSrPZt6XLmYHj26yhr3anOHRNW6yAdBltZXwRasFeJi0D6GOSMXIAxuWjwP
3OQWOX6SCDXq1a8fVPJ6lMfSNZcLWN3zOwDmtRPIzkmL5ySO7g3hAWMwBtGJjfTWLmCs6tZAU872
PBTuD/RFyhhHwZOj1ZZzNr97/ePaeNgx9K0P6MRbAzjVqWFGZCBypTMTf4jxnx0tX54XZxszNs98
YK6L+k3+resvDMUxcYkRXr13JDw0mC6m9aT7MyOsJMlAUMplB5y5tIiaEOm4N11s+18REWU5m6pa
VvCoT3VPoqmdTx4rkwqXnTzm9ViW3Yb0Bxy+A6t6zksnpOXAreGmp4Dnr2XulCRmVtioaKE05PKa
+AljV5mQ9ZI/SXMGOq3FCZITsEJ0NGLUMyLZ5DPij8ppJPbIJpK6j3PnltjEKXHj0kvNI+ipzJDC
pLX80GlrJJ+LKl0kRTeKUhyL/AC8VErx2qmxtkjDVXFzz781P56ULUYQcmDaP2TPhitNDfBq1NL5
0gT0rQBo/oIvtssEch39bs6B+o/a00Z2DLaCyE/u72nWhA9oqfYxPvY3qF55ijK6A1utbaazhD55
MFdgeQATNZaOIcM4TCLXl3r1yEnTH92ZpusvtNb6kFEZVmS15Re5ZKv1SinZr+P1wMlh4c3hKefy
pInvvusuRomPQoklzNSRCkKAVVUTCIR4vmZj4Wm5RWYcxaOC2uZLrR+LgA6HjsYmzWtMn3aSoLzo
YefoW6n1hZvj+dheHHSQ8wiBI82r7WTkcFQgiMZaBRfy/NrmCqCU+pqsNGqKJx8x/CcUc2o+lZj8
IZCknT4jVRod0cOjNrqCmfkEG+9OdpWfs6PPDRqrZVmv4zMqTBaa6+garlSb/GbP3vsMZO1ryHS7
dbsp1nX/8Ffczh701lR2GskLuQNrkGV2LXjg0uPUtpeOyXra1zism32NqULx4acTkNpZ5cucwd3a
dg6t9nW8+y14KPg0mUB9thWkNKIeF/5LTD3b2L7DOCbWOu3s0F/7djksdQKC19fM8AykVuKW+0Dt
XyyzvzptLhf1B2NPzaxFmOxFREaCCAoBI3mXBP1GhUlXvPTLY/wp3q0I5ajq5xZwLrdldglYzVUJ
TJBYtCM6L5eQkjSowyE058KOGXdRmRr/y5mk2Vlo0I9OGdwTR5LHSt5d+JVPfbUkZaqDohvYbo0R
eyp1JA12wdxf134rkZdemlmRur41D3gkioktHeU3PFcHm9voHL3ZnNNlyuE64x4I4cTd0XClMHJ5
qfMCLa1vxokdJTD1Ste7hrPS2BF7kdJKt37dyrOyK4pAp4AP0GKUhAVESBxYcesJ0+OpBo0YgBta
9jROOsunB9k0kpntZJzGRXeF2TO/xhyJyvqsBf5hyauP28mZxSgC4y0BDsznqhKOp6a8CKNp+7RS
BW5pFP/AuQedrbDVMfMNjFdblJlg9Z3OTi4PJdSF6FtaiRg8dq7Wj1Ajc5z6OCqw7KfFEWo+GWYs
7/zXuV9tf+Rmocw20HdFp4QjbPc1bAGGw+/1NZLCSeD0HxcSHCH3eCXr2M4VW/8B7pqtgjDGohCm
Xsw/kcHtDiQQ/EHMgBuFv1ErNT36zy6pYa1/AkCRSFVLtMdOi1Rjws3nTB7+7d1dVNaoYHaTOHB4
/+7lZkA7ZGH719xbaOLQ7QiFD/MX9P68TgtgCwUZiHz9C3Gm9zzXS7ZwlGAK7Bl37X14vciTydbn
7mA7o4O+gX5hlHp7TIvglT429P+VbVWG68sFYbi/9FdM1JDwNbNaPanS43fby5vbrWWmaNiV/IPo
yGQY8stzuA1/bhf/q/jvUjL/0z+o6CSpJvLXyXLdGpMPgFpd3T/XFrKVO4SqIix/+bKgcY6YDCe1
sUj4uIqMhbrxCMEjr12BYfs7fqPyvV5i+5eAXf9zCHYGjMKFAcG9G3qUET+eJWSihIxmkqvypyCV
yALBDmtInP9B82byhSBhWwIy65Ux2ZZj4ZEkzJqXv9W8C9XHHNZLUy4D3LdRK+JL2/4VBCk9TaAZ
R5rE7gBjBgbU4r2qdnkEYBz2x2mRtQo7n7zqUNkmAtsK58YAZ0qkb94Eg5Bym5BdYQPuUSo1oGqv
vmBgWHxUph1SVnVt5SFQgUatR/SDEWMnojYO9LMRMvbIqMXKZq/3SNJg07AipMAqnzdS4m0NrTXS
XpQ/7DntqE3l8RbOvHAYsHolxyN838DjIrqtK8/2I8wbiZcmuOhriWCUq1M+aQOmk+kZ0eQ2wXC4
Uj+Tm9A5CtOpND2kHK+EN0Er12jFdnoUHCW2+sttS/BPScXP7uY+UcZ28zTSZeENp9yaO8ItkeKa
+weut2IV49PU3F+mjFieG5nqO9nkdIvfUPlYJwahroQTwAYB3RIN5eSnmtEowKKnouOYUxHZGofO
E1iRJ7U/jki9s9a3iNJsaAHYRKbEprgNslCzuccKIepFnOZRQgO8xbJKO4izvaEGQe663kOXM0ou
DH3HnXBRZvC8RHYBOzJs4TO3g46ZxOHGzAvXKeIFiC9XNzm+YbE1xGhhWC+HRdu4BZRc55BO4uRq
MU+NK3lTJn/9qexa4wXfFAxM4s4meJCKJT50PkB629YDVQ47R/7qaNSdmM16NImut+wbv1ywbX+h
edLY83K0I4FkVf7+VNfPRmSfEmH6oC7FiUylNJbt5jNmtQ0vmPehWThWP4ZA/L78234MvxLygB27
79jFemRfC/JM1rQxEunrk7dvxpjwXdHc9Y4ebGxmcDxnGJfxC4zxLoNGw+UZIgVLgY6opbtko8lF
dtOzy0nRsGNeOk5Ki7fG7n49yFNd6IQZMYwKZFxnRSPsJOwGhl3PWjK/iASCsIjTdXwZhJB+ZeqT
Dn+Z3CPM2dSyeKsWUVZH5kp9BNjYXJCNg+ieKCFhn7nDct44EIOS449huOcatm6E9coxDhayu3np
YpO5KjPDSNo1jSMxYxsJq5OKToqURJUp+YVsyyen2IYfDezoT6jk1YJ5Ko8yYlGFEWa64dXTsTm/
wYIa8TfGDLSDFWyUVuzgqS/tbY9/8vLwNpAcGxp3GZNqdJlyXfhRy8iCDoQ7HXuI3EGATivD9+cK
67cIO2tCxB7pddzo7aDDK/ywd8FnDWGpoZZ+j8QqlSr9OjnwChOQRuxCD2ImwJX4alTYGuDt7dDt
kwIH7YX2hBTjYm9t8HuLkZQxiKZrD6ivMaShBATbAPUMnS9yuz2UbNKyGfeFobPZQcP/FJUyQpO8
NmhrprwfWwb2rTFincXfWMwhUJU3LmZR0PZkK1RTirmWaKz9+HyMF3REoIQtsXUKOpjWuuFJbvc3
V9zcOD1TEOyfoYHitWQKg9xNftkmWbDsYD+RI7AhKVT01uFVVadeXXpRs8cJ7XB2LiMnq+lL9/F4
AobYCC5viy1RZvN1060uIQZqrodFMQY/CwrQN9WrCw3iOXkkaVfXMyCr/PlXimuymB9e4kWXF16i
q7V0C1FtBnsprrQ70e7y2xv2uu+Yz2frA+MipIHSc+01ISJs6OJzZIAn4O0oe/GtlrjUKjZh9pYZ
9xZVU6lqYuNcPW+23qKYSPI+YQ9QGRx6P/FENkj25tGXO6PkRYwORQwWUI6Im9Gz+LfxAVJtIv5A
jDIxGYhhvkq07JGiVjzxn5t4F/PnhTSF1xE3VHrMNsCzUreAtYbAW/NHUbwLsvgfP8MuikPKtEh8
kGha+P3kOKDuTZ1QvXBLmTF/hx5SgQDFL09nBHEcbDbk+JXqpeUjKzRn69JCf96y7YfOTXYMW0xO
8kx2SecreevGaSpoyIqetzpLVyBgZvUqOufFcYB3v4PU4ibA482oSy7eUCpXp97KrUgDzs9ZGTkN
X1uzdgClVdCn2UAUvlCzYjrCdLf0Ix+uTiVtFFJmhvz8PmjWpXHya42lXOxO+EnN2o7NPK9IRMSJ
0eRgjGXaCUhE6UbWLJSpJmhak9chNJObb1HCsqF1v9Ny3X/IxlkmXpXby64KLR2de+QJsYsVMUBM
/4m7ywGrYYukVoVVE2JTrMZFy4Tgx7fByUd3kV8rI8ybSHxcin3eWeSN1mnYbBRLmdZ4ywbfdzeg
zSaKDF6yHsRsqz9567UpLHjtVcic1lB0r9lNIHGJ34/g+V3zIA0bIIIWgiWtquAfoWAEvg7Xr9pM
amdIGbNKWvKrOVWShJTtZzY/lUzIi5Rk/5np75N665vpSIIMhrylxu8VwB80HSozQHeR3wKLm22C
s8giRVwjs28WxtqTV6qo/zkJdEyo3kBDwSDkpYkK7POTX7zIz3phEpw2RU6F6xjkWUBo7V4pIsBB
rIqaliIFw/MD2rQTMbDWxYnUuv9ru9yQV+UGI+oKaqb7Qrya1X6feS8taAJO7ZtGCnVwblrbVaks
9LyKoEQauWTAZ+9X+wJGRzQKWzFHZuO42bZvhrDB05xD0cRqKQVs1lV+ixVEAkj3Y/KVLNBN0SEy
JtofuBjGHFC81GLpmx+VraWGNjery9gffxl3bjPXZSHKrtg6kvK46StZI3yWxqfZ+Cq8VevS75Tk
zZ436krhcpW7Ndlqc+fkGdolIEY1otJw1IZo8OdzgydPeB/rMPt+9wNmKym+i4+0fTnuogfJd2qG
BpJiZY2WaAJ0nbZYDx2Rn9u1fv4loK//IDAdoCvyeEwBtFXoPdRSIFxz4qK8xmix3xQWWQCHS67x
4WmTQ9n/J2UgvFgZj8DbLD64pac7WY58hkTWOCEIezQkIqVW+wn17KTyO2G5rYWty7rHBKG9dLaf
ww9cVOUx22AjT86LDMgRGQC7qOcS04myk5ICz0uEY8Q+wRUnGiMgCmU+arPisNeCjnnb6bm1CpuO
2HE23Fgs4G8nPJz8kjMSLX2pyb/dawWJqP4WMUMS6rz0/tiDejodJImW1vEgW0Xq4qhzOKxsKDY6
WuFOj9i6EtUGPJW8ex2rvYQIxDhAwKPKIXfqTPRLsVVTkBD7kaZwIdugBAYX0GzGV8gIOxDeoCKv
jKjuhztlwbJnoX+RA/mfrQDWCbpLmsgWf4If98XC9G44/xMRqJojjKyAmvo1vUKF73rra5a+69uk
nu85RCQG5uaGyc6vukaHJkdlpvcPIPbvHszl3qr073QI30ON6w3+sBNK3cpNw2r63V/5n7fErnmX
TD3cGYMxIzPKkTzj6W297z6UuO7vq5EEZsm5L7csbhL4Js5407M/cgjTLuK9qVIYB/tK/0kEH4Pq
3HWAyYSWMhdjJGvxjSu0fE65VmpdpjEO+ZTJW7ilkntpD2rN5W6njA6haqZDHG0M81fdq9YhOHjb
qYid6eZSee5W+vwObU6eQIoS4uvhiBdo9R6x8XT7VuT4/4lTK4S3hw2ixGvYRTjXJzADgwzhIyTY
sVTtLt2sFqPbPy+clyBlnrRsqEqZDU+R/x33wThyoZV0IBHiQRxqadllXCHMBF5QPcMLJWlHGBlG
DGJKzvG4LpQx+N846NaQj88dVU+rPsDv8dtGsE6HbfB93xFdt4IcVpor9e3Tq6Ct4B3fNPybC5RT
xxz1iBptwF3sOOzaSUp05Zd9zD+F/r2IXDyYEKmGyGtXboSpHx2Oe+Zitn52tF77oSHa6FCHEz11
DYEO96+VPjbJL1m1rvjBKqxlP5dqXM7pDk1fChSyjJ1z5U/uT1gMMTHHqW5iNu9dXGjyR6+rFEID
B5Ng/qsYI37A2QY80Pfr9GGcPPoWgjgyKZnhrVSIIQqnq6dPTAGr5n/JGlRfLuTFXAVTdcPhOmlR
6biMeLReh3112yA+2kqehPmT4LA457tcPn0VJHaefWeu/wXV571MA/WZmOPYXJWcRqrYAcjKb1/z
8KreyuCJkSQ9SR8qydRDyj7N4cMnjVT4OU5Gs+VQBpE+ovy6uGCNpBsp5PbRb2YZu9TLuks/pPuo
h3P2vT8A0YwmUSH/ioe5QanrJviGPxLNNZ3yx2yIqin81BwUJ/4py59daMTNUiUf1NWSAqourea4
acvuWezYBh9TQGLkoVF9CHsw4CXOCtpoAak6w49PvaeHk1Yq7If0Pv5nAo/S6WKSdxZbG1vfoC1M
Dk52bWYbOHHmZEx3g81dHxVKW/dp+t6eW0CpdowcnevexJw0H7R+LBQDkflReJ6Jv6LMCijuLCds
3c18SztJ6HYGxyPEhJeQHPzPM7zwGTe6b4Ct1WhWXZVhhMf1yXdR0OaOHtiF4dCB7dBs0cu6xq5O
XlKCnnEcEyGRywFKMQ3xb3Bq6se0yGEPXV5rxT0IfezfROGCi9bySa70rTPXNjetv3tyvoWtpY4v
A032jSYeNEkl04xdeKiwT7B8LVchmbNuUS3jCJhn0KthFqTTrUqwcDOKcscUf4lHang5nzCpy/cR
D7mIoYMU1rsrCb07xoyua0TMXxHdI7pfouiJOpyuqS+SexrjadzvQ/4GYsJOCDtP6V2PZKgdWmxS
lUg4wu6A1EfQ3d3PQlv80e2hKFYXbGlnUQtG+NL8OZqYnzwaLgIRAvCZ6jzWoOeXJ+C5IQ+SizPc
d8Wz+RJqUorS6aTNmAuYDTMMEdPo7Y7jPY+KSROLJasTu+4eRDGHrXB1xkgwsszrgRU8LjZmuCUd
rBWCuZSOvrWzSqNdSF6g/OLxmm0e9o9vstvUS+BrVigfRCHNlZ6iO/GnnCSpCn1Ioh0C9bxWeW3Y
/QWj21qBHQjD4ZT4maShbuuLh0XcTxz5ziSrzjOADRaGXHnQA6zmCS0bURKoi9F+kyWN5/PtHOk2
UyBfvvEWCfF11VjBNVax+1nI3iDhUwcoh2JSTNBQkH/T99Op5ZxM8uiXW2viJqpf3APDFzPHhJU7
gmY03QfWkuVGfiSMNRkpHcpSHvMfe9nP0IaYncUQgqef/4TF3CtJJ7v2MAFlG213u2noPzOtPhH1
uurRuV8k4moh/Swaa+L3/cz6TC+O98+93tsGLzEF4HZ3uzpUlNEsI3HTMDzfKXmxy4EQdioMntvk
qukPTMWN7hHpV9xUUBTk/kxL77mlY4RIzR+/16NpWLxU4GfAVuaNwdgBD2Glj+snNh0SQqFFbO/z
XKQU0QLOW4QOb/VCUBLviB1BB55LalCWBlSEtMTsRj5mNA/APbOWI5F/gVA+dUbEbkDDZNM79Zi5
1+CbJV381NQhcwPUFkC3K3UKmp35+A/xgHEc6Z+pKJmlXO3y2JXr3nJlba3/+XSYtXVEmor8xyWH
v9ELBiFFiWliHI4tSpts+c+nGROKpfGeCdDuGTNsqqihNeKQqnIfwxwfnDMKPeyYPhBVZ72m/gfn
feXtVh4n/CaEObbojfxJOljgJ2p3c+DImSZpa6zahR0ZMqFWTaP8m15zs5ezT243jrhBNf3b/SVP
KCKvTzyQ1VFqBumuIT8vF+kudVPlEbt56YXoRoiakUAe/36zRerVBkdlkuR3+4L1KfLyXh3TNB6f
rEqmJFvsTT8IhFPrIs6tZanvesiii+ppD0LTms4fRzFeOfDdswh9ujJ0VBK8tXIQ5/qaoFlaRSTz
fBPe9s7qrigD0qRqBedBb1VYhWoBgz7r7Dp2gy9s7Ig3ard6WF7E6aEUt00LupxXxInLrQ1qZIAj
CfdeVhBk2D6UoR3+P2btzdN0cjL847FE6NmUV/UKieGI7K3dEd46fIfV2l++Nd6qEwYNAj+f7mw/
V1hE+CKDJBuMeNnuGjQuwHUls7F3588CgzaG8bHhwebx6jsfNsrPi6huCUWpGY4HNhKm4yg3J0q/
NhdnF8sLJolLKrzFG+sE06VLs4UG9rwPDr3qWt+1HkQRb9k5IpFdypoQ8gp0J3uGZL5gJG6bNT7C
lOWgwceFRFQRF+aFh6ECj0/Vq08PshBdhrayqUmK+/fCO1tZ4j64gh5zSy0dWgQm6Tx6ORMbGjp4
CvvJue/PsN0L0qPSAnjCdftj1UrVjcWlR7sdUXPtNIJk3nR/Gw4DBcOW3Qv9MjRwUDkrcq7oIPip
tzmk4sSdB3s8otwN2HI212FVPmRaX01v+8QfNVcHGqrxHthsI8bw1gPaeAUFg8yys0P2fdCE2tF+
K9D9tJ8vgCoGMBX83KOcQiCW15ukc6LzEEQbXAf8EqDnADR41+j7+IKVn+7JmYd4I2Fp4UTytElN
psSYZJmxC+99xMJtzzH0Ap+rPR+/5o9wxAvdDxnupsMSQy6Xbcq+t9nqZObjvCWWl98fJ6iTf/y9
A/9Qx9tcV2ekqb/YcgdPEHr1FZJ76Z64oUkHP4iYgmSZ/4lgKXpdYGRr9EXDGNAYMJGAekxn0XRv
VXQDBEFZayWp2j9EO7IierEJ29tVk/BimuJlP1nky0JFGqT3oGcRJYzIm7hKFjaJu6uJfVA7H/2r
Q/Tqu682CEUTNJrFyXoQ6c0/YqBshAnJm9tqLkcutT5UYpZIfras7IY60pjsmhqcBeIKBp5yQfZr
+6yAX3oIAF0yaWi49vLUAeeIqCKFJJ/fwSlPGAjAG4P4ZZG9fvAU68orN/j9iTWNszTiV1Rhodz9
C6iDWSzuwNHn5JPs48c+AGcz8eEfKk17vQEsGZKlP5/T6hLsr3xnAPN4quIGavQ6iGIiT6XOrevj
gfTO1DehPHKskh3/bKja4HFFF/aJnz/9tlUhyN6QxHAvnttl6PHf6a3y7r7suQzcVR0+lv30xhsN
lacWqiDzeCAre5jFRVkZYLKnUy3si6qVYki08Yew+CGvvyHO56wIaZ8stFGYeOJV07+q23p42MrL
r4FctI7S3CUCOhnpjslBdH9NV3cL4LvA1RrB67Znd1E+FQfEJ7BIy5gGZGVyO4VC8lLRm9AxyBfQ
krSEcHltScOOw3exJjKp7RhmAxx03i7/1as6ub0c+L0Ec4cVWRkgnXRmN4sm+dn0PIJdk96Z+f8N
evJe+SAeHBdqyVRQfN9qm7fo64T7aPT68FYfgnxIxK5fJuw2+rgDa5kn6DgraRiLes/4Sm30Gaoy
2mB1vpkZHTmW3SUbSJKqqED1sKWPMTAe8loU5waaRmG0yako0spHADJXRE7YsNPzghyrmLP+Qq6Y
vMKMso6TPU2eevgXrHPoamoZTftXG9bEOdkS1pPAPZ6IxOKVIOSC6wx93OKUC0EXjFfFNTBmFeNS
voPFxlkIlwhKQeWjHYzXNfO1QzSVKdG+D5aQXpWXpvjYnLEpEZoHnmH0P+zpkXAftXuqbUzqw4eU
R+UX7BRCXEJxDxhkdFEG8Qye9iesGgBUtigz+S+N057Uf/DXk/LqEv7qy34qxE8z01qdmnHnXmVA
AJBsTN3lThIFlTr5OlCkRvYFmbtA0SzDZMtjwAH3CIqLykjCcNDgJR1DETznYUbmOvAgrVrVAgdv
g6MimVkpq1Uz08/1zLu2zu0AGyMnQ31Ykr0GWA2gEH5oO3PxTgK7Edu5H+uGC8VxsT9zybToQysZ
doGyp+Wl3JRPbndI+6pyqBJmVvBvlUk0YbHaLTBB5OB0boHsAZD1dF2d+EJ8XSj3XUjOq6OhDEIy
L+nVVMn83ydRhjzt3i28Kbrm7sbeGIqFtdrqbuzl1IrItcoadaqcPNxr2I1pBlWrswnaBoghnDdj
p9v5ubSTXS1rNCXWm2jCOyer3Bae+u91TFdLqeYLJEW7QoJH7vTlnincAAfrw+uKty74e9s3S+AZ
hB2nGhV6OOAvHgwc/CTwLSyO+uzdijjA6yc0xMFpp7KPSkcQMAUjoxLl9t4Zkyt21PRfU5e8pTgY
klOo2y+cYFHZUSmqL3Cl5JzIzt5MdFlWYlAtRf++mLs3izIR0Za/b2ibIdB7XHHXr8WaS4dovZRx
gw9J6EJjI6sFWnjC3QjeEnJ7lPPTw6WmAhvpVU5BrTg/zGbsMtRJS4sgxw1bDHstzYBVnMCnoPJ9
xP/zYra48r43yxCMYk9eNu4XWdUElBesWETWVMVmAK8BhdznkvU2WucFjdqeRGDxcXN/Bt7gWl7m
qCPkoOv51ZL4tNbq0AdLFIaLg5eeSAGmej5ELUry5eC4tVDVUbGOLzpHnQpjpZQhsKwD/0LJDxe1
5WeHdl2Z8V2a0itzlOC4iNe4wZDxHzJ9J8VGWc5dKbQ0PPwNX1Y0dZR1DFCX27KTZ+X83dc7jH9T
qSHXL+J+SLasayh7hN3t0co69++1E0Tl3guNIpaCBNsb9Pe9PEOMDPwCyZATXBpK/sY6zLvQuntj
C6VmIAD6cbWR8KBWJA/TKyTKcV69KsLH/ggz+EdCXbZQHLIsDojwUgSK6oZ/Mt23tJTgLiEnaNBr
rpa8cNXlWldhkmyGvQ8Qg+BUfM7PNY7TEpn/75/jzS9/CdK4zUJ1RpCejbVth9U/EQfYCNPe/Rlm
cSItE4Ef5JjBx1NjiDB3dTOofyMG2VF48C9PvJ3ThfhsXGF0mhTaLc89LUZXsdgKpVMszJi7pRJC
RqOFa6nsbsWdTyaorr6yFMUeF4wnQb8hax7nIYmN1d13wUm/uieaQhS8yMLSQsSIIUKcDq7EuHwB
vonLWAsaVN9WcgcyiQgxSNH7xFPFIFuZtc2CBTzGToeL0Y0n6wMFl6gK0iFeEUmtP94sRSWMvahA
LtyuiiMrbjsR3mKizyc+FOopkFNCIHbKUY9DoD7kgl7s3gRQPpuoLG1ikBEWdj/y4WFyNsfWjH/w
3riukNIrgAYws3ZN4QIe7bbCrJ4XoPFLyphtE4X7d4g2UTkP6u2ypwUHvnhjAEwgK7Kn3GonzG54
NvKxXXVjaUpepreFz/om3HNJeTPZqpslKcfq/43ruIPJ19jmkOnvJEaLAaF1zxk4CRh+u89uMQ4r
7laltPGwXE0g2dqSijYK9uv9ytGS0jSNXAmyABy/s09Ge9lbm2Se2ItTocqN8Wn8Zo/r+tXSdNPi
dS+2DqmL1upXF8B/oAYksDwF+NMrtCEI5p6KTANTSMcSGcybtTSmIs6RaWnlV3F9DJqCvP0kGfUr
fkCvxPkZGa2UZmNNIabU8bNwHO68mkmF1FK6CObyO5IVhfdIJSJq3a/gFzU3nBoMtGxiXBDaUhbq
9yJnbqbCSy/kY1miySkLfXMU1tb8NKIloBqyrhPxlMrFxCkXICvPZmD2UmK1MsHnRwLJk4beLRHU
wrYF9BKrkyRrlQdlKHpgpp1Z6Z4lHFmu5MROT5FR0zWmqO7llDpppsnex8v22mnGk9jKm0Ozdv1U
2AwcA3idQLS5GmhzU5ELBVy3l6Anrdmz9vGBM0Anx6XHTKbbL/MIFB3Rehfl35Vp8kDbi6d3o9Ag
XdkIXUqoHQKgOIku0jK9cuV+wLqNoqu9Dvy6GaMTx00BViB2mch5SrTHFuqli42L+dq9y2WCcGta
s0AsgngJ5a7tVxZD+09tcs6+34gTWUOjpTRJ09lTSvqO78jVFd0Z5KyDBGnY3vmupfjkh0D8iYrA
Eu+BcSIVZHKC089xsuW7VEA6P2/QGYPbNd+kKJ3bXTvpYXtJHxhtfMXc35td04jLgFmy1UssRMeZ
uH+w9cHEYSw3bmoAkfxX5pa3x5oO8MDoNgPV62PZZpE2y1BODQXFUFXv+QutR1KrYTx7KvufBqEf
XAGHLCv75Qdv7cXH855PftldM4HpJzo3uU65jBnJwAcWE97SJ19FSvqJq+A1IQm4PqNnLi42jaXi
bJxKHLZW+UCMO6YdBGUdbdzidTG0ERJ/58vw71w9Jl3bUMeW4HHtJ6PgcpHIu03iYBwUZNgz7+3S
UBKgsWsSrjoGKS9XDKxgY1f/KrGZ+ozdLsv+O3IuWiK184P0f7Q9U/8YmKQgYHPT8Ioykjg+94La
MATFq7axgwLBpMDeUkYK/aftJm4nz+KOxr9okRxwrqL4QALOw9duQn+qsqy705MdKNw99D4Vzeoy
sRGyrs3LDgQxZswMq2P0NvKjaxTftU8IOPylQzoAWN3l/VI2QylIZsZLpVcKjGTlQtCoAv8k3PGp
cxXPN/FV1qAhGM9VgA2DlR+L0wxHQ6Dsd3ka2Uu5qDsQvC4gxgx44fUU9M2E2IlO8kMG1UTyDByu
O+lMTliXkKi2YmfjGHzoDMQthGjxwci7VQ/dt3m661qVIX/fil0/wiWeS0hXOWKKh5/OLS4So8M7
S56fheoqZ6UTG2xfO/y4nw9pSPnOatZDWxEFGdGhY1v6YW76u7VO3LljWSAyRdtiEHNvIyeqztcp
Ccavs6jF8Rs9lmsFvbK4hiYJXj4V1JeoELjqsyvFXqf61opOJ1ZxXrElb/Mgon+L/U9zz7gVbCcB
iPSYUESHPWQBkAEgtjS/KIVLvj+2kDx7ExtkJ2fbliHF0Vf1KJXIrRZpquRvEiTypKxH8l7NFQUt
pvum+cvQyKi3A0RPv2afvi3Em06YXzBadaZEUR//AJNYh7QpTR2f3uZa0gNf0/QeJ9lXfMOrqqrH
fiXRJf5bajAMRAEgTqhbovegZMySwWo3/rm4qkwh8r344+Jhzn/3pbbpkSsZ7SuCGXE1S8DKUTz0
nsY9brKRk/pV0uVUdvRunUdl5qtf3IV4A5qDtSh9h2GpsRzWauZV5oVCwGZvnXnUCb0v6jPnQ+mn
cuu87TN5F6e8VzxPyJ3NrixLTgZmkhr6w6xurR79D8xTK+ybUBMrYfNLWWCpzcDy+tikY6JmbslY
Q7iwXvIWnswD5QNEWCOxVKe9rugIN8DXC1U6BCfKyJQGWu9ObgGmgv5b9FU7uE6NDfU7xdbEfFjs
vt68lNtetLdgzGJALajUbVUHn0s9PMNELWnQWPb5CWIuIMtFlkIHRVsbJVilvTSjw/1q06e6KXyf
m10zqH7JLV9vKIyrgdQoGq6Vcyidsy3OSOTQ/u2XawuJSZjZNjVeyjL9AbLSgFAg0PLbx767VEPk
2Js7ePbRLgKQerHiCoRlc15R3OZDEv7hat+k16mxYLp4iX51hovPEyry2RRlTmKznR1spG6fzbtg
5y3ApwVEzrN4UGnt0UimP/u4URURt3BHC2pyXfAL4yV6MCy7wnmKU3b/0/v75I99rnDcqYmxiuDW
GkY3HfqDEK2CHBJpHN1VAfxvVyFaOqL1iBLQ01935DovTm1OyQmu6CZQn4U8hjBIUwoVE7rIjsKI
5qqYeicvfzJ5bnoNpxNtVuUNOstbE9zGYpj9tmg7I1h2OVq0M+68KS7VqrVILSDHGxdLMMqf+4+Z
htD0UgMpBn9ImJZgIvUQcmcThpM9L0uol8r+pk8x1KvHCz10ujgzSAYkT+S03zU39C+K3/H9bKKp
ZMQ15iFVkC2bBZswEADdwaq1SU/He05h/zHXbbtvLLTVF3ZM3uNwya/nIHKmfL5wLx6RwrfgwBRp
240X9J+iO4cJU4F+1/hyXN2zq7w+bAlK6CGDWFeQnA4mXr8Imm4Jyg9T1KHBKrhEk+ch+UBCBV+c
4x1ZyQXShGVrxvhz1kqRmnlmzdULL4ck31OzOAqVvlhFfbzFDWRHJZEZs/QMxfHys5jnEHQADJ/i
SkYasa9fR0JE6QB9og4uZW+6dnR9BbSIDdhYdnzwo/20nvaa04/b4FglcRaDgb28KD+CuIVe/Mky
ji2x+mrL+uGDzNY3oB7tqQ2nB0tqL/+85maIpO1Cysoam5RFAOYFkSCR+2ap+JzuxF6Ju4FYS8rE
TA8eZbLfkSmGhobE9/PD3OU/DZNgYuGxonV/DzHOERbHDkQUcCx9p+xrFNtfvyxA+kNkBvWk03Jq
UH3J6PCqwxvOpnM913TbvFRuZRK9cQx6px46woAQTL17aUnvMPpNtRECLRE8sMWhXoJkRjJvjb8T
Db9Fb7IHmNK6xshLxnF5VxpOGFGeAm1XU1oZwO/nZjOm/db5bwCOJ9mkAwhcBIBGeYXo3eEB8zgP
S93Sguegnm6Edqjg4lgIGQPe9odAlgps19Yj5LvJoCK8cZVRLczBXCA8jS2LUvGGKaG9X6g+zl5q
6ByKFw+rN8jjh5CVZx/f/x7AFG6whJ79hj0JkTqj1/hAkc2PcJOEkbYsaAsHrP34M/T7vFD30k+q
Kua7Yce+/MsoyzwkB5Sy016ETELt/J7EOzzFj9wrizoEc9Us9YjGTMh1fzWf3bTWHvgVX1QJoF02
WAK7ooOtBcbTukHdJ98pDaO7/0NbXs2xVbgiO6u5HUmElemu2HWMCeLz95EOLrxKiX+gUBJdZ3ki
E4SLapbXxzOalDLqLLbj6sVFpJBVxoLgrNcoeFGocGRHXOCIBORel77HRVqNQg0HmrAYnXfNFzoD
DyRyh8prQ+x8aFmIPENnctvae444p+hD+s5TZ+ZhrlEI5fJz2C4XAvOkcnA6AykkUrJA19oUuk1G
oHrAv0SeRkR8P7KnFiclbyDQLcfUYdwDXkdVvdxB1IDaNg+L6JSa0t9PEPpJ9J07IoHGXQK8wUOR
SgT/eVZABTksUDJ+sXIT6tWsxh8lsrzkWjwXhjZjnuHwhk6egSMYas+ZAKvBR+lcGvj77Eq4MhlH
8hmrd+A4JAzTMLPhF6cqlk+vaDqnzJ5ry6BdyH8D6L8Ao0W2vEWzs7JYxut7QjC6c/I7q6zxXPwo
kTtr/3/IkeLZoo2vcIe5USHLo3Yonlj+PmKcSJGIaex6HwqjsQ6t8vDi0+NEClhgoWruYxawE2dt
S34n0FwHZKFWY5mJj1coGhJIk3ZWWtp8xHQJcnoUt63CqJENBHSnjMlJlDNorFOO6G7/NJJoh9Vg
gWMqVoZamO/Oc6nJYW3pIWQotXIizMx/zAcPswmtaM2mvvbGOe496TSsPN8kXjJxYFZJ1ohlpxJo
gafz7NhCSMGxaJ88uy6YQ4YgMkl3xTTBHqSRuZTFojgnnkPO8PH4Ku0C2iOxoE6nVKV2uzktvtS/
CqRhyyXc4YkSCjxz5RIhynQ2fQdQn72z2Itx78t6uYS4+x9Vyv3x+LKL6ru3C/Bo9DMRq6VEjTSv
sLuER1FIwj4ugPjdpfp5lk6y8mgdkIOswJoW7eWLZK27QR07DcEmudW9HAqtP3yLjqgliruH0oNh
LdCxN/hw4/Hrv2/5br2/5dGL46rdIfghVyM0xyA4j3XgC9ajcr5U9q+UmI2bSIS9Q7h3s9IFITwB
6W3svjimhm0Z1VaqPAxfWrOrPQwhY22wmrqC59ggRjC4XDFilvOzT6Gg1b4Z38TcRcEaDhNje21r
sy69vep6IXVvKrVdQgEI0Bd9BEPCo+LgkNVhiCdbf26YpdBSPQEAOaLnfJzSQsEKTcviRK1tPzpL
YCzUZGoL27fxfkAWhB1fn4CxVQezPlT3c6EmfhPAKLS1rFE3ncZ5fJlyN1lgoekeIfEYt9ztWNOw
nAsQAMdTkWVIrgnWTPLLJmZQ+3cRrKnkXcdq9Itf4abmYHpEpghD66S0TYkgDs7DtRw9tPIPLYED
2XaP4G3Jvu8EcyNaw3kcCytCaf2UgZOeIU3epTh3zX2aAgbD6rDR9b1po5I5gj66ObCdzkvFey/X
FsEr1z1lU/IVwQkQgRbCWJCXbU32xJcODOdJjgYAnboK6J6/HIcTelqdiFhmJ5bwQRFBg1NQizGV
AlxUxnuCjCarTbJde0SinuBvz8L3YKieZwycc0PnnQ4fao0S3kked07VdzipcdTqOdAZgYw7IRy+
aAHDd9lFzQX2oPi0JLtJft90lr4tyudNqQyxFgF5cH5zL+Vv46zQz29uBI28ZOieSUK06dwL+agc
pqI/EHrnu3Jy1YOAL0JchaXBhdkOwh7LKKcSX6WWYD1SJLSXt+1bboAduLUfd8sPMfe8G06BHBl/
toMoCqOCS4DxZWcQeITIjb59ztOCoQ+pVFBp9LKa98UTXGI63JTVYrarM9CP2Cn4Ns4TFKf2nDR1
k0z8rCalK4kSzhCnV457gupM6gYZMRU30JoMlC3UXIX8KSsuN9VLy8Q5ULzylS2NZj+aC1NSrZGU
OewFeCeuSm1v7v+I730CdmJXBNYzGH8PTIJY92m62ecalDa94adUKcWFWSlgXWts6TJ3ip7fh1as
uJzeSAR++MNhRfBWVP3mAVYoYxyhX71mgpae3kO9qw7REeo9iWTIVQ4k/+I89v9Pc9BNMkNGONok
D6ib0d809FRZp7DFZvZDsQU8G5k+UtUiB6YfCsLy5lUp/4nzEfdb8G5V7AIPydkgTIRc4gdb54pk
cOToXIfkZqcwi2BYJSJbFm2me1nlu9EC82jtcCZmCZMa26avaylgIhH9CTvKnMWeg3b08SimQNtG
ILCk8t4N1X5ML6ZaWLGw3VceNmwWxPwvEHH1/jF+NrSHeLqyfKQjXMMM78iDw45TjoP3VMQGJCkr
DGMEtfhyKidJRt8fs2f3KuOcCmr+k/4hz9SsEDhPrSloYteS97zaw+FvErpYblLBLDVs45gG381A
6qFNHOgLAWfl+T10rejgqpVWQgrP1PVtXUhBPG1QJZg6j8vi3P8VHcfVbx6dkfO8vlzCQgTGg2ft
yL1z6dha2oKJqR68JmVDbbsRUJaHBKDaKrGprhLwwFEF5IzocKTPQS+6FjbX6PYNxqXOZeqMzJjr
tC9yO8w6WBLFStH5XLKyUK2/Moc+iO9/fCaF1SBh9crMzk2VpapE5kJsjfZuLVvx+/f2E6xeT7MY
nHZykNM44pX84q8ICs2+gNNutm7hdPhyJfNE+X3whiQRJ+QnCEnzqjk3gkfWbgUzXMjBHZrOrhzx
Np+pD1kX/KAXZxfOgPC+8yBXL8BfZ3XgVdneT0LMa9L7b/jwY9pTdXARKTvbTF0ErnZ0hh4y07Ft
W9gBtN03Z1OcJexXTRdasuC9CiPAGyG+NhfRxj8HLM/0J0xEbZ96VeO0vVOm9xpx58PrGJ5bBxmb
2ZZbdiCZ0/7PP8AwOfqs3aYEr2yYmTmqIKzosOJ/xSPHKnRS/bxjr0nsFTQ5qXHsPRFTMnKBTMqd
cwWPrZNqnqmmVdfknZMFy4ltbyBG/cE/0teCw2zXz+0j8EdUqsE3YlqTBFPNJtRiLL7uxi3oYKFj
5eB+MKrc/PF85xjOX/OTFmDO8pN9BRGXz7LS+e8UwbA18gRP3LR8BY2dbiCRrXNaRl2crN/rQvjN
yD6tHJ1hO+ijkRY6+b3r/BsjGJSypnpMOMd44wnDEQufHzd/eFG4gIwqZ0ToKDXZL6PdguIaWa2Q
A2OEYih3y7MVMfbVpjrCcgYcQkVR5uwNrKRs3Xvu9mOWJRKwMkXI1oEphleRWFaNCgl9Ge9MJjtK
MnMxGjC13/L4wmBcxCRmTTI+Y/TM+Rtjczo29MflboBCUGPBQyTFRlbuAKfJ3InBDm+a3tLznvKK
It5mU8ep1+ehXHL4IEVjqcCQ+tTHR+qfmMIeaqzX0nlD3/bv6Ut/nlPWFzocEYtneqp6lBF8qtyg
ZRjaRtMoyPyASAUDa6Yv0gypqXMDpCrpsR3nsJU8vx3Eq9yhAAejSfxg8VQiSq9rVdHW7NhqOI+s
Q+ezstg2Q2yL40FnwRh6GZ1g1OOghti07rGRLyFrxaXwDd+43E07T+iFmpcM1Y1Ug+So+uwZMhiA
AWJyf3j5i6St132XgbliSqBxSQeUAWGHW/6ZcrioTxDbE6xs8L1aldxK1m6bvh+wOldvk0m/oW/e
/zYmiLRGIRxKfdtS52MinjQ4Np9oamwphkTHETi+23ul4vRhAH4n0Cb5oMVXyu5JTMCgeVr78ukm
9pvKgve8cQOrtk23JsZm4KRXrd8dg460PRk4r0aYJmSdR1pzUZr5GLtGcgozgzMCIGeb5LzpU0NE
29VJ7YOKy16tts+PcKLwhtEKg7KMuMcc8z4eV4iwmc0fiE/mF3YmM9qy7LuFAunfUG0WAa5vlPe2
QnPCwyAEfOun0yZAdjL17l+ADIcqW49Xk74QoVi3/NTKaCkOyuINh1k13ZoGXcvptDxROaHA0DW8
Tn0pVB9WIy9Qi/vIA54iDgFK8+TVFnEmHRBfwjG36UeDL4mzBEe2I93xnFDN1SL6tO0HSWgeSJ/g
IOuC+YuaAe/NQxZ5O1uXdzrydeQrQeY4sc0eJMoOF6xzBeRmaP+AYevA58/4q/pnmgeZTzSXofhd
DHwPSIps6AZSraRiUdaFuynO8fjB5MxTy8zXtDXN6Jm4KUHEbT5xYRfFb1zoAEK8nFN1QU0Pk2cj
b38SmevJhdmW0Ipv2DMa1XzKhQOPEJjzFbtRqDY+sotTXNSyVD+oMXf+RBM65HRu6zW/3P5IGoWH
kUr392R5aEfuNi4s8M2lmKQ1Oi2Sv3YKbmzAdpKrMkH6OhcEsvjoFJ0QWE+hnSHCK9UfZqP1twS9
6lX6CQinSvX1+1IP3/UGW9B57qdM7qLa1eawAJQBDu+esubRtZ2bYPIqVrAFxEpa0mr2+Ht/RB+a
2ySUIbv4lTT8D8627Navbrj8ZaSKltTGRQB8pfRnbWWowZRUG9L5tiMQuZaSCrpi4TaAKmixIY6f
Sp9D6o4SR9Wa4qMpeqPrYO/+3BB/ovx3+KDzcrMmMEBoOGjHGUqzhWbL1svZqf/y1nL14btHnKJg
YfORzKqWoTV/IBocvfyDfwgo2GiRxSHpXxiK0Mxq/x+L4GwASuLTlUIALsI4H2yylgy2O6hCMCSo
X4qFUi7KajDfdBFnAXSFp3XxGohBaOnROwWlJDumbAFZCMWU714dXlIk2MaiDlYMuwkxgIFwfuj5
8/r6Sc2pDM1bE9ksP/+2pwK0teM9ogfTVWOqPVaLo9MewKVV1Mrm28B6+qr4iLG30gjDaMslaGS2
nchFXtoLif6TU4yWuwBeVlOOyicKwDrhFHsMx2zJ1Lx4aggelRHGVpz9Kj8qV/hDl9r8QH9wOABr
dJXHENKFjhMwwem1K3cwpGjQDBGto7XjL/UrcNl1apMIKUVPkITf0VBgJhpZFe5F3glVgNiVFB4Z
GWuwKfrmFyR2NMsuEaqVY8JLofzMXUVt0p5pBgMNReWoq5hyIDYO0b8gOZthXLs7UD3n0kRNKZw2
conbvryb3a4zdl51szqYTZqLlaaCtgGDzQd8LTfiLutu//pafejY9KBkadpv/eK4PsU/rRxZIfjG
iAlrFWI75iZgz0yNX7Vpjp3tBmej2dyM0lxuGcTxOSpJ7IJGa907vLHEnIHHYbZrCcUUl7mlUa8S
0jMJNHVM7YWFPl90CeBqVzMEGYwTZVg/3I74j/Ei+zCZ62uciYFxrT7jf9+3c1cPZTLCGTAdjt0T
OGRvtx+4QxloBfo5EZba5WzuXI4J/JxLjKvQIeVSq9Le7l6xwmQ3CCZTqjyVjbpl1nytFo9ncMip
YljdZ96wzZsOTKM/KA9+nayFSvmWl8LIe8erg68/+3qGmU0aoAwO63uCdcUBQAvZEejPT5mV2c+c
SrqwlV0vMkv5OKo6Om6YwBIj1fhwM2xPJ20Zcb359+0hJihQyx19kgiJS7bRsWC5VNitw8h/vCtW
EsWo5umofruHzUuozXxLXn7eZQ0TnmLCgZ7Os9f6eii/a+sCSR+x5iULeTu1Yy1x6VhRVgRrVWsb
/PXJr1HexBevAqycu9TkcPpzmlQ+bTXLvND3RuNrIQmN66kDyeKS/j8KBZEFPIub32qhnWvVedl+
WHqtuEzvKf+puSxilrRYB/ndh36Xm7yFldKNj2zoVWXU9WrGA5WIMmOsSw9oV+huKA6lgLDT+KgA
rE0exGJRQX3SWMCwvFYwZ6Tph44lMsnXmg78PGQuFdjmVXOpxC1kI4TKwQmRA8A9SKbaJxFeJWpu
9bHiMQfzsCAcBR19QNLdAWr0Brdn4D9isNbNXBlzM56feQlk1Xom5+HNhngPr34Vyp34ZgGJ+MPA
LFNoe0pH7d4/3MPBJ6WgcXSCuh/c+7pO6zCghiMFsWJ/ucRpzuD0KqBolhZwjV0iMN1X/v7KUK/Z
Qyjk+NVgAes2F3ukK2VKS/hJIpgyh92jVtDttslUn0o1NGVGh58u0vXwn5R4+wojSErn1wkqxCKd
tw+31UZhNyzCZ4cE5fGohgfgjYMvOLDBwdbEeLR3hpaojovh5h4hJxrbyIF0Yhb93BFhszsMoDDK
2B1HiDNPlb2jziWVdc2QkRAn116n+CwAjY5Pt0VxZu3nkAVuW0ylFGY9DY27S8+hPU/Yx7aAmHPh
Jg+BAEQGCbAWQb9D9nRpD1h1gprq6eafchqBBTlDC1wYHN/+EfRw8xkr/B4gSStr1/XYeAkMIHjo
53SEH7GRxg0i1asC6Z/SocLVSgTvGsTRKkWCXGBw3zQtV2QRD0UshEcTNVLIr1W2R7EbsJI+LxiX
8FCrCeRaFd80KB2jipo4YNgc3ErhX2qnZj0C/2mzNsyVJEkF+e/pofc3rMjScwL9cSVE3HVFspX5
sO/v29bfU6QaWrXPMrMXBTqtvCmaYtO7Mhg6dwXBQrgPYrLDrsAUCv6RpTRcGsp4IoOaAH6N7ERm
b4khwQh9FAyDlYCl6m9A/AMOsuVTqonTgbCRToFAXGOEEnZnMrMC2QjV6rv/rgXa2i6iKJsgRauU
8xCzA61Vvytq0MlYCFsX3BnMy6VXhxvGG1MVg/S5RjHn7h0Xr6mlkDLkfed/UbuILgtbUZyKlwxL
QgJM0UC6DBvXLscO0yHSvZcD378StIgRWF5krHA964vWj458nDzh95fKMm6nTWvla1TKcWvrnEWn
JSNbiHzIDmbPUWrjl7dJGInnataB1/XJ0NgLnchEFKUiTfRsGtNTHx/D8zAGxGTifx73ejC+b5xF
QnOjIw9V43KtVin/7ByNSt+pLnlgcHJcDFnjCltXeZxN22ah1seE15EnmF/HX6eOFJfs8fi0OCKp
YFCqRayc5scmiqbnAvubResVn65r0eoKattSn6817kqhvYiYfl7aMepFMqlIN/NAEMU6NVvS3WKX
bSmRP+sOe31ntX5EKysy5IIXp/acBBOM6aoUyyU7zq9BYPxiRE4txbzJQYnqSfIoSWTgrp/rVWlK
IPmZT697yJKI4H6E1ehrDWtQk6W1ivnqJhAcOws91TdCAAe5MslxBZgOA87rRpmPrbKQTCZwvW8A
rO1fNw5V3OG/Cz1TfoVxXh1NM89Hx1cyRfvxpUva1Ziigf+bI52z1oWphLnsy8XvbK0YzYT3g399
GGKpNXTW1W+pVgjSwPGDiXtT6eRvH8aUcOMeftadxy4qf8Ok+yVeEIDo0iENSXR3fe3YNbwxA+Xn
R4qKZ5Evdt4Sn1cmMH5SvABrjeDddz18yxpCNES5P2zp56CyEUXzFbL21AfGdRqKN5aqrFBj3JNc
kpd3yM37eI0ZNWHgLIuWNRYnbO6DNjQrbf8yGhH/+rgW3DlVXIwLk3uUoqfixK9h8s8Gz/QA6i25
R2creFcAwZWa368JVpxszrbIoZIqdiQx7EqJ0E2j8Cq2a1LPbrkwA7psh1+/luDBxqWpb9dYkkVB
rhgloNLbW0PQM+BsX4w7m8QGTJbsZwNLFSgpQ1Hfvnw+hzcCLM+7dyxu/OshCo1NaU9NMwckogdJ
4gO0KlQ/rqZzOXg7OW9QnD5PgH3ugcpXRrxvEdDBoe+Ej8F/FoNEH6ZNz7ZY/L8OMufo2SdzUkaX
WbKR18R3YGiYl9NKG0lma98HUTukFNdYv6LxwH80HlX3ttbmXT/GxdPdtc4kTvgDBwmZMjSkyCe4
ILutwY3Ilr+S2NvNJa8rRe9XLx8ebH7B+NXSTkzDupqgJwpWQ3+0XvOHl+p59QeHMmuTeKUHyD1c
q7H2XnE4Q4nmIk3yZIbsoJieTsGSHFheSjGgOn1mxZIJfWmae9yEOQ8ecmh1lnUTmboeFTtnzAln
ZvLOhwQPhyxodUCjaXVHWSpTbNY0f9Qw3eFVKG47xXXa1n085DwTJtE6wdxL5oWAWYv3n5X5RUMG
odbJO89DIQD11nlitsph4R5sUFBBQOXnktb3vwS8Uaz7uUn4xz4PV5C7IoRZUHDA9LzeFaxj/Pe5
/+8XxZpLUptxYI3JWwbAahNovgMM0gOstWaKgOQME7Ze2I4qWFfTC8drGO3QrBM8edo9e/uX7FXR
qkwcbwo0QexrIWQIBJRPgx8XEIuMgq0jXDpHau59eFaE86zjXZslaLq+Pz1Ot/toyapsdJpNouCP
fqWJ0DnHgbTS5By3DIf54rtNWgWXv1J/OftaJqCeGZWxPRdi92QBtyKj+GhzOhjLvJox8aK3T1Jx
OH0D+quVO1gR8NH28sLnajCwpkQiUCl+jZiFsO+x9YbJ5HeGyNKerdNRFIW8tPtR9unp9g4g0t6O
ZdW1tlGfHvtfJqSMbT7cJqcQRy7kes8+4uj0Un8zxuArBy56a4FmE6qSCvy1ULGkJJ6GmFzP5y08
fGIIYQvK/o7jH1RuxDzyxyf2g69VXoYE8+N1LHbZ6NeCZMXJe/V5/RopzYJNgjgShjYbz3o/ZqLc
tFT+uLgKoyyOPahzOmNeftFgVuH2yAJNEi6WTLrcu+1t+Cq3XbbcWX05bFU88bdyqjP8w+iVpd/F
mXuVOD4Pm9TFm28mSFkgXlUoMcbMo7k8b0YUrX6tKZpC0FbIZMwqUyQZvUQULgP2aYbYc1wktPGr
v5UAe1HRZq9Qb/22vp2boONI185amHfZnLdhZzCKDUed/7gqj8n8o2NLh9piPWikfRixcF2li2R0
1cn93wocOv6t7tS57t0l2NpBgYkCRbC2EGiZ/6UQCLq9Lkc4dS75dA3xOoZEAE7SD4+urBiiXYAX
93KLb4BzJACF4SyiLWBDszsnBnJTAUO1kiovkPJm14AqxpA6k0OyDeZdMQ/ii5wiJ5gcGNTd1SCg
YhPlQOTwTqHyd7YrcyRf4AaadcLvvigm6sA6TOH4kI4sfp/XyRCbn39OBHvL0jriGzf6TDDVb2tz
yFYG1NTwRCLyXn5u6ZsXl6zB3bajokQ6nUlf/ZicRUG1i/iLz5DiSPCgf61OdnXNtpCTjjVi41qr
cJnRUCyCg8NIxQN/+awow2gIJyfgJanHJUYkvzwdzuB0zboGRkv5nF/2KAEGkSNc8GdpNCEAqIdt
V32HKtQNS1UgSjvTB+Gy7da/jczM0Ag40S8yG1wBBcEVKnSBEgLWgg8IobYid/JVbIVylsS+mlle
A1ca+yhdWZMl9vvGqCxN8AqE3CsKOX8cHi+7M6L2p1GTS1WAaC1oMg4GQWEWacNyQIyU2Oiga1WU
7yurp4Gd1/sM59Kk5LonOxf0n7ZfKLKGdfGBUseI2ph/m2+rlhhPoiUXefyY8EQ3ZgEHRTL1zger
mC+pQdgnoY0JtSMOSFqvhwDic2V17/ox7f+l7ov7j8CmpLjpWZlK4kXde6uce6KDUdlw33iLLIoa
3EmE88m7EYdKRD0rwqVUvrR2EhJy9uM/fB/wmmEfDhu3gmI1bw/hoMjxLP0Cjxhy0cH6yWKJVVaG
UlOaz2nCY9lsLf0W8N2hThF1RkvOxsNnrjVJfcaRRHJGBjY+QwFHo3FmXcPVJNJC5DurLtLq/8Wz
Clogeuz95Kz8Wf5QjzfPxkt7C0CAIMZfeHv+NV3BIi99h5PwuSekyNg46/jPpqHC5aA8ypcU64aZ
7YyNvJYPxDxEqAKJErfNattzPk10mOdOiw2tNiBJfRKRmnZFNnLhlf/kEgy/1g1jm2k5Wgg/aeK4
LDSvxV0lMuXR8sZ39bPA9dMA+KfBTzk5bOHBAzQNWeHPdcp+vZoX6NnbV4itfbeFJBx4V+TpHOwP
fayza6PyeAVEG654OhehSbqQSjHVXVtRgttEyXDR3BSxECUM6lgfzfCw6xclbjnyhvJZ6af6H8s6
/D5ON2QMCPjB+5hF5cBmXlf+VXO2alrBXYS2bLyZz1hTrUPsWX8Zm4uUEob4VRpTsZ+AItxpXjaI
xxcHj5/1nRRanbHazFMUyZalKC6662nOngEsaVeqK2Jpfoh9payhGTNV/mNlOijLHHlEPbG18rSx
nYDG3+NnObErjeX2JDWZn26xEB06kOCxYhX35mno9u3xE4OTnc8tvU04lfQscxN1MB66wPtaDQ3B
q01cbaXHkP7SDHL16QBGtvZTJQo+iRcmGLThAhSS7pqE/L6mkBinxy7qmpmkX5IfP34Niad09IZb
WGpH5xf4qWq/B4WWR9JEGXwBxj2QhVMRnNL5PlX12YaqMuYU7WFB3gndxQRXsVqo/+IFiESbyqIr
+4uXQzcQ0o4XGIql2sXOsP9KqKMhBBoVBFaWNTPbqUcF49RN6tQvhuSMtMKLgjehgFAAOGNuVd7M
7LikyLcfZgpp2IKAStsTtLWioXysaqNo0WdAJ+nwJNafgZZ+g8u1r8GXHv4asigwX0fzte7CCgt0
Pc9pzpIEkP+F4qICvhh0l3So38JFuPKlhhoaBG27/jNSQrc9aSWEoatIJRDGUzUjHHcqI34hpdzW
TZMHVCa/92reSbWHY1DCMaRMEo/OHkCvevbpyA/IL7bVgUB7cMcAr/JJP16pJV6jU92f9xqwZGEu
WkdKbgbcTf2C14dXKSFNgqo5aWWyuyIyRGIPF9YVOMbHhnQGzpdI9VgW9RxxpUwXsDAp4K8yS0F8
atDk6sqV5ycgw89dmG0vmwHv33Bx7fOx3/ExjrVLqY6H49g7cZ8YJoIXKc8/2x7FoWpD7XjkwlzB
QA47iZLA6WBIMkQbCyvdLX3DhKvvNxrxFjuFFRcOhC4ymR+KRipElrf2G5GNpxRKCKHXR/aRpBgG
7ZjzfAc3tlLsAKVgce2IM7CYCyIhGaDARxJ71NlcH3xue4t4d3jmGOw3EDfwdJ4pbbJoQCFs9xKV
r0YDauak/qFppD1idUJnYjR+ue2dxfLNCOq+MZDlIcGSCXmWhe5XTUEx9WeVU0fD9aEAzGnMbcrB
lWf2CQ5KcCN6+7qBQ/jdUxrqpuSDVIVZdAduaE0dd9L304q2J8xH8jTckF12zuHpv/w6sLeYGLmZ
LBIdjlqln70Yk5vSp9cBeN3hezfPEQHFSIqwKc7UcC8WdMmGRsTD5yGELmWg4LzHE1d0kLq9QIB7
CmUJVzsdXYZBxJbxn9319zxiDBM6B7cyCRlntqddyw7a0i7HpVKELv2BE7QDLYoyMur+HIIDD4HZ
+Sq1bdLjdsCa/jQrURNBUqtpkDK5JLMgqJj7/3UlWXEsP/3G7pwdnO33YxnmWyUJLlns/y9vjB+Q
rxgWOypxWNEZC1iRDvm9CoM+M9mSssKgQTHvqImUbT+r/d5bdu8aHoWEo+egiVKohpgQWkhSOvCL
OehrzhMliVvqaKpjzmrpgvU69N19gwXbXx/QiTnkKp90OAY7WnT73PMCssJ/LB3t0LqebWcYyqZm
Xs7zGW3LCu9Weh+buqtodZV3jYdBN5q+Ovrkcn6wvUWyDanVJ11qnynoGuRB+WrxD1FkKaDkWJHQ
FJc0vsh+FhJH79aRfWEzNjtCzwXfknXFdb7plLI9J5omtecg9wvs+1cvkkxsMJUzqH5eSvwFUyKt
3yvhJPESn2Cdf8BByYxRU74U7vHYT20o7iEvGPXu9kkiJhW/4uV65fo22weMNEBWQZ0s0T17YdJN
iBZdu/YRbtyVkn1ZMtTmJRWgNGzTVs6ecBe/793F25lbfTC8jdKDBpmWB+ezdfRjJrEW/Fn5uCpO
PS6hqv8lUhZB4ZQoVajAGvSFYWqvAHbEPugHCjrNThUuXR1G0gK6MOcwxaSjoSHW6TAuVwOY+uFC
YrCFqAxXaYGhOKGAcy9jzNQseWmvE7yjaeM229PIwFSLdJrXO9FVlvygk+7UF3+5gh8zVOQp9vmi
EtgeMkPE6OCadCjuOYHi6JMhlmZL0POImowLLtrRBXEPQBKDSoL6+YfEZCzZqAW5q8acpFPPJsG4
A6OO34QO62Ddzue9ZyzAtQUwWDvlnqjpf627h3c6SLHtZWURGTb3vCl0xjA5CP4mO118jIqz7gFN
pQwrX3epZZPuNFbt5GfH1VMruE7DWcfkXiQJIqp/eCYGoHQKPY9E1BfTCVpxJxtZXNY6kcJZdAbi
aUri3bFAcqXxW/4LmpfXnLEYq6P+jpZEPLXWDslkeYcj3qBwCzOUbF5AQi/3tEjrZrwb9fTLlsXO
wKVpDl4ob82lDBqhk/dj6AeMEYTurPqY4SVlIKFv9YXNyTui/aRgRLdmsVMhUndWL7URZFIojCfa
eWpalCuYbLpTwmzEp3TGt7VCGgOAlr66S2wy7CVwlNroEc4IEOkZKHG7h5yun+DrIGKvhRM21IIF
WLckeX/pobuRmmrWDpJOFFAordwpud+Rn9yOXKsWcz8n336go118eQM8h1LAKdyRt2httYB99KJv
OfpNShXOgi7R/0yegSNPuo1x76m21HU8rUYIQeG6vxdLEhChYWDMGZg7r7dVdoy0D3BT4/rWAASe
nXWe/CvloX/aQdudXuEPSTKcl395EaRI/kDMtq/j0TAT+GJGQqzQQlxZnSU9nmPbtkTRwZ2UtoF+
0QOEOpHkUHR/Q6zBNBXk+VjkaDK7klBbu8hqNboU7wmcVS5yY/AxmHuHZU8OV8wI0CGbNY9pqeJX
xbEm6yqDQmy97TBjj95RKKb4qmbiNqvqLO1YmoVLQ0BudP4DLBofqdXMyUvBVteoPBACMDJDWEiQ
8f5z9nC2Z2LJMR6nQCvgAbAiIukArK8tj/6OdE7lb4ZLKPvd0JDjn/vgVAJ1BBb1euau+Jx7ylvt
BIOJEJbDzMtWjKBcB8pyoxX7OY81eGDCQxY6Dr3dG69nAqMJR2Q0VY2PG0MNSMMI+qgSQI6m/yzD
ixMv8UuBFw9xunHHScbthKcinKIKU7jyIf0xevfsgenyS0rjjDJcfRYQiWcavbEZYoTqe7GnXOiE
ZFxOiD4sP0ISTe29NsClRr6zEybGe9YVlSverPCGe+AFEqW595T967godz4xX/O4oPc3F2ZUkaWW
XhKMxta8oXSKAT1dJRUfRT7z74cY2pz5t7IcYtje8WLlVBNitU00a58wZ2zPdmDocdYMMPZGBoop
o94zn7cQ6ldBKOkb4OmfTykYhg+SUno2iSbuJjXqDKBOPi7rLs81D/Bv/F3cUIokLNhIgOwSklaK
JfX0XagUf3e1DITCbLgyBQK5mnekFfGnhtcG+I4nEOmY/9xmbXakQIIi9RvrQrSHU4mJ6NIM0XBE
zKWm4HvxyjuGdAam1dFRPAH+iDL78JgjEPaxDNvWuvQ9cI+vlrOZeqdwjdkCX2RV9YayOau0bRpv
9kmiUtikZoAZn3yLJlJ+kcVjftHnA1WTejFsGzZkZ1YU1R3jIbDMfdgY94PY4rdwSh+2hpHQUIu8
nXiHcCJ1TFSUTH7AsNcZbVOA1oJ3+OMFJbLb8KrYjyXAI+luhHyGbTickwLipcNgMQDpgHSL0slE
qFFhr5YS3RL5kNFBmhDRDT4VK+ygL51b8eXPCMFqZ1ePxvwtle0QO2PbTj3H9fHBWQCQO/0hEEYN
NRsTuHtQv81fwASh7qQCq1wPzCcLAiKHtlL2SqRH94RvJ4aZMFg+w5WhsY6um0jUW7kCF3hL8jru
Dn3Pm+IG8L/Tq6AZXTeqBaJbbsF/IEkNKDCgugUdJ46bKSmEoMQ3RYu6NY6bPhFHz9DsV6G7Ijo+
2p5S4zCS5L06e9W7uYgf3QGASJtmEIR5mQ+H2rWwQiu4sl9/oRVgWEMcWyRuF/z7PKLZCfRQRske
30fdCQtcPYveHp/AQGl9Ud9mto9AjVMWcGA422r+fFiwqcdKlD7KhSANeHFnj7vBP9BFaEHVpOoL
gkv8ghK/PoJXSKURoJy/OQODLACB6oozXZ2bHTEL0IWy41LMYw0yUMhJB1zmYMsP+3S3OdEI40L4
1AJlxQbFiI5TTZDfCKRs+SCCg/nuy2QvcV5fxHcrGKstfqXV+yxzzFAoRvnwVg/vS3/rJl9kOjOb
OI/8MaaF9Y5HyrbeSPUxC8wICCvCBygXniHkqri9OIN7+vBmdPQCq73Xa4rDqWzjjVNmGFBIjb8r
n5Phy0Tf3FvaYBoYgx3loe6xNMpGgQhqDBASFdxEIUQwYUZ0QL56Kdu+O15/yQv/QWd5WiGObL/U
mFzdiT2we/OHunkjkzsDkJemiIowI6zjKHK+5ovoiEf5mn2W2vbBl8AQs/hXl2ipgj8JmQVpxpDq
tRDG3XnTR7K+kOTFIDEhOXxQiG/WFm2BXDdJcpTIswtTzSVeKaBCZxE05CQaOFZZHBfn3NqFX+j0
+9r3Z14V9w2Gg0Ua2vU+YWFt7RW8TviNkkU1bD9i5gyoLiWxOGfb/HlgxoqzXv0eo4zbcUpZP220
M+Vv0I3HApYmNxy6ra6x+qXgJwVa4gPKE6Juv+TcDgrrqO9wta59qZgYQRKMhcWkBu8dDbpFHzwR
SyldQSSV+9kTkIRr5apScmG/Nm9xROHu08y/Eg1gu0HTi7oAbgy0JjXggk1xSYlUI+54eGeWuN9h
UwjaIGgJCLmv72DAmxeJXimxp2iUKxoLCbWkSgbOyaz3RL5MdlUJpkyqn7W0/KcukYYxBvi1UFPH
T6pSrE79MXJL0A3E/0nLHql3Frg/2UOrptHXTkshpm6puKBSo7YIuyjX5J2HMm/zFCO+GTxnL7ig
rJ7pa3ONLwPCiKUb+Ee2RH5wcWUTIlL8XhW5pDnqDqajtpdXIf+dU5QoM0RJIm9CnR2X+e0l3G0T
5zbyx5X99z265NzJB/m30Cj17/DZ9KCYFNsm2Ng11tN4CcwxXqrdCFSszrrnUvPjF6KxcnahHubd
VSc94rDLRW0gAK/k61BmHVfXQDaeIjp2AsvxBFz2tyCKLfOBW1D+Ik7bS1QvXbu6HsyHK5T5xOhd
jMPgtB5UOUXdVxaYz8vdApopQ7zvDaahcwi43Sq6fHNERZ80S0vMYWf9l0n8BdkqPISowdJV5z+M
Y/v2qtfFqNonQ2+o6ML20233IFKRhTUCLn1GKu/DKuR2V1FqCpTFlH/wprJAssRl5zMZNKc0GVKG
6XUL5Ao5bweD07Cls30S0oQXQPwanQwrabXpRrndcbmneODycjwz/paIcvU8ZObYZGu8raeAk10b
UmPU0TpKe5suEc+Q4zc/3WTGUcAXJWeoSXfu51XiF3t9HfClH5Xu4T6y4j/c2Fu5HEb//QJ3XIsW
3FVOrONNwtV5orrOhzqfJ6VjUIWYSxmFxHRlGGEopsAFgRHkD/L7sM+nRUYJyj1Cr69i7OJOq192
nND5MW2oBn4qOgXWQe4EbA6FiBE19u5riUirFl02mkroB+3UytZ+xhS73MsL2Ck6x9s5ozQ+Lla4
dBwC49Vm6gt1BBrZobdJM1MrVQbdr7OAWmb2XcRQkgmAM1oELLPm7LNQnsM9/rgnyHr7TNXmgJmY
BCJyZiEuyEBXzzrsiXuKNxDp6BszHhuZQoCX0BVpKbBLuHsJVYAl4WpzkkN6SLSqpwNczgaNh6Vp
1l6TEnAqt+T5bv1xLTleGa3e6kqSz8zNpU9zYpfv0sFw7CGfTlvpRGBgiqB8sLa2RJ97RDPY8ZaW
PMbt65F2woAP8W7OzT7dugvJt2XZayNCv5OEfNx9ra5ibnVg3/zsfzuArlyfjitu5ilGx/2SGnMa
G7ZJwIZ5jhKY2EBv3geNqqlVE6ILgcHP8Oc3bxUI1hfXYPqrKZ6UUhQNU5LiOvYtd5zZPNnX2BXf
AVlTgVpbAVrul9ExVbyutPdjTt/MnPUkP/pSq3CYAR2NbXMYn+TwuSGcauEcsZY82BLOlhk1B+mO
gJwknboa8aDscLr30+JI2aGq0ip0ykmMtIb4nYNRhw2Mr7n/jkXCu14E1bC2Wi6/nrMwUZkD1/ts
eg5dyeAElZ2RbmxLnWBGHc45EOlzqiZGvlN8Guggua7iAfLpExX1YVSBmAHoVfayEeJUdyDF89tg
ClUwUrKrCzESCkQ/3EC18IpVEoDNLQ4HWWpk1FGUk6/G6I39khn+A1A1QjpMkdg+5n981xgQPUbj
Qnsd+53x986OzlxUPIB7/bRO9jPZFi2A49axjRl/tE8Ko5LkUkY+D53t16BOj4FTBXA4rSwd9Dbn
osJAR1j9kqP5AjA2ikLxAhQA9cDeUiyVnld/8EdSZi6wHUvRF6fTGxbpeeeZarDbNRE2Ed88+zEV
4BDTloFk/nE56yHk0bbeWLXqxIg5ge0MaZUl5B/fZh9ehpGhiDWT4gGc5NN1f1Gr88R6MowTab0+
pbX4EPJ64mGHI8hcRBkYgTvl0mkJQjViGwfApzAWqV6cFwR84YTzWLHW+oeHJPDYCh4MHl+Wd7ck
bWkONhFfcy5Hpk/Fayda6uz9kxGOhJSAyj5lMloVXnsVmUzyInRRpwQ5wTXR7cQSjndqrOyItogN
KeCHu02YXJLCOLO9NixyUtnIg0wxEQOjMUrGIuIH/bZ/5zIm++xyNNGg6nxIjqOfQU4JH2xUX+rh
LqmkHJv4FWEYWTy2yGGHDIaFfZbErAkxD+A/9F6qbtTr6/fZvwvPEE94lyrcK8fKL4OMfedpoaY4
gFdMnlzf8MrZ4lQKnsz98O7Agh35dKz4TLgOaOLQ0cVRCXoSYwJehJV0DD/3ypsuveTzFdEI9OuA
7pGXyoOmEd/jNywNVXB42CxoVdcyCrr7+wRySEBGLwLGNM1atRkXobpYODleEZHPQRetMRS4uFqB
3Ah+YBxv4W4Se4vDdtMQ74hb9rEcZ8IY1f9pZs15/0Rd18u3HZNpDov/h3U0w2TCUD6TyC0ThOhf
HZGMuGSLeppfkf3E2QJrI2dpBNl3YbWRK1MwJ7VeKtcTo5gDmsFSumV4uPf5dNDJ7/XUqlZhBPKM
nYsEpEdi2KU3e20bnNAEzK+XzJ53L75Kr3SBrPRzXTvmu2jX7Ga+5A/9RzQm49ploxrNEfWWV7JM
WKO5llcBLzYy1/jyZht6Kwjbsk29wpKz/MvNKJW0x3duxW4+bTcflBmcuZ7mhIrRxPcocLl+0Ct+
9L0p7uK5H9zWgbJ130eGJyX3XSOBDQILzUGa7PMdN+2/7K/srLSUd21uZTSc6OI3vf6uy44xPIFZ
ntJqZzrQOYJuWM+P0QrTCChuTJGe/pvN2+Xd5JcTa59JRdS70f1kWWHmKrmhzhu1I78E5ji22o/6
r3VQjFf+qaMYT96QYFcr2QZ7hPU1P2XR2UCdHm48pR3De/omuH4Fwd4b4iTaBAOPHutEW17sEY9J
HR5D3c5uFm/b444rBWP81qS6adpgTBakRw0o/45Z+mPE01v5Ld64Q9bx3PrYWOOjdEPySORd4fDi
yvwFzizqpLKPWWRU3JdN1TveByoTgEqYu312nzMLcVhkNE3QsuE31cgwB4ACkEC3drXBEdtMfKhz
FIlVsOdbHQW8hT0BaPl8mkOjKwO9v+RkSfjMByLz/SLME9j+Tl+GJRXzJ/x43J3Mi209ZBFJYEsR
tCQtjWZjHZAFRDftzdZENQCjuVd1s6uZNgcTCd1Iaoz9TRtkztalUcW6Q5VCLHE5ZV16AknC3kvk
YIWadxGNnutV9sJchQaf7xDeqran1HbjO8DgW/g6/5pfjSIg/vvUZ0uh78wKQi3PcpnUk5+ECDhz
PEixMRf1idq6xhhoXQQcxGX7ExzEN0nESTn8tRic3WQI7XcgYD3LkgS0nF46WMWH3WxTGqsWJHcL
hhbWBem722ZXe6uifyTQvrR16lUFEtE7rnE0fDBd1cNaXKJg/glBm2rPKzDmso6sGrIxBTcgmwf0
b+IeJKnJIkWlTyYib0xbZ0XlbS544P/azIJdqQMCLkThW74vAzBREtp3FvGJeN8pB/Rwmi84xVoa
sFMAHd1ryGOIxhTK1Z3KuFnA69z15SeuFkrRSl5zqqAQ2EUd/9o80SgcD6sGlEebcyB/2HeK3+s9
xjDknvwEwusfH+uC+Qxy58QqzjaYonOXo9pym7aPHXWTiAMjexISE0R+gNh8QKSyjhhNU/Z0121b
BF8yPQFsjLmXhb+fKKTTksrX8VlUvkhrLhSiYhlu9YEfogYJ6nnEk91IYdz7sdnBNgo5CzUgXUy3
h9I6oyBVrwDgcDoLQAm5Jkbd7bK6XZG7NADbjkIVkOat0nDhtLbuhj0jzugQGc0TZwPQ4lMyhNUG
75CeeIazcxCWiYKSBUI23oOFk9ihFi7lSHeoiTEzQQkAwZxjeNpMKz10YJgMIYhHYmAppkCRFuwF
+QC2KgAIFze0dCnTCGKRiiX5bUvnIMjbBvdcMQKU0/ROQ95PQeRPGKRjnb/qUO4UevKdncjj1zc1
KpPomu5jY64BH0CHtiorYMfWtGUfHkB+l7+4cASlOk1GwHDfkia8uhxSKDZEMmmdSTWCnm476/vq
LvyTxndQNu/UXsnUUxpWH02LT3oUWPUb12/QNM07yE0PjxxDL8AZfNGWxDv3cxRm+DQUaIPzaxPm
JRNq3CX5acOAPMDIT2f8bRmhWlhC0l5bMpKFwf2Nm4n2+sspb2oGMUxcFhQc1SwpB62GM5pifNTd
uY/CpQhmIlrb5HLEodKRlbajK/E0oCwXgDXooBmGGeK0uVNkyi4m0df+OQhcWXaiGZnHXt3NFjSd
MyDrdn6Sys3n3ExoHoBRJUJXToC6Jn5V+JPtwIS2FDrN8WI4HQvXccDEExwf528X8YAqDuIprHcQ
JtN3EaxYmDjb1Ss8210OOjxG/acop+feuDA41l7r4+oybhIGEnReZIJEZtZs3UodE94ue8X4NAXY
hDv9FDn2lmGvSYNJJVbebwy5pyDNCdwvH1GFrZVstJQLo35icquwiVBLWXV9m1SNLQZP6PO1/yJb
gnmXRU1HEO05uX2JN9hWVxPIkSyvwZerN0B+5KfGnhZy8zOQzgnSCPw1XDxPK2cjfmPbTaPK/EHa
5mA6/Oxprg2MNfQSi3hswdxajDrHQuVV1j1fA3QzDfPnmRfD4B6yuO9tFGcLMGp4vmTEWNRL2pEj
ro034UGWKY1HlkjOFmjlhAjDJY8sv2HP8MH+G7g94QJ2WQhqSd2SF7cUams/Zrn5W89u8DP1wVrm
Af9sNhk8D01HjmN6tNVfBbdVIITlOAbY+KKMJz8J3YUnT2Ksr3wE2Dzf/WwTYJEmTwkDti5GkCGX
AlN1oROw7KDU6z3MfzPD5xCSw6T8Do7T2qLcXSQvAT2p6LP7J4ygy2wa26c1Ew/oO2omcEAnf+3J
S8hUNT8Mvp7EhN+cAC7OaFOr0qAvSoWvemlaWpAsufFanpPKrwqNs03uVhxBMDrH7c1lxzg4IBaG
xzbAnNsZM6zgh1nZTYcpZh2+KY8faVayNXrNLiNqxp0KZo19hSlWaayvQr/frqYfCXoSuGxQ9lQ7
ivQ7eFm6Fq+6BOVP03lZDN3srEfmtdLi4AbELu0tdRcSiQcu5mzUc164e+mp8ptzlUI2vfPk22pg
9e4Xopj9W2aJa2eu+HpBYWjgQ1qOymmYC634SaXaD/HHvnMQM4qN8iIqbWi2rDFx1u+ZqQyp75WM
7q6mSJt+NpowqcvJW5HhjNIxj6nECDq3gx5LIO4QYbgKFP3ffbsImX/YrP3AfFONl78d9suepq62
RkO1r3E0aiZrhxUGJ/FYtDw7HdKRiiJeKNVGskJguKBwwILh4bbyZX/K+Iqxe/73qEIky9szJtOK
VTlbnn8Kvtp09FLFCK/YDJQxOuCWFrQW9mfvOY/kwiokjtFKdcl9t7kA4aZjwfV6MFUcQQUTIMEJ
9IASWrEUKu0itwzCm+WQvLl/cb4d6Ooe/kOaTuUnT7g3QYeXX2ZcI9Tjnl5aATJN3Qz+6o5oTe1h
8W9GxHtJJm8FEFE8mxJ4fNYy9BB5/YfCuknYYLc62wQFHlgE6XbZhJ0jgzHaIYlq/hutaEYVei+c
XM72HQf4fPMxrUN5s0QL5GafkWJLdJWxZsspKok3mx0uMGCskm+OHHvcDD5I+j1HupmRW0S+1bmh
KjfN6AsUBZ1mmDmAMiqtfK/7zYc9gfhaDByW40d2iTbPRlhyGqRMpfNng+CaKTDxFmgEGRvJCLoX
b7LeNpNIPujZ+oINfQwWfhKgnWLi2e20zSm44GsMkVuARQiAfD5RyuOjjCHszmwDbFl/L4fOMH7e
NxqdI4XrQhxoarZiM5F57qDBKkgw5yxqKFjjZiL2Z0oPr+yVbNHthFyiikXNoXbTnIRl8BdcbnOe
BGe32TrqBQ4+v9PLklNDZlAhncyjv7xioydsJa3RZEDtd3LM0HTMCYuvA9dzN5kignZBLrzjjY0w
6RUTl1Y7UQfLWvJeNzuSODsMYhKMildMU7qpQVf5lVNCmTiedpdc4MJj6cYovcxxaTx49pPY5/Ff
l8WC7nHzqijG9RYDxH7n9mrKkEhDaNfEpHhgi+jYRWeAVJNej3XU7ulhg1zY7Yio1erkMFdMWbsT
T/n3I06JtwbHkmzpBZxRGB3yc5UVyUBG7RLHWF0misDLElwWf7dbyC80hVLIu71NFccz3yO1mAci
CMTO8kTul4+c14Es7RcNg8wWphvRFqZS090dGtuM1cF8qKce9VN5BpdKbJQZODzA1F2V8g3B5dC6
d/pGP6PbIk/RyAzifRDEKq+TKhazrqcJ/xeBhGrGMSxuXOraWYxEunuCxjszSEtv1nQ2wPMEMmPy
O64TckY0lpEnRyH+WgA5oOePGNgb5xuI94ULyBLHeBLKeZiN7gmOugUZIa4zVgNq84V8dkV5VnIF
1ySawohsBQNmzIonCDqiRgGIGnhecqKcLgnT82d/gpW8T5VTEQZ0TuIT+GploQ6Tbqb3bWjaK3OX
Srjuj90H/P2kEjM36B9Ex7oAkHx93en9XMT89QQGzpy1S0yPfY4TjbaiNuYfnpCY+DvN8huVpOyM
DGDpZVPIcwuaaNuKXwKN15/WwtSMwP2UoAH1d/d91PVW0zkAq2INGVCiK4wcglJ8/kGUUr612crl
csapQMB6CnnHnBgRmnrdfCmrGj77c4p0MBvTsODNTt9T+uFSvEJxbr4xxGSemg/VLHarq5mglQ7b
F42pshAEz73+noWGRT659vSMdvQz8xJTsfJk/k/VaisKXSBRkfc/FGF7wQ3stIedUYyoBVb1FEFO
sIUy+76/4D5ji2kX/rg6yEXLmLHB+UI+j1HqTDFjD4dwZFNpV8tu4MTYwpZZxFC2XA9Qld0mJ6to
vQg7VCepL0WPzHsll+EWGAfRWwwTtJx/QrvTaNbrwz0xpzweAK6cI+4AkP2ft/4nNc88ewgWXfu1
8AsIfuI9RsJzJDpSXDcgO1BJRqGvYKNlyy0qOXaOxFl8qJneYJdPkHKPIRySZ1fIlkdbQWTP9kGc
mz13qA1tgyq9kkaEReMl69WDmN2ryPKoxPBEDpmoZ8fRFZhQ5Z4VzFklsBVThgsrwFmqN4wX3c4/
m0bDz5zSJN/AW6sX3g4dFTRLWEmL1U2vAavL+pLEYfMovhmygZPnr7QgNuU4ae+Jk8Xd4vqxnSpX
hxxTHzrngxs0+PBwICYHGTYitxYvExW13YC2uKdJWWlgXEmo2MMhNVOGCmURlcVtQIdbX+SZaeJZ
tS4lLg2PzkIeMwW2lp5wpUuAu84sqBR4hXKYbpg7bzgD263NY1hHKWc1BtWLkQzJBZ1l6FmfqV3F
I1dT+Gojwmc0JaLXc2e+AO5vqwSdsKWrtVwe2gUz3ZG9BRLrknmDgzMb3TuL3O+o5AFKYa8n1je9
PfRzAtXhfVOD3om0ExL82U3AzYsYa5gMnnHiFiBFr3yN+v7rHZJMC7ZF5ELWKB6hvzEBPV1hIDCK
Cv+By0qdTkK95rxPRt39WiOFjffpVK8QQ5p12xwTlA+68EHIFhep249VKRyBmf7DcPD1EWeAzT6z
c5vGZu/Tlr6aJ2DphK84s7wyYqALmwvg7E57gPDi1+gJrxucONhhxXOYoRfUsk0hEKuHHb/KJfVO
KvEGDh7ZDHe1tknrRvvcLtagSBf1R+trI+rJ3PPCJcSqWfkz169vy5n30Yf+C1FM+gsNEIIR6QyO
ecNNZCiCG12EB8RuBHYp6SC1UWSQ2gB2nLf9FVe7/8x+lQfV+g8iqBCtvb/W4PCXYWjswtZ41hlU
GGCs1h07hgq/DBmphSTqsPyGyn77LugIUxDi1miKNQxPqO38I/S3G4VGRrfGGAHB8of3WLGOoHSM
A6NWk7mm8GkpNMRA9QBYChy1B2g1tCiXhS+LcDj7HT2TPEVdvTSVpzWLWukxziTWxlSdSlKZp658
aMIXNZMKUwUff+1tn5fcEXobd3asBlM9KcaZDkx1D+BcJhgPuC+95ch1DzD5YfBgoBDOHZypJ7sa
shFegfo0HxbSpj8tJgUp8npHQgQMzJv12dhSaMENKpOL1q/Xn36lKIEaO+5HMugw28PFTU3cxmIE
rf8kX1Sxctq+H/sT8lcg0iNqGM0Wfu1JMkFv5Kiy5ruzHZ4sU5ExHJiErM28VDNmh5xZvmKpxgUe
jZphkDveHCTpn/ZgDz4M9dvfgpmOJJMkVjIKBrFaw8c7n0BUmROd/vDXyeVh3zDlmevvOwN71z+9
xnzyv2S6pCy01AfmdTT/Z2TyOhv8qFGnUfDVBk2ER2L6bKp9QVIt+vduNIyVhGobZIEyPH+aIvQh
pMz0RWtyaJ1qPIVThvaaU3gdEYpUT1C9U5QEwkBg9yvgXNVPkVLHGq4ipA3n3TiiTOpmUiBjfnb0
KSAaJHilMZsLWdMTQ/dvDlldslGPFSgq/L/ipuls7hftPVZ6NMp7BrdPg1JIkOu3v94BLgFOMFFO
oqVIA6l0cX5DGTVM6+2WCsD+do+0erhMqY7WtmpSLmsHkRAaAnD/fDRBuLJZxOQjKmVfdMF2t0p6
Oa9c/8hOSgIJHkkASOQT2IqLgjSIQnSdiSAJAwXgWHv9C6SFgwFcaF4oeWse1Y57do54DEQvd+wc
NYKig38JFCrWnoaTFjCZ+89cgGkO2eN+NUSnGEX57YmvsSc1tgWgwsm8zovLdbA7D61c/4AGBd4n
kTx6UTHod0GxSWTSLuktb5Oh/yf1eYZ7Dge5BxCNrZHd9XkDjB4Gs1SpF9NIRnOI2/duG1VuX81J
N94YaK5QFE7DtDsgmFwEn6kz6cEY2QT495wUKwsTYQHZXhBBZ1FInn8NE9oKLWRk00XZnwt35YeA
ZH2C//Zjl7kPKoUk/rU6nLUvZntkKHae7rueMU52iFwwFPnjvfTKGJ0RHWR462Y/pjShNq/u1plH
ViSDMbGEKwOjIWBxWK5C6SbbwroPZYPcNHHji16UwJ22w4PAJz5M/ofDBqsjenUS2/fhWveE6N2G
vRAk2XLf70/uu/kidE2D5HlfqZt1ThBNv9QMZ6hoDJJqhJ6bzr8C/I8m2J6iGrXOrlwaQNow9+Tm
AKdTzW0a676HpKX/vhYjLZBdEHig1siuKonCP7i/8fDEkunlkZKJhP+nR4ZXx2+3LJ8K37gOn4vb
zLKJQHVx7W1kQsYo9DbO72jD2qLCOugu6WGD4MeI9fs1MsGslEOynnx1kxBazbMdg4Zd3JIi3z8G
baqhDYjmjh0Vrvm4bmb8onwDQHtQtWz6ZweNM69PQzLE6fIbZRAsSKRndC7bNe7U1hMO2jk10LMT
NX5Xo/RDCzRSh2nyGs8nRApixAs9PF5o3SjZxFPEle3LE1cVhTj3Lj0U9W3HFvoDFPfhVPM+JJD0
QK6LMrIH4iyYMClmUi6QK6ILC017GyA1ZhILx7RFUgBmwV+wff1i51Fes+BMBIZabPAqyB7HsLPc
eBRHUaRpTQxg1BZrtOnMtZo0yUjPOJT2qbpa8gAQxReemXQ74reK3dWU2Tf4tPUDj/mhWYglpjey
gIX99+t29VWHFhgMvzT1twejgT/nmJBiMMVVyjQDmWnseAzOEM0qUaCa2VwAMZFm50PT2pV7Up0y
T2P8rnvLwkaWMWuGMVZbYC1sqHaKa+8c1K2FD8nI/j7cce/J1czNQg2grsgZRNEU8ybA8GfaIClF
7P1SLVkJ7tgdxIBUcKrHogFCYmyI6SWc9S/UCmGHFoVc2DX2m3oTv4OzRYB1f8drjmuNyPG9ukH9
dmbQFA4ShY6pwJY6196dLiskWxmI1PvaP6zeWiWmnV/pPsD+IutgM1u43XmeD5YTaZJpwGi/kQEB
0HvW3U4dYG/zcwSapUOAEcbj0jyctDbbmkz79oAofe5nnLRfd38o6GYCPSeS1dOK2MwTsAyuK1V4
B6FKPjOKQL6kYb/VZpNBcCPw2R0Laxs+y21VBYUZ2P/5EcJh4YLvmaE0yHLPIgotVkbW1yeVKwzo
zT+j51lZhqWvxt8oGHcDSopQKGeFNtdCnNHjIqU0p4pE4HO+Vx+ugL26Ma9xKpkLlPJgsEJlnbmo
pQ0OunedWDV0RibtN59/UdiAvTohOQ4oAEu9e/nsVdGNMk76xsP1LtgcCsfh//kyJ3omA2IKcWte
AUblCsiPeq3elYBgVTLk/Z4NeINjjHqlKltuvOhUn1YcOAL5L78qKC3cohgAcPOJM9/9dcUNpmML
e+7LaWBawWOc9pKeb5rRmqvoop8U91cXMLtsMPKjOXcp4mROKj1D1pI3rLUVnqf5wnhCDH1LZp2c
DYqsgXSCZqCbDt+lK3ZawZBfWeT/hwzAMcgVrPCVWn4qGvkbM4dpRmhTivuNotJNI+Yxto6OdPoZ
ujE3BoWIxSe7et6FETtOrOhpwi/738jQrsAcLJlNd4Z/aQN/Zjd2Pw5qkZ9+dqSUwCyIxaVd/KTp
rsqrKqGihawS0kbnclQpFosbIm/FY3q04Z1KPBR+ZXSlpTckjyLX8VT9RRE0ZKG7/iVZvK/h+6eJ
6FuPYmiJn16oyyIhIIpP3/Z1GBSV+z8D5QwiEAp8xHBxT5HuBZoOHz7BqVC9JlY+5IYq/gSLwYfo
RRnkkNrKwdomh5clxuAH26IfWiCQJL820yuO1gJ+XJ2Vcf3NRpjLHV+nljXhTB26fdB5jN6TQsd3
C+riT0/Pzvwi23R1Kjr/ealLQoK0rmVk+Smitui52Rnf+RIs69gxu64Z83IbMwDSgVWSRwpKfTQO
1Qk7IShdq2LfawZAKtsQv+WM/Y10Dk3lBLJG9tm6XAOmp9+LratIxy1opVhBEiI4ZosalwbVJOOk
27GAKfVgNajdPPFLcN5jkTFbpxeP67C9hvMdrMUHCGqEW3xEw4c9Rr+PfUeRqq21eohO8+udFOr5
DC4qETFaCKbfQa1mHII5dJiG59Enz5WL3BhUF+xiqxoU7yo5BPlO4XUtanjBueMnZuNhXXSoM4TT
oML1eBdzSaKLgmkhnq8hfL5fZbxIm9aPHcBzydYfdsGhbgNylhp4WwGVbRNZ7y9BBxUka0LKyjrZ
/MZrVvoXZpfaUj8iWGQxwqNOtjKOVllZiyJHbU7zGzLnqy8SCI6g5WIRPlFk9OyuXLJ25kL45x/0
VJh/1Uci2cBwVH2++v1Rjykuq0+B+iubbzwjYlhg3ion05HRrF3e+GiAsqx27b8OB1HoVYg+2qVJ
2karz8NIW0KP4OgsRrVzf2c9eB3LFH6rk77dpfqJlXZpXAyloOF0pdOR3WKqBrGQ9gmgnqpjSQqi
qBxmkwKy2D8QGrbyIjj5Pj19QO8hAGgpyjmmTEEYAOojiAnupJ8Bl5g7AlzWT+3l+mB/y1mhjoq1
A7p1p+zx92dndd7xyV48WoIFSPMsqbQyTpRFAMbS+zPdtrlOCSwVIWJGyO4ODh0454DuEv6dB6AT
muc9bkZ50QE3XT31e4xbh7q7mqBt2Au7wh+iufhku7IHvvj6I6Bqayp+7kgn+GXATy9POQSRHAW0
Y3AUWE0D300ela47kxwAD+RolPy+Q9/mX9OI1BLu/biCmitGPXjfMjoYHuThAgQlhJrWz87ZERs4
yk9+LShfHqi0aXEWRIDjpbvvz1NnlyNh8ji9lTBl0smgrOoLyN+fpxJbAtGfHcDr08NCczGQ+r2c
bkPKW8FnA0YbV2Iy44ZS/roRHdzhCazlKsnc3rv8nGYrsli7Ow/VLwK/xP2gJ1t555cncVfGVXS3
p+vtShQUw4cb9StmFsYhSgvw9314mbkJLX94aaOYD+/czvv640PpW/tU7YidIt+w7Cgws8R4EhWF
x+Y+GCv9M8rp6ufMfqf0HlL+roby3mqYSjxFuQRmeoxgwCHul/C9uFN3PwDamBj3PBmXhnyzop5T
TP1qD5/3M92vC1gnmu6xYYTiWDZwDqFdWrEvEn0rUZN6qvqcaM77lQYVyzAap0Q1MmV1tiE9LM+T
d0OpfOENyUy71I1Rsoza7MVINwEHYO4G3qHTIeDS+bWs8Iv4AFjCbm1YpPLSSbgdO2zN8Y5OpJWC
zN71hmErosoH2aIiUfSina7dB4R3v02vcbEYUynVv4jtkiUv/OI9AbYj8AMZ/tM7mBmUraiBkVzs
Z0oiWozuiZJnen/Ec/eus+aCq8nQ6PLHWfpGNCd/5+Y8RqwIdXlTOiQ+XgoC+ZLbNnMf+X/3wmt9
VS2orTDpOTkYi2G9KuJo53TsPAZBDyHcRirntLfl+6hC6o1wOt3CIoJqtA6kwTxnVIDBQzOEtZ9z
wOq4Gtr1FihM3O1QG17+lbwqckAAgsU+i2YqWtCQof3rPqHxQe1a6ObaCtrLWIf+fQs+KULplI0r
/e/wD96vRzEfQG5xshrazW8JalUtEibN9fajAapJAURA87JCY5jvV06Tw7qiTn7pUeeHtLQxM9UG
Y4nm4KpzIykuVXLc5Peu/cWWxuCorS/5VJFhs5B2qhANGAV9wst4/2lFRH/f3490Q+E0PnWtEBck
jVTn8OVDdDFiyn/DFYtmfixEb66zrhxlScgU29+vtHYkd08zH7D686rtCmEJWSQ10sMrn28Pc49E
hWo7/4zEtA1gBiTZErKG2e1l/a8//VtsRyLIXqw6yzy/2/Gna3j7t26SQGo8LMc+/Uph8jwDTZvO
admTVYlcEnY++99nOsrryuf0zhmPe2GgtB6uIakJu9MXhbszw0iScTjgDDYOK9vNojRv3iLtF3Az
QmCfCwGLbVz3WLdX+0Dgvi7OTpXPvSc+Cv6aPp63XVwlBzQbPgh4IT9T2J8YWstmwrN5HYhbKyN0
Tf8zBp92raMpDhir89D0Hv4p7f+UsRfmZVVK8kX/KhQbLniUJCnSTC5Sj8pugdDSZaXrr30/Pr9c
Kf2Y9h4aRpJdAYOcfKlDtTcZVIUWUgF+ai1aq+lDjbzmID1/MQBz+o2Nxn/kznQiV1w5rfT9Pwt3
CPStfseJeeqbKtp6KAnaIGB6nfJGe9r3d//H/lyRnUb+JobAdPu8/1htBgEZukXB0rldXwJqFKjq
uNC+GTj0czBTPCiSpoOtjvdMjwk8VnxWbp/63laEandRE6sIup/oDgkuaBt4qcJc7AVAJsiUGKHh
HdQhg7Bxi1W5xWiFPEfz2zk4MTEFUnERUi0q8q1HWUiaWdIK1yaUCh0A5IHGpgN7RcOH91Wwefry
v6o9UQtjsBcNToP5VqLMgER8TeBsuFpHxh2PqRcHfvdk47EIrvTXLnjJDqtoZDdr5Lp6gbBdwdIq
mTPDUo2rf+asDpJHEIS6b2mmkO6nuiDP74zoiLJoZ2cn7ighp8FZ5vr+grII0ByJXjcR/2Gmc9Wg
zTtNo0X0895v+O18Vg8eUherL1/sgt8mO9garSeFokL1CInpmIOlj2YH5/NFbHjTzmVSuhoEb1fQ
rySktJr4LZyxjxurkKSoyd/ZPKvShRSALaBT9OecXWeXMnm3Wr+zzqnDmjSfpdkg6YuKZTTsKDis
zxjcF6cs7jY2rxIyAGvXsBICyMGI75V5bPCo2c92QEo/oeruxMG3EaR2PW4EIodr4wnq9BtRYYrB
gQEp1olVHRyUvDNurfhbJbD7bVwk2lzwiKk6vtk+EobG1/12rir+YEcecDt9TYQyyS+7OqyjG7hR
a42hXLdLPDh4l/XCdgQx4mBMEUpH6egzzdLF+LCX9oP105aUBrFmMN5GQ+JFqMbXZrF1LrbYmvoo
FJsccopbj3ROo20h+qM1I6Ui8UM97ouQRLwdxmdwbi9/bWjrsvPI2J3SojUYYT5QWpcJB5R6rmc3
i9fOog42uA9hA+9Jm+OhMRQ2BtnvFypoQ3dKiRej4ZbY1woQW3T0PQ9cXM2AdrXlwgbLYfo7Bg1l
ukDT5ktReRT1y6HSuZL3+o9LkCfWhV+04/ppM+3imDQFhth1yUg65ikAPN2RuGkSgQC67qGZochv
cBMYVtRlxK1EuqKVxY3+zS7y/jLN9QBiZVbiDH5+Ll4m0DSxqmoUmsgnx8/gygjmk40Io7xsc+ky
ia4GPvxCof8kqi3FfkU9BsscTyGlLRsVHxWhF6ADednhuSzv5txOCnrLFPF952l3V9lpUcae57nt
ZcyXucgjVRCf/NgFCEsjfEOvvxOTFNrq1xI3/ihzle2cfffGLOHEJ4+R+os8u7WscfQW88owhr+x
TWms2/ZcenIYvckulSmJcq9uEH8KPrl90LlvXQxrMjL+RKaZhbEBodWQeS4XhWTeMQc0dJjRQxJO
iST6SwWx2M0QCDvCzE1XsiJEjiI8fkngtduxWGRhIpWAQMZlVGYoUj5pjwOccoUp+5q0F8c4eZry
VOGKSSRFMn8eMRnttjHmlkRGHBLlc+U7UUnWUxoDEco32tFo2BC4yzs1m0Fnvnp0WtW2vrjigmr6
Udh3CvDdxRSf56L79Kj6bLd6MKOYBdGbW+nZYU06iM6vqECKAGE7O/l1ZPU8BerpytkQMX+P2flc
BvNPJYzur7Wq2+odBH6WP124DvofuucaqC2uD1Wt2MoShFTh6euhjftVYTvbFfjW8SWiXqjUbacO
QRpaEWru82kUJ/bLFqZZfn2wV4xlaGT5r02cz5igugqRdDWSCsaDmP8zyz89U/aswIy1vtnJ6/Nk
7emkDsDOO/jEk5X8WRCZ61cQUg9phn/Q3+z7HFWX2EzWf55m2gEM3LgIEVnnotBPJb2OH5AHcbiX
TbP1awQ6tRVBWaa/zO7+EhSflxWho8T45nZoPHHITMW3g1FXBw0ux2UygbTFC5aZH5TiB1GhLTDs
eyzpzmIPmi4HxJn/Ozw5UueXm48GwKWChHrdbjnw2bRKtf8LxmbCiNG3G6ITdj91uIXwv728lKHm
sN1Dq/vz1NTIi6OtMg97RX1C3R1lue9o2tBY/Igra4uNBvcPaFCoDIvxJPcQTaq2y54zOdbtlQ6R
71OVFNE2uXtI1p6zVxGwLoN9vNXBJI+apnymyby7A1MYab/ZukWgx2CpPwSgjpeWfdCLdNY2VSQF
e4k4b8GYmLXv+vg7eIZpyqA9juqedYocT/dg/bS5iT5P3860d7i9cJ3CITbe96uCyQgol2NsMOb5
FCOMKOY5D+h4yrFZERwTsIctmSlYW2yRWrCihLXvQ5eXiCQGnsE9iugMYR2y0aXfyNIRr4BNIWci
yd1XjtedHHxOpvCL16exMypZes1M8sxq7/J/kfbCXK8p5/NAMO30IM9eQD8Ec0OLEncVnbRTfrUl
SunwoMTM4lPeeZq57NsKRZRqZcgtD/KTrUh7H5yOBK7LorQu8c7CRgppALHvT8lX7LmebzkZHgE6
j4vv+NnJ83169uXE8gna8psmDnNKboLIRIyP1TVKs7ku4fCEQeB7hxLtOS4vLI89PPe6TeV0RQBw
LW1j2hIOp1xaYpyQc2utTK/tgToyYme19lxH5fyAtzWwWqR8GBb3A3FC8vjG1eR8bkZ+V9ooPiK9
H27pTWVBZtE5M68SwZ81kjHDcL9qLsljSLsHr+b8qh7C9DDng9ldblWNtx8LAGYtOziSNDE9zfTo
R/YWrg/iX7lvlM/iPhXj4jCrPXdtAjaqRJtP4+z8AG9rDifTiqAqjhDjPEOdH06dlDlllulOUnci
Rc8szTwo7UKbhMBlMQh8ARdgGRFWRxb6rPc30J6zBOOT0ATW9P8/Y2PwF6M5J6sCXBOL8vzFd2F0
Y1JYgEQTJ3k2NNFdB6DTbpCFI0FcIrTPJfJynAudlYa332GoKZ+fjzofByD3K4yDyvwIWz2YXiPI
vhjPsSvVGSAEo79/rZbCjFpOutpZmNfYeuYNTuUOON0JBlY1wx1zGBOUqt63EpgWsmnJQq9xoiLt
2nAl8s0m7ZlpBwrABhzqg2slpCMJxZ9kaR6WGzIlGzLQhEkGuJFxGiClDNGzj9fC/rzvCnudt5ca
y+VATSkDVNnq5vq3wyD6/K1nL/FIo7ojXUkNpqoxbEIBjc4nfNKI+Ypp3dio/bzzfRCXXOR84St2
76oPNpioJlKVeh+jCrEeWOhgy9oHRsbcry4z3O0CjfwFkZPfAN7OLNL0kOlYk6TKBLVmWRf01k4v
e+TwYYWrgwsgrRC576YKbUJm06l0QDc2jOwRG/XpoCjf/O5v0hMwsuIqqyob1K2eNT82jJ35YPAE
kQfgk50kliK8vLIhrFrOOwk0Ag1nmV9DkhQIwa+tNBT3XYE6lsY7jed68CU9rc+3bnC8ez55eiO5
Qrd3hnlTCPafxBQj18Em2Eao5ZEPSMO2KQtm67jk6A4m75YHyo4NybAWhYbLOBIXeEPPGx9MT2as
YDTLmErjtoF0QOCtvQvTuvGHy51u4TzN3lp7rQojR/gSnQwd0aQZuVHh84pPS10CgeA18HSa4xE2
VAZ11qV9zg59a/RUcL/ZmBn+RpTj67w36q7ILgWamGq4U7w8oOyYnhpmwSMiTCw5iv6Ri7tF7bpu
tS/XczjBX2X02rW7xFKOnX54v5IT9CuUZ0c2Rgk+qbUmkH2Eorfd6lnhX6KbadJZdnajdHEbFMih
BcJ5IDx/T9XjwZ7uPgH6vDbT9nMqXvJVcpVTeUpwuynvcYZU+9nLZv0IVW9tJImOU/Ph0VeGt16x
Qze7xoqrNnC1pXAhipxD+Q2hWKIYKQC6YiJHmBTP/fNeu/V7SOYU+DfBNp5Tzspo9EASwi01hWJH
4TsMOqxQUnDExlruv/T5ix3emOG8eIKlM+dHDPPuGfCE1NXgcnUd+P1Y7y+OZ21Mv0OpvkUECDGf
mIORnTiIpKv4CweULnnc/zI8lprOfxTfYw3X6w4N44C2Ha7C1HboCwdss4t/f62avXZFkTMtAPWi
5VQLA/1FBAsxYjB63pYr68wQRpDcjBqQehrvOozerBxKnH/Few/oribsR470qmh7bfm+fZCG1CIs
ScbBKeQj09eeRHG7xwR2cmjfogDXBZ/SBMmD/ZYrUuJTjf/SZXLkgsCmKDwPRMi3TigqSeKkl1Zu
Z3SKONc2AdEX5qDNKX4FZ/y5ygwmQhpdvXSvx1U/nlTpToCjWOg5938emujnpiyRtcUTxuvsVFZI
uZaX9zjIU6qoZlrGlt3Q25+UtQXdvt+y//ZGpET+wmBWnuNoPGfA4HjppF5PUbXN4Tuet+jK4Gen
PSmN9wwXZKdry+lVSCtUxSgQQZPdXQLrYls89LBFXfNWs2WNvNQZqApoM4fHdYSLQgV3ic6qukmC
r/+XZhNAEDKNxQqJIpnwnAyQEz0w408MDI34n6P9bCbaTI9BpkEFGDtuxNiWCL2PkIV2/VpdOPmy
AHdjdite1j2UVoqcW3tlmTs/EwRWHYrtFTVpXXW/+tTSr87m6YU/SLVamXAXak2FEgUbMgKS3hr8
2hopQAYNCp4x69Sz9Br4Tk4yQ/2ELvOexFJzf7IqBhDsPw46QqxiknwOTc9vyZ0foqFP+cPiXN8Q
i7JkhSUubQGGONP7wfeDIURr0kGFPwXk+3LQ8r2FvDkNSH5ttXPf6o2bVNHNHEviq7WKCCmc6wjx
J/ZHdNRipD55tNrH24PUhlB8WKxOeKDajB12efxTPauSvWDMKGzmEHhdKjVUT+6pgu3CWo90sJa0
Jna5TRW0u0RGz1xTtcp177+2aJrF11clZqs4nSb1BzgStuigEElPHnj5E1wINT+Ox1mkbjlWvHJ9
GOTlnzogPTFBevG5Cb9EFI4ABUzqCgvf6BvvNAWwpsyvDEcY47zQqGGJI8YLKEPsGMjmAlll7eJG
LuzBUefeuTI4Zu0mMe3bH83vgzRgr76W5qSl3PSSUVQwgqULCSp7C7lnCpBkcJ/+nyoc2ScOXH4I
n4B9VmRIfG6Emisow5kA+G7cOUIgyFqOrnEzynRwex54uIshXhneOOvyiRNMWhEGpXpdLIykOLbU
Pm/csihD1EHyFKXC49/QCDwtgVRepbnJiyDYK1hCSAliGLv1MUNS9Hri7fmwPcFFdNnzvjWsECsx
blkS/gCh+gPevCwFlpBJ/Pr/Mt4H1BR6UFqsY+Jk02dNC7cRJQkI49k99omKbBnyR1Jo4iskXEK0
tXI/x9q1iJXwzUPqTLqcm+widaMS6phkdVEzuYGFZoAwGuf+RRvxQHLXb+1yRDeUHkB4i+KBRoEc
jPsXi/6cPpQLXu9pwfvqdxN44y3L2kLZSRG1xScbYCpZjlD2TYQsIDNYCpIFi7wUGkAXHHEDFbiC
VBX2kMZvYZM1ywkjEw/irhmije2+jr1KrYFt+LbZkhrn1/1A3vnODXHcbA6YI4bkYWFcI466ReHe
vqQYvV86gTJf8R9wBDxHxxFC4vMEkNO8TQeAS/OajoXlvIz1ML0FIGUCxaln46BYqtjE2UjhufaY
ZQPwUvrNGGxyB2TYbfB3KTWIHu34QTipd3Q1acuh2lHdIEorBFZjBwvC91SsPdEYWY0wEdWV+/i9
prqj42tAtqK2MoWz7Ef+jTvOEEPWg1rOj6BuX3xNJoQ0EqRDdPuRIXZtRlTyBgFO1QOHE4MKWbFF
giCGIj5fe8AgSKHDGC4ZL8r9kV+p73nMMIFu3YWvEKddehSE8u+nFV9V9j4uDVcvJK1OQXSz6lr+
lf6lOSarEy3+C7dWNWMJloNGust3EmaXq2880Udbyz2aRIes5hO1Ndjk+pQ8zf9vgqDdT/pUWCek
Qd6px89YITkW17FcUlvtslg3gm76e8tVXDu99Sf6OaVrtzNfJb3+vBk5VNvRD34kDliQ0zld9mxS
Aa/JD9Ipj2oWEuW6/GvYCNms3tCHFRPwCgSkYXU25VekYEP+WMapA6yiTmR798E9OX+8R/qCIwGL
Gua9NZeXPX/gp8UBiR5nPOltYm/KoAZzkd0OdWXOUrm5y9XeVItaCF64URIjotbosWQ9dDxxjh5v
elWJC4yyy5Uq4Mis77ms4LWcO8GM57zI/YJQjiM5z3aYyEy1T3uQFsNReUfUm0TQn1XGZlp1yHye
V4Z7rtitPTQwftUAI06MR/Q2ZgPa/G+9X8uS4dl4GmZjO8wzZdDGqauz9eSb7c1uJerQLArfJhlK
VSlGv5bnwDTkv+vAtH/vJNHERSwJCo3ebHPSzuk59lo/dzRYz8ZDleZCkJbyfHs2NGuMA8E0JiWl
in0eTr6fIXE3cDrKadlVX/yfyMyj1sTtCcHGA+PGJPk9GlO4LGQVIp+F7SpV2funWq/Tq40Mz0r9
PaA6IaFF5rtkXYsUrMl8lmtGKn1ecfynLFq/tnMsgaMKHRQbdVyLshQhotxRMSFPlRvY9ZdaefIF
ySDS8bo8iD7nvxLShEfC1A5LBHLs2jG7W9X3HvC+aACSFxNS7Mbx3iqoMW1okgYD+BlMV76uVXyH
Or1NFVIYyOjptWjXQg9lfPh2AbdHFAWBSRK8t1Fj2pITDcrqECqKx9pRFVxn2pA4DzMHKJu5VhRE
fnqpKSJKMIT7iVfLkhM+LMdWF5KvB+dUVzIljqvuQTvMS9ymoCW9WsYZ1dtN+4W/DB+i5wIMupOJ
e8EzWhAN7t2lKBaoSFGPN1iU24Gn9UQAnRPlg69ME/sjpfLTsJFXbsB7CjS86MteLfHaACeTuSxQ
78EJbFGa2JK6UvPVcClt9UvSfDDyhEAJJ+d5lO3qC3WQI0xZJOt6r0dK3XxXvwL1CucPtMxP40nC
3JyAEb67ivLkMqMLuHbri0pzJq15I8I3IPBohhEj+p6hYbNDlTAMNVwDqDeIaEFD8x/RvIdrgu08
NQ/TdCpNprcqMnjuw+4OaHFeQr3heC0tPfd4wtqIy37pQmk3DFeDztGNkpJF26be4IWfBRNzVWnM
DJt1SC/ZX3VPbVh0PRSyWPOaF2VlX81scNmKgnJK2UESD0Z838cEAO3HbJru3iPtNLmZh28RXULV
guAGiFubXEpodFuw+veNn0O/i+oqDF0rNWVU/wOMlKmsgFPJ4bJazGgr1NdFqs5FsynvsqxL799c
r48Gf+Zxo0poRXAgHmKnovwmNVoCb5bAv59XMfTDmbaf18b8tPr4aleuyQRlv6lc2YfJM2KEY6YT
F0lQn7eIs1Cn4k9KvSEFAjhj5u/UaIcAuXaHFaZ1OvZU6IlLdaomZ79pZ3VnqLKRG71qYJlFuqr1
N8yNPkiGQe6nwZz/p2gvUWz1oiJGnrTwibUcEPBAVcz9CpmQgVWkSqJXvU0sx2G6Utm4EAHpA9Cs
yAZoaocw76srxZntECdDtZNbde5EcuNvGTrTPSRFv8em1i07LH0OWB29+h1IyAXI8XkwD3+DHHO6
H4FlZ22dKnjqdijrfotaGxsqItjvvBKjZln//VH2DveabsqLVRWUoqlwdJ+wjOe+psdkOEIWKgGn
RxQOWyF0E7nxYPPNi6tZj66ug7g5ueli2hJ2t5o/+Yxe54W0GlLy486CQKnxe9JkMvKV5HlcqHhL
/Q06C8FnhTkdf2luq/tArwfyZ3vwxp8PgMxap4yzqFlhFQP3F7Vml/ti3aM7WLA7Yaj1hc9kkPxx
+ybiA1pL3KWe32OstQpbLDaPR6FlDqFfX3yL8K0KW04sM5ykYEC1nExz7XqG1CM7jzDHTSXBIEDu
eYBdOLmO0NcTjqlgfiDUGTrfYiVmRMR+6wMdnIb5a8kEIEQmCUEr2vbApHzJ9bs7XSYF1DhfSRYe
gDcIEsZ85hyWtI8DgLERDJRumy+wSxZMRsxL4D3OLfU0HLKFnKYPl3bHuFV8fKj8aUMovPuzPhnm
QpakjxbVGgtuas4EyFu6PLCg9wEBZnB2/ImL5+UDI1GWLxe2p7a/tUA7gdykBz4ECVQ6Kn+wIJdU
aZbELFGqp6j355ARwWc+SQJNmaGWgfrSGXvwAiD+G79aCm7ZiNzUTg1R4KNcnSC0jg9a892kW6ed
GEyHppRHb5MSBU+Ct0MB0PI6Wo/YhM1AQM8UwJHCntDXJrA4bLbv5+8VmPDngWKRnX8kmDXQXzQZ
LFu/rZkYhCOqlRNmWOxxm2iUTxUwYaG/ShU+iuBqzB0KoM23LujdkIoaZACXfAz+95cbUtqTi+lN
dBklRqrjcsv/jLhwUkBU6oT7WiiyxbFPesNxvYq4/WisQfaRv9PArStcWksvIzBM6w2WiPDY2JAt
GTng0MA70aKxG8wcWJ5SodfH7LDNUiNPn/HOmSQHZdUua5zd2Qo8+R64iFMQ1pqLutKxFDrWP8Lr
zdHeJp1rRr8F70QgQX6kP4ORHayE072SBjLPkV91V/GOyoLfGBVQSDD1EA8mDYQ8tJV0sYwzPBFL
gAGjZRAO/Iqo9HBB6OiJuUdlg4m3LrKRZoKFg8QTx1ivv1XHNopyBDQbkmUHFBkdlSgVYjOfurTO
3eNlpyRGAbNcdKniaf9qjWeQHgl4D6T7SakFA2T5qgOK859wFXIxDRxBuu5RKF1xja67Gnv/eyvA
QWjlWK7zZw0FBy6uZKyfJxr8vVRDxPyD8KfhUBSZl8j0zYc++p8rv2DGfQr/vx1wxNDubF+oP+5S
b4ycH+fgC/VWF/fmxHZl3a/KjZq8ayawhcS0iWirBvAAla90GOUHjIppC0KcRgxpHow+3sjoS0c6
+ksR9qsD2J5Igm68SczyQaH3f5QIuF7OextlIidD0P3xPUmK6QCoHIR12Sc5hOpO8KBSYVn04bHH
pUKWRvlTnS9hvKfG3wJw/18SRVJjxXKJpiO/cHsslPhdlBAmuoZNOx3/PSbzYmdSs4kMXTvmM/dY
XtXlXlq26u03YK2TuBql4KH7gOin1tKUvv00AxMmvnkBhAYUhKjYeiIutUIsEtVxymPyReqTUcsW
XzdMS/ZBpZXs0QkYrsQxJ0ExZGKQlDnCYeVafv3YspySK4vpFIgrQeCu+xVVAGzBux1xQoJtz4PZ
/CQXUylv3LF9O6aSv6Cq/l9TIkWmxbrmIXziWugyZivci5P5lKE6q0WQij8FyJNRxHfspUQx0loK
NYLOmIjJWhflJITjyq8DZJiLUZnGXnz0YnQRi5CUxYtMlMTGMxo1D62yxlmLlLCfnVJP+04fFcie
Mm0sDzlao7P9zBvT+jDVIDHHwJoFdfsmlF3YZDK2biXCjs2IKMG37Pc5l3k8tMxk2C8ufGG8fg9o
nGqnogErLXscSfc0DqPp97MDRYzw+0u7EHbJpGluEChzGV36ePBxsrK6A2qdX+OgQQ71xHZkVCto
Ax1TC5mnBYKXh7jnwXDc27SnnI93+0dWGyhHYCHgeTkYLLRdEBNuqFMdIOtJjjnPdNW+6BI0Tth/
W1fvHHCwpjdjSwgOtd95ZNNZhIVniBzN2p26hYrHqgjzG5BsvSWlkUAkvOfOgyrs+OFGhKrhj7JD
THZLh6ce0PvJwms5tsSmwtRWyDEQexnJSKTk8/SbzeVC5RbNqqLsGm9nOf0Ilfp6g9l99oS+4A45
bxwHKjbc1JzZHxC6XJQfJEkT2DCcd+u1kltIhRk2L9D5+OfuRvpuCmakkF5SH/xla+2W8HXIOsmg
gtEAlFh0HID5RBvvChAeLF3ICmnQGONv2y5KLye+g5M8P7W8m/gpX50/+gxoWHS1aXjQ3xtIXV0O
VsFAKmhDPaYyC6jQecklu4T7/xl1b2U5+SZykcUrCfc0AafsWf1ptjjrsADBnxizGokCsmcwGUOy
upvO0OoO9fupsrTUx4H6Rsx7hCZhi6O3NlKc1tJ4PVjlX1AxKeTdOGpeCDCPLhqvbtyHl2L6VLFx
Ga3w/LIKbl2fDYHiKmmC/YBmeMV2vTBjuEgVYiB7Ta+/32eSOs6TioqE33lkX43HdmPeM/Yy5fGk
IDtx0At6k26iSNnG/XPhRzKrhp8cXgsLxAwvaUeJgpeyyUx6uquuf+N9bDOvKHWzXGCZVzxgdt6x
VtW+CpQf3CuBWvj7+jw9hVFS7JFyDK+Vr0lMzrnz50+LT8GgbeYZqsqusvbN4goXoCSmZr3rbyCj
arHMf/hO7zdpxmBpNkeQo/FLmiCFVN+d5y/mr5sbNIAcix2NTdUl8/Bvc6RS0OfS8SQj/NOh+ZjL
DUMT2nDSRVBHSBInJwcyIhEmZyPP/Fomy+QgulXhJeLJR4aVKW7cGMPCygDQ/87TVvcxyMRyMaG6
W67tnkipTT4XMlwVOjcLYjWIrqO7HqG4c0bzh1jPffT157pZhiDl0UpUe/dzgalm4TXOsWnfZr4w
eJbzYYNTBlfQn3RjmLhaJty5fSkqDYPnJrxNjD3JWpviPvuolAVRWdekfj/dTME2Q3q+zjSuczab
u+k0tu9TnYTyIaWRXR2AVSctZet6ru9Dq8GaedfBj9RoORZZYmlFjpTj62gbpDba2dC1TpHdNmCJ
rhJaPzoaPn4zrVSkEq6HOAEqrSVbb74iSOzekwzQNZMWEcxcwEdPPTEXk9n8kU57dszPmKhbko6s
qRwlUneIf6/qNDS6rY33wWj0/qE4dKcMe5J3AnIywEJ/5aH+T67TKZINpgKj+j3AfLNXCzxMl5a6
gxUfU+c2bUXkIV+PKdW3/V3lbh/rHtPESWz+nb2InKODwNP3HatbQYEdrs1u4ckG2W1Hnu/AQERi
4nwP7e1riPLhCnY1zM9UHFRfDgYcds/Llu/r9ZClKaeloF4upELk8f0P4CAuNRmz+ir+8vB/K+aM
0YkdJUp3DCgj1SGIu/ADSKMpb4X5EyHOf929GwRimzgLYn771PhB58U4r58ST10yJPQKt3n+obbC
8tlRz1ZVjELhCWAMaMAICHqqd/OKbccetCUHH8uC60MCxz+6wEnNWe2AxYifA+l+6KhHjqfKixl9
AoXtsDkDAKyd4YjCfKuMcMvLU1e29pbQnb88nLeLKYTDR6rXmeHwJ8+4FS0ABsyYUEyHytkDDnoT
UR8tNWz/stHN/K7/FeVKU3+yLuaHFFTabOxWvjK2fpH77h5aTyLoioD508QzbpT3dvGaAmXbNI58
w4ZiDdt7gtWfpKMYKAgqBHutVz1GE4dtWnVq3demwi1h3CEq/iivUy8FPrrc8NyxRoOTXk0v2RYP
3JfViS6+Dpk4FcJa7kTJROiF5cUNMijEjkBq/3IdAnSmah7g8aHzjkHZDRrJn/VHJrb5iR4TGKwL
VpIiEgxsx60JXxm8PypIOGQlFpIxDVDkkhbh13aJp3Cna/Gz4s6Wz/VHS1FtXm/yJIPGozS2uPzr
Lmn2/1lFaiKzuyK98Esb/j+sWH9HwoVMoS0v9VPeh+K+GYzxpi04UtgwAL2f5xbu4mYhTPa49RP3
BTWlpxgV4zau22yV03DeGyFqjZSPT7YowHPz6lUDwGm2F8cw8VmjNa/4XR3UADdQ1qPv8r2fQvPe
U1njGDF6Fd1frzKKwsun+NS9BqgvN9L5JRsfl83onwHFBkYfsrbt1ltKrLtoewxbpS0PdZJCPzAb
d/zbHv0hVAmetowhp4zP4ys7axXFA5rlt0v5msJZz0Rx0wn6LftswKCne+oHi351Yu5gpR1m45ab
TfhBB4sxu84chAQcgP/H1nkklhr7rKLKG5jS49MFYNeQ1NdsPHBSjKczU4pwXIl7W06wpNeKZcTX
1/PRfHPf5GtIEJztZ/9C2mej2Fg73OO8g7xgcs5Q4mYFxMfMwbe1IKpOcd1c79acELmbdgD+k6hB
4zbN0Aac0+fhFJd39zlPUJpnsSaLfTLASPquQN+6EkyRcP5BXLoM9C/Le2SzG8IKeEK0qum196FX
KUCwx7FWQks43bNSfjdaWizIJPVHE08vScp67IL9oat92084rsUW3H54aRtCDQ3kPAeOD2yZXvBC
3JRelTfAERZtZKwKQuEFgrcgIxHJY1JT+FZy2Ylz8rSeHbZ5pXie/9QfbWyXpFaps7CE/1WmOJ/w
0a9emOW74tLPZn8+Tg4ggWG7LFpkGXt2K1Rw9bGvSxgExOF5hyuoK04J8MiynH0EpciEB1TAuymG
gTin6VrjKFTNvGTbG1XidREEY8GzrBEsyYuvdZZ7fzDZs+j1BmnN4GC8mnRCdvvYxDUw/57OJ1Hf
97h7T6iKtvyYfPrfoCJ+inNcuF3jLFjD8ziEgx0r0QE4ogqWkdzHwFGad5y9DV6ddqq6eRB4Bd7B
CGZYnNyLnN9SpL7S9S4sPwrxtj7iE3EOZ42NaGcJKn2C3FDZHXn+Yj/dazyRYaLoC37s5hvZ7wKF
Rr1w+7c41OLVwjOlSz1vFL9g+DAQW1mH5b3URuMIphKXWdYrAv6YcnB8PPn1IA3ZbZbglqhOKVWq
kaU6LGInXVtKJ935xj8SYweTgVCb33oQIgaguh6qcMqaJruFyPzT9LuKCJTA90XoMMNWevXbxQKE
BCjyvHBhhHbCkRoPuRt4g3pYH8AcvWEcOxzxXAxdCuzTSmwiY9908Xk+dzCOi2E6wK1eS1jZsRIo
OO2gyhGyNjJiT5/cuKMNj/o6XHh8KLDujI6xL0Ftx3lMd5FIHY89zqfS64sbQOsjgPUhdNmiTWZF
zXBg3AfoXGDTDa4LSZbHmAnxDhlDgEritVbH8uCva+IGZMVD6fP7Ao3+t7nPI2Kry/IMWh9MRuYo
GWpjqsIQneRC1hA6qc4+UTtPldWkGtq7tdDNWIJJQJrGJhtybueV5TWruYjCfBGkP7EbXjx7r4Zv
I/3KJ4UAdSLa+LrMKLgphTs9NJZfIYoKSHRZrEGCQ7Iw26lbVieQ8YNyacxfmOVHrwwj6uVforPK
uvw3aA86y16sk0RFzbG+7ZCbQt0tMk/FNTsS2OvE85w+v6idwb6/GfWtJumndOtcZ8KHU9r/X6Ym
QXjOZms8Uw5ot4RRJ7cZTpkwXy8Zbc/asGjFke+JIHnJclcaxq++hgRDHUXiWQJdlJaKdOwe72cU
Djtxdzbi5wCdylm04xOK1qC9oC0VlxR3Eyxpj/3tVuX9qrWnP+lXI0Q3RDUvQS378X25FI7rtLQu
RNnA7/PhFa01BAIKWAom2yh6r7+i0dN0yk6FlazAOLpdWSc4IH9oKzJpeGDjGHMGZT8MYYFOAtkz
xpGVuS2lrxQwVD6L3zjg/SnGeBCYFeFbKXx1nHBYsswgY7Bxe81H2wSYqnk/MgcyOtzR4o5eBCXC
hUp160C/0fFpIV9vVsq95AJqCcXCS967vKXnTKeP3i/guTFFuxjYfKz0D4rzIGnScRgEbz3oerWM
9zgZNgADCN1d5PLV2gJCcXK4nXtqXxKg9Gxpf8XmEYnD7lobTImaD3FRImQX4tuvX95XzZQQMu6L
jZfuxUb2g2+NK7GRj+HloSuPfJG5PTjW2j7EycRSjdNFmXd0XB+UsvUk27KSpXHb5OGXgPJf1ABg
mHew9MSerahwWnKdh1bGERt/PpKBOzbXqUScQHuFCb6pgb4WwNsMd1/4jlj67QY84o5tRPmxZreK
jViNhMXbNxUvVMWPD1NwND5zORq0l8+F0Ad+VwdZBe30VyqCeGsZyBMg8nUoUM7wst31NlqrAWEK
eCmdVnJr4KimNs8voKWdLyVeHwYj5ouaSjKizV027J2ICFwSvxSR/yEIoy+PiGfh44AOazVIMwNT
hApGDAmmVJjoUV2Xk3eEtE0xkbg2E2FmG2fHG+qLmSlHO/58WkED63JBNzAeNObl7CzTmPrSQ1+K
/AeTyMXpa1IhTE3lCKjrN7rP9ZxtXfjdvNCvVqHmH0WLmvxciPZa3DOmODCVlqIE6P2zsmSgnIWq
b8NmAKFTlURdDFU6Db6KNUWWPZrliPMI8uiwm4dYNqKUUGYFkTjKMi3w4ul6dtOFDSp2OLF2g3VN
W9F2n7jQHiAP5mOABgZCFG0dQiTURaOnv7adpeMBmLIF1PCHpjlSbPJcc1nl3nYm+ZmNebIrOMPl
QmKaeegSo4pgtJwd07REPsdv6opFYUJ29R6SioKGK+A2j1bGiA79ncspFepavwh5Ojyk+4UANxwu
LNE6GXl9U6hHhp3Es/23HtnsOO3d32+3cVEGgq4WFDkDwAMdtZZGT0YhlM2vJsDGj/Bv9tnL3r5E
XLr0ajjrzLLsMacAyQ7wb7C4AvMkqhAItw8KcaXqZqyczbgMraTr/I/dwF6aNKsYtlEAZv4xUH2F
W7zGh6qBOo49FJLi1/WbSiSkOKXEfUGBrmTZHlJt8ybG1qNddt7wKEFxg56i3BWv9YwlBeRHx1co
K9H8Q8VwHPsjXQrBRnyjpGCfbGzm9Npag0JQc1gUQfxqd8kiyJuCGLGSqlGFXj+svQS5ip4iJLIR
YeethxPUZcmEdIVwG5gunhDLnCOS0Tx6vIOusoG1G6YVAaZxBlx/hIwCShyjfbShn7B8ezubi5yf
J3NFa+q7AJUbK9kfzVCa5xRBo0EptyFVictBUjfMARe+sbHTwePygETTmcLAZ7V5CE7m3L6BeIL8
nNb8nzT9+AOSsrJjaYFLp1C8Qq4NF79DuOEPItocA6NRINb7mTFEw/g1wdCwfdJBOhuV1mvqX44/
GTXzNAhN9pfmWpscrtyMmyrRpgxrW/NR7fxGd2xXnUqNnXDs6B9BlaBVEmlwkGnZbtTZx/jJhFCS
ZGOo2u7AhJE8CSBPLao5fcdD55iMpjPRcQH9TQozbHNGEQqz65rNGyS7Ulj4DvD5cofvfnQPQqNT
sMO1r7gwjmOb3olz+tkSQAmDEA/OzlVSmcPUMSXoN1n9C/qx/qifZsgt6BAplcEBu03tXfi3yVGF
eT7ONw4m/0K/fTSUE9eldT8y+WFXPJNCttsuHfq0A1tL5xf6kCylYjriWg5vLmQndkSxys+wFzm3
m/GXjsRA8fqWfD3iBtJJFgM4SlL5aHk+5hsmlmbosrF93/aLyyZpF0/gaZmaIMP6xLIMCEMZV2Nt
cOirB9y347e3rzaJmX3rT45FvT3NqAM2Fl1o3bmraMNm5Rqi0b03hVdMkmeq+ycUaWubJuHPPkG5
UtLsk8XxIa5l8tbEIW4sRy9/pR+bNxktoZ96a8FgtCGf4JcqDStqwrhmUtUJ7uAbYOwYZy5tLqjF
x/VP2pb/KEXblhjGFcreEEFc63vjR326AcRDnt6oeNdTemgXJ4rVaR6cfn1xdketZSqg/PU/S0qv
2XSb0eoNq9bl4k+RP4iEpGGnRtpC+Vk68BoK8+EoruIzf1oWDVGy6s0V81dflIMlTQSkcV4uRltb
wllPYSEMbn+VIC6Keo1ezyrDg6JM+zurD4DOd9M5Z54aqIaq0WVdmtMtdJ+eLz+zviRXRYwd+MJh
9q9QYSzErB9u+n8Yzd5kRo1SjBRNFzgJNuhqGWDkYv+Kwr7xFAxWiMvBy/O5OYToaEJSYX87pK2n
FlFTOhtvqq11Ieui46Hjfs+QzTL+VBjZXEw3so0OUT/hELDXatY/sWKAxg2RKoE8ZcgftzmIwZj9
M9qmiJRBXk8e177BK348yH9qNYtUD3gte35Px6ZGx/OVZtoEaqYhlsgE1KCY19Xw2SdQY1s7mNl1
sSVgZdxjdlPeCqv04Pt4JftikaY4a0k96sAidoWRnb0tOVa+r6V9EQ8JDXEE5dbK/HNd47CJQLnX
s33y/LbZQ3jUm4zcah+P6sR3ZrM1D+6FQceeZFdgwhxVk5aeBFohvn/k7vzDF23iEC4gpNadaola
veAa7JH2VQw+h6Q9dKJOA4HmQeGOK1LUw+kW5E/2RYtILFqutR1aIacylrZ4glbuZ/ZKstxi0IWJ
vBl1ZhG7o+GuxrpQwvJMdLofut5uNt3qjhShMntlbhBj2Idb/eMooXpW1hz+UM2U/KexA+mJXQAM
Oi+/f/EaV2n9KcCKdHNSGoB0vGfXzXBErs6FcgDPFG3uwmehY8BPwtu7Zg3xidMYwXcTc5x6XrY6
G2u0qYH433EucN0mSDVkY90iDCsnhZzbSksBDebAa6SMrtQZO9qX/OSuf1vxLNgwri+n14LsLzeI
9nDW2m/wtxWPvL+4loNG9cCZ4zlV4c/b9E1QwqvLSMUG1B9PCFw5GxEeRpEvt5ZG6SKhEy85/PZT
sDEs1LUB056wO+l6EQ2nZs4NCUbzkT9KbPbuZmMkRPkNKNFv95uBzCmJrtCiPcXtZur8sbW43zvw
ghi9TeevsEWQaAwzzWYTCJyrEuOZ6gg0p+Yf/HgHUaR0r0u+VWKTjdMfDyelR/1sWG64Xe1dHswx
iYoeVbm/vY8c9MIJeLJ9BcFGa4nWLNVSbbkgw5bBPpLX5syg5pxIx086yBeqxDoKtN5DLBSDltLk
kSkCk5KJqKGUqvPUOfhC9NBzS+b17rNyGe1gPPKRCd/1TSnKEhBpCAuAJbXd0udZXSPZOttXnWbW
UprHPCVexcurQuct0O26+FZILPsPBXn7xLlY0Ks6PuBErCtXlrJ9S4zvXkZ4ZxrBz5wn9QzJ2nuD
hcPXgDJBJN8fZRKtKL29PEp+fWAah1oq9/I7wLXlTcIDO1ElQ88K++LeaNbf7c1aifDTlLmOpc+r
f0iir9Gc1S7hJ90+4jn8TdR8suAAW5KK0w+tndfpf7tJ7ld5l2TTgW2ZPjttJE5wD3B39qSayMmr
Mnbt/bfDgUKG//X+KTARGeTu2ytPt+N6cUWk0zR1kw2fH/lLt6GXeHBUapqQ+9c1JnjNCzDXnJ5u
rqTELuageTzJJkW8xUAPM/Uoeo7NauWHHcH43o9Mgl/NkIQ5wIZ7i+S8q6ORVnZwCnoQ/q6PEaoZ
NT9mKe6+oDGoCrAL8mOXmZHAJiwCgk9yWQjASDxtjba/BSRk713Fe8DKr7LVDi3uZINNo/2IzbYY
ICWM0VgewAp7HaaDnfY72IGv57/DpApxyrcVPuvvIzrKrGwO7/D+eJsGRoMdHQYcw6EwvQjzuIM5
aDaj/9hlx9Px418uNw2M+IMk89wTD0WpToi7+LkeQU2qXm4i9oBES8aKuUHNjji6CpsNDjJJNe0Q
0YpWigfaxu2wSlB+KMY1EerNVcRcNwFjUwuX35ayj4cvpSg4pLFIiqctngot6A7LfH7Y0Ih3xTS+
ABdSDARJUtXWS4vHxLXAgbzlZrgqQtgcWrYDp8sW+KJqSSSOjtCDvAKcYBXK5i0he8eTzhPQeSuN
1nKWg9BS6RS5Uf1eqYClubMHUMMWj49ZwWEHuwRKtYfvOE7HzovL3XC521GGQwE=
`pragma protect end_protected
