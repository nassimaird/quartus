��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�9s��	�si�(3��Z�^*T�1�6L��
:�c4��� �>ѷeL�x�����Yylk����cm��/���(�T�Ί�hM��Z߁�Vj�V�M��im@�F_.Ei&>�/�f) @J�H��|?�M�1H�{-%�j_eɃ7tI��䞺x�?hC{�����pu����;s8�rȬ���e��1�
A��SJJ�e�j�[F�X�T ��=;���-�&ӯ�͙b�i�>���
���1j�E)��z�|[�M�'8�y����9w�[����2�{"��6��l<��KqGM�zٕ�� �	^H����'e�I�������B"�{|������SՊ�>U:��������D�P���_���w*��*�u:���oD�T�>F�ל8��T@�kh� 8OC]�V^��9G�1)ݥ�x���}�(�g�K��bd���YT*�N�vij��U�D�`�yx4H���S�zl=P���M�����H1V�W�l�͓<�t�42r�#Z�H��$�S"��$\W�MiݏRT�����>d��s�DyGNt#:�����do'g��OUd{K���'�R/M��p����z_�hyr }�?*�2jiь���:(8q�V����)6�$��R���޼b�� �p���z_"DOg����( w�G;ƾ/�?��4��K��� ����[�{7�g��@�����a���2�����!��.����PB�0ǭ�+�e��ΙY�>��!'���I�I�B���C=�>�C���a���Sq�x�28���>ٟ��gQY��j��]���8���A �f�oA��$�?_�����B�����]��%����C��ji8)$S��*�����U�3ѻ(�9�v����?Dc���=X�NY�D�$�C�|L�0����z�B�����)�8�����د�σ��=�P9�ЂNƈ����w:@��L�uL-�1��nXF��.�}Ψ�Aiﭯ�~�![��I��8��K;Ֆ�c�P���3�!)ő�֋��7���Xб;���t�KG�m?��<kMF�4�B?S���6�t�h�6W�m ��%�?&CI�=Mew�3��r~3�3u=��OQW�^�؇�I�(]�h��tT��/�S�����\M%\ ���E]���� S������#;:x�	���`��Ǩ�oe�^{V�x1ͽ毱*��XI�g��G;{
 �XH��u��Ƶ)�+]���M��ׁ(t����v2�!�������!LT=6m�L�{(�X����U�!����2���Z�R�jˊ�v�`]�%%H����^2@d>d���.���R2��8�����8���s�N�
���`�l��W3�pi�虿\���4@�+%*DԾ�O�����J��Xztb���q���� �h`��!Oě��1��B�u��_AB<&�=q"��:���۫ �#�݅�*m9�$���ps�)�jc��k�ݥI�L��ܢF�Ҏh�R�3�����KZ)1�ᅆM�PcXz����Om)��c	��0��b�PK��.6�_���jb�I���q�d����R?����h��w�/g�ؑg��Y�49����0dC�}iv]j��fN�h�F��iyF�`���:���bLB�xW%ؽ�t��Yz=�[��
���>!� �k�Z`�$Zyxv���C%���"��T[����Z:J��H~��Ք���\����6r9���&����	��r�C�1�:���y�u�^E���&\~�<�Q;:Ė���HӜ��h��.N���]�����hT�9��q�"I�Ҟ�_�TP���λp�΁��?ςS7-(/��y��S�Zk��h4��z�Z����{�e-���P�{ ��"%lT�����)�f�G`���Q���+�=Y��O��a���r����e߁	u2��H���,u��0�:(�C�!(�\�1�W����F��UJ�	GA ��s����Ig%_�w,�#8m���k�?qa��TŢ�;�<!��}GL^���d��k1�;4�q}��(��	^��I�;_}�q������|����=�(��B�1Ta��9؇�	qw�PQ�	�.$[vY]e�h@Y�.�2�tJ�Q,�������!M�0�P��l����6��Cz�9�@T-����W�B�w�q}<��8���4��Ϻ�v�w��Wm"2V���3?�+�d=��Q��1V�K�o�Old��֐�k`�K`	�^գ�s�
�5��ٶ)�i#һ&1��Yc�,�#6�~S�ٿ�!|�t��+�5���zp20�\�;��94;\S���)n�6���ڳN�ahK�A&��@�h��_���;��I������"����� 0��ƭ�V'���C��$Q��i�ǝ�<�`z���z��
��af�ʻ�"�ya.��|sR<n����[�P���5G-�E�L�=h���?&4�=�a���Q^����*zC��&ƎW�T,A{%#�=�զv�"=�Ui4�g �؟�>E"��I�He�{6�>��_�*�6��Ak��.�Pb]trl�zr�_IA�?���8�j��B4�K���DXRՓ��P���@�8�o�kr�����R��k&N�I��#��� �S��*���/@uqi���%/�����
9�]R��k��>F���y�L^�?G �#*kY��k��B�l3xW��;�7��t}f|'c���V8�7�m�U	Ŀ18�<� ��#ҞD��;z�8��m�a�#�O5�ٔ/.$�M`bјfUک�4��:�Ə��1�u���A���v�u�F]}���&��F"p�6+�o5�|:�tS'�;��k�Cpq$�GaZ��Nk�D^�� 6dh;��|�?�3�	TV#`VTW����x>��&�o��w����䪺s�.,���K�
������.t�ԅ�@�r��Z�Ii���"G	�B%��r�:�Pӷt���^��MK��u��\�UFbwLun�p�b����y?ވ�&�)����Q���ZF5<Ry]d�!��\1l��[G9ݓ4��T郙�7��l�:Q��*���~\�t�������a���ú+��a��'�ӓ~�?3a�\�[���b��G���(�|Mn$�:�VR�OΒC\Rݑ��z@�NSe��8�|X���Jf��z��s-��Z@b��_߫�>g{֕Ey	�q�b���g����9�)����86�Ů���>R}|&W��{����%���W��}��5�����6Y��	'�A3� l\.Z͈�i���F�Y�{�W!W{i�;H5�1�VٝTؾ�͔rѸ(��p��Z��
�K㙚����D�B�<���Q��v��b*�˺�Ёy��fp ��*�E9��my׆��>޹R�O޾G���rN���w��q��ĸ�"�t�.�E�>���"o /L������<l儣�J��{{�.+�D��N9`vQ��T�;w��X��<�A9s\hw� )��o��-�~D@i;��χ`>����a�X$��2�R@��p�6Z����R��`$ �Чf�qz�6Uδ�u���"-��ux떤�L���*�� �, ��:c����}�^�d�Az<�q���+��8��7�E�K0N���v'/�ع���΅+�v�O����yē$j�Q�;�����na�)��9��P�J�����I��;�Ư|������N&�SW��Ok�7��Qg��uq\��oS��Z�.�@n٦�Hu�sq�n>�E*�S����K
�{@E[ ����D��YdD<9<�E2��%# �9&).�U��A
FCS����kzØ+K���2.����b�m-��/��e<�R�!��DE�p�9�ƨ��r��Yh�ߋ�6k8�MA�R����!xnN��ϋ	�o�^tm5x����ϼQB�&`-r`ar�a����b�d�E�y�<�������>H��S���ȗ��,�}�r0&��~4�Z���A�UE��;�A�qr���>�(�D�M�j'�* u����49�� �~�J�R<��N5=`�����}�ڶ�Pb�H|}���/��j�s���p�L�؟_��PT��8!1�&Nd�)��cj���;�4�RK���8(�hk@h�)�q�7�TC��ܲŚ+����M�|�M���ox�1�ي��fⶉSOg%9y���#='W피����[��ߜ�\	��U��������5=���MM4�����Zt6�m2�X�����<�Ϊ��{���2��-^_Dy���V�L�O�{�N�w�50xS$���W~�u�����nJ,l)|k�x]��������'�!��b�,g�"�]Y��⌽�q8`"9���m0bTF$�+�$�4M�����Zw9�/}�R��F�@�=ET��kl0��yϠ�@q8˜�֯�w��Z�|��lܗŷK��ε&%t=Ǵ��%"Jqo\�Bn��䴜����\I�� ���|�HLX�-�G��e��0�;<<)�e���%g��hy:���� �I�ˑ�.�m���7,�L�����7�z�Sbi�6�؇:���k�!�/���o�����u䜾�nc�PR��h�r��-L!�n6q��µ��P�� Sv�ζi|1���~�HW�H5s~�XOt�D`�֭�Jɀ���y�[��\���Վ��R7ދĬ��\�~Fs�8� ρR�˭��N���p������q�������l�\��N���v,��6t��f�Q���UE�ޘ�j�T'~���	/�'2i��#Ο���e�h�Z��i�[�H���}��L�B��w��O��N&\<ј֧z�FjQ���1f�ۊ�K]:_��$0�/��ȲV%HLU7+EbS�1ƶ�����3�^�xk%�be/�r���p�:8��8EA����Egm��\Q�r��>GQ�s�Y��-��|ߚ��0�p��3�$fXW������m��|�Gв�����B�l�����c�5�� 7�W��K#x'����V+3���|���l@r�_d�2��%\;m*��#�~����w���X�a��r�f��T�aR�D���+A~��Q�V�[������i�f_����2�#���-LiH�^3�4����Y��o4��דBF��w~��.~�������,�_Ͱ��XB_�h��긟���-k�:{F���۶�Oj]_I�����y.۹�u��P�c��w�;-�]0O���7�I�@���b�T��<�&�Z��Ύ�f��?�u�+�&mi洝�R��-��x_��ו�Y��=G"!j���"M��~|�lmK�8H���$\�j�a� �#�6���Ŷ�1=�����4V�b��%G��|����S2\��"*�p��y&�8wo��:�
��^e���1���G������5f�q�`Bܞ�d��AOƑpД�`-9��w�G$C=N`J��]Qv����@d6�~�|�!L��h��<":w� 뵮k���:��$��(��9�θ��(ܟ�,M�/����saUR�G��(}�&�}fM��t�Tg%Ѕ҄�@t��d�1nkI��e*!˱�II:��l��1��#k:�e��}p'P��y��b*)DN�2�>�����DG����Un��eJ$��8�sV��g`�:u�Il� ����^D����q��� 0�}�l��ϣ|�P���Q�-�f�1y��^DC̵�-q�f��6�sUJ�k\ t'KԲJE��otѽ�%=Y`�&�b�I��f��������6�%^C�?ip%0���m�	��]��jS�o-�A�B"��<�óc��	f��0�[Н����:�^wQ/"���E2�8Y6>.a|�q�-�����(."b�vW�A9ęȵ�TR�A�ˬ����wH��3v��W��C�햆�t���Y6t��f�e�!�=o�7�r_Š�����F�h0�������������)�1�����$7��d��w\oz�eTB��Ʊ�nA��|gm>`�⾇>c*J�gp8 �S��!ߣ�jFt)��s��ȝw�%��$%o�0�ʌU��g�}����{��S�<w���.x�Ab���%'c�w���d�$�{�UA����<!�"�0E����#�ŏT��b�f=��1l�/&����,��!Dz}���u���>X���j҅ޅ	��V��"'�{
�����2�/�C���?T���5Шws�$.U�C�,C#x �X��Rް[��& ��@�6deu�Z�4�|`<���5��_�%��p*H�N���t�hT+�W��O)��q(?��;�;!�~}��o t�nrD>�ב9E��UY�u���@��e���,"/ɧ���)�"Lj�/D&/4l)�+�Sʰ��Ɗ��f6k"d��,�a��R�`��KO�C��=��h���|�eE��-�>R[�!'q�����@�ש%�yNAD�zga��[��VeW��x��Ӻ���a�V���|�:������C�PY'�6��Xl%zs����n�E��֊�((�A�`���?�1�����뼓��izjY!�Mg�	�P�k"H����i�2��4��BB�L��g��E�ș�	�o�3=U9cᠲ���� ������@�ȵ)N��~~����1���m3k�Z�@BX�t�s,�U�W ��!!l~�q"AW��78�?���r^qpM��(�%�x��Od�}d7!�>���x$s�e@�<i"�gF����$-|eڕ�`!���)��kRc���siO�.f�s;=tkP��� ˥�F�c 0:�j0��%��j�g�nR9n�Ϥ�����>���+a@�!���xi��A*�R�D7�"UĨ��0؛1�@�s��w���!t��2r��]��:�p�e�)���l�Y���]��]����������~��?b_��)��
��\�]%�>��l��g4�^�*���]t����	�B��Z�Sp
Wc�~T]]��vW��d3�J�3R,(����S���W�Aql@��s��Ǖ������u�g����k��-vJ"���@��(0EE�����$̺hh�"1��ã T��B�ҩfuê8�lC�fs��ls`�v�L$ּv_��$Ӌ��yC�6u�/��ݣD{T�G*��#��ݽ��]|���C�����q�d�+;�����haR궬��IPG	W�*����m�X'��|d+d����ӆē�lG��\����iɇ&�� N~ d��d�Ǟ�I�bwu��k�����/����%t&l�M�����T����H�F���e��O���Yn�Y����Z��L�3!��Sv��,'y��&��3*�*1��]�F3��q�jj����9tXa��m��+��\->k�&��Kc;���1�[���`�(n=���p�@�k�N�	U��S%$&���w���z!�{���4c%��e4f�k\:�i�XQ_�/,�js �?�&\�Gr4�'�7c�������a]$�a"�=�lS↫i������@�e�P�g\�"�o�g�s�ȒFw��]���R���d��,:������vsl���
����.O��j~���ƻ֝�N�ku���*�S('D�ūrBS_1�@�ɨf�ॵ����%�e�G��N��5K!�07G�p;�~2��Qp�B�]v,M
���
>X�Oq/YZ��kx�E�l'�C�z~��]��$A�z�>��Yi��\��?���h�e�uJ���k0�M@�yd��D@�Av3x���x#���B����;)�p]�����NK�oC��iэ
U���,�e]�P{\�#S��LI��V��X�<����}Î-R��#�O��1vP��|W$�<���T�ڶ��Ac���Hנ\$�~0O|B'�Q���b���h~���D!.���R1���tIM��lvP=����
����������-�M�n�
�Qz[�BPH�3�#�^&��5"�"~S����z3���u��a��pҥ+�D`/j�3u����=����W��nɣ᧊� � ��C�k�x���ZU5�E]p��gU������4K��zժ�:%�Y���)��!�v�*P����W���,�JAeOˆ
�V@�[�-��r��j�B��5�ٺ�5R������/�z���oֻ����Y8�Dw��/�[��lnn���TW��{\���v5z@���+`�!]B�d����k����=��엸��+�ê|�{��AQ�`-�-i��������7�?5�V�kP#��g���j�-:������4�DZ~+��R?&��{�U���=�ɛ懫�x0�g	
$ː�K�q�2��������� �8�ƣ��0}ƹV��N�>�{\OS$�c�5�Q1_g{���\~��)v��W�,�����N�����"��k�Կ���hߞ��I]����0��܍�/<���+n�[;F\1L��������:�v���B*���2���kO�����%^<`��J�4NR�*=�i�,��A'$Te,��Y�Ϝ��X�D�Kv:�謃u�:�H#�n[�Ȋ�O����d�D�eG��7
����b������&���13?�8O,U=���h��@����;\�ׅ,��Ɨ6��)NdՓs���ƕ��]�V�M@��x���a)��l���d�f�V�zOl1W�N����.����9�^��� `���X�6�+�{%�MW�����.�O�օ�� s_���jڦ����xƯ�h��QM�'ןc
g��	��%mQ�n��h�TT���f�T+%�k�h�8m����� &��x���f
�dz��xTR������u������.9[��7D��	��ēS�D��P?�H� l��h��[�o�t�3ōz_�V�/�!�
�O�zkZ������Ж�g�ܔ(z}��q�:1��qn��H���r~s X�I��;���SYK"}�I��x@\�.j\�X��D�'��MT��ҟs����1X� ��@�8E� �P	k`k�i�Ъ��"R����mm~��fc��3?L�&R�� �S��*)�`�������	��S�P�R#{ES�5D�~��$�1��|"S�̭_�앯),�<Rї�:%Ce0��| �)���2�pX��ZWo�@�#�;�����{$BvHAɒ��W2<@�f�q����hl�� ֬:<�@v������Y�}	�p1f	��&��f�i�絋~�-��*��N��7�v��^���-V�mtt�8��2��U��v�szZ��L|�=.�V;���R#���~@~(�nl�LU��7���k� ���c930��T(��Q�\�_��[F����4�|����0+`�Μ�uIdH��r���_�FǡтN�=M��nbnb[�b����0��W��<�v�Oz�8�e�R�R�p���>�V�B�e*9 ?ﮗ��k�$�X�rTP���%���ʨ@��̎s�g�!;��.�"i�����v��QҼ��6��R��ؓ�p���O�)�$I��v@��H�wT�F!���Y:�ds��׆� �k��5��_�;��t�$Sve�]��Vo_%(oL����,���A����[|y�Y"�zL[�K)�̼L��%��Q� s\���]z���^g�w�bP��9�]���%l�����XD5�&z�Ԧ�p��h���y��4��Zy����B1^��G]�,]it>H=}: ?n�cP�Bp=fu��3�����J�����NݚT��,���D�4B�
ہll
�ࡸ��r��s�4l1?�o�7�;���c���h��̡b�������Y�L۴}hC<L=�D ?�L+^W=���\c���E�d,	�=�D#��N�մwT���R$��^���i�T?�Ĳ�T�B��m�ZcGnb��V1������B�����g�AəX$��j8���B���L=��e~���Gu��Ǖ��C; 23�ڟ���z��]}횘<YJ��L�b\��b���G���'^x�{�"3Z��q���s�1�	L����&�y&|��0�љ�k�$���yQK֯,�L�7Y��"џ0^�^���>-�feH���H�N�1HX��+�~>	q$��t�x���!*#ɹwJ�U��hGV�=�Ǿ��Hfe!�Q6�,a`�X�e�俯���
A���8��=�m��}c��&�}����7P�z��ܘ_���r��h��b�a֏8��7v�*��$Sř���B�l��d�.c��K�\�j�׎[_�D��Y{���@�BCn%��x+������rX&�}ɓ�����Y��,D�Kv/`����s�I���{��k�s[�1�;���;z��i�l���r���LJA; �Rd劀$�ZP]�x���ڦ���C�ֹU��� ��@HGy�a���S�_��h��#{�Bb�q�jT:AxJ54�XML�\��g��5wZ��12���~��ˮ�2{:ZN�D׳�L���7S��XG ��l=�E^�8��Z&�'��Ǻ����j��3��Ք��C0,�̐���<ֽhD�:�ܤ��kT����lK�n�P�ev��r�\�^�=��Q!�]��=O�F��t���QP �{�Me�+���~R��FɪX1,^�E�F�z��;0dZ��֯�(Ho�K��t���3a :�9���( :�1�g��)uT-�^�R6+���]����<�(!���8���9��0X�Y,�@*�P�5����o����8����,�q.�Ȧ"�^oM>;S�ll�\/m�%�v�l�qXB��m\^���o�3B'���U�]fG��)՝�����`�[ؚ
��]ßv֑>�hH)�{s��Mf�:�6�e���Z���^ �A�*b�s�;k;�d�wPP�!-:c-X�B _]7ֺ�� ����X���@�*��n������U���a��]D�? "��:�÷bPI�X-���4�a������)۸����$�X1�,jL�e^�x�s���eVpiX'���/w�;����cY�ʧeN���G~Լ�pYY�u�W�=�VeA*hV%��W�{�s�*J�^+�H�k�Gʠ�4�1U��:~hUMX�;5L�L�#�!Z͵[P�s{dԦkZ%ӆ2>�H�3uE��$*�w�eclD5w+�<W���������8z��/c�J��f��H�W(�Z�-���������r&��4H�QB~oR�y.	р�&����w�����ns����kv�AD�S�5zr�[���$#����yQv��	���.���vP�+&n��xU�g��B�L��\�����z`�1���B]ll%'ƨ��L�H�X\T;��?)��$:��$_h[�g�'<�Q��?��s�k߱��+� 'x�6�JA�py�#%�$���J��h)�ǲ�OY�1z ���߁	�w��9�:����WEɁR�-e{�J.�_����<�˳ܬ��B�E0>x5����_�#"�LW�璘{�/RR��L��~N'���+�(�(f�ߦI�����j^[�F�A�'�>5�<��ݫ�'��Y8^{�$�x�|�x�Э('�(����lD��K�r1������~;��t�*BP;ؽ@ǥ�M�Mi��*%�S��L�ИDCI��%^۪m�I�B�����ٸq�5��԰���؄���F���+Xƍ��Rf���P�r7��4����y����t�����?qm�I:�� ��d����:���ڌ��w /�m���f���he4YV�jK�,��p��Q:pd��4c��̼a��J�-������30��v�z���m�L֖� ��`�62�k
��T3Ψ7VJ��P0l(.�}��;g�8��_�m��~֕�x�F�y�h���a������7���/o��1��B)�Mk筇**�H�ˠ���G3�5o�V*?
�G3#C��*�| x���/���y���٪>i�oQY�� ���
;���4o�2��V�_�R�h�I����j�0\}��/Iߞ��S=��| H��i��<#�>5���]�1FӖ*Th��V���V�ܠ~����U|�ӝv�f�D��S9&J-H�M��j�ؒь�L���G[�>>��E{����
3��	����/���
ԕ@�[��)0��C���@HaS�m���?	��j�s4���d1U$���ȃ�&2��k��u�z��i¬\yE c�6�;����sk�e���'|�6�x|�<Ȃ�VĄ���bBԠ��i��^�(F�ߌ;�}՗� {�w/D�Jj�,A�@�{�ux�wiN�M����li9������5/�5某���p%�d<��lo#��wfǋR�!;�U��B�*���-��^`�t)�Z�I�я-�S�@-'�sp�\�D�X�݆ �O[d[5mՔ���	�����J9�H	����m��&��W!��AA��֯�D�!�:�s��Ԁ�tTL|���x5U�P��C�����t΄����s��1IU~.��� ����"�7�r��9(On�B�BGi���ý�����$� g��3��;���e�ȵ�y7Ј5F�7��U��2�2��d�m-��`%`��_�%��ze��HT�~6��2#gP$ދ[e�U5�>��<<�
#d���>2���էq�O������#�J�k?�,��������1�jo��F��X���;���J]�רn[��q�Q���\]��Θf��|._�4`)��We�N�3�Y��h��ԏT�4�;�`C1m�; d.H�Zbr�FHK���.�<����+�驚%4_��8X��(��Ę���A�"'��A�z2����YZ,ʓ��$���P���Y	��K�AK��Q5�f|mFƧ÷[5�>���*w�P�c޼�X�w�2��N%Q��4s1S����^���W*�1��A�>�!��N�]J�����h������{lMi�kd��w�U��.�®.M���ʵ�pQ�5Bq]�4��=��T��ǜ���`AuW^�88�|��i�4�p��}K��??�<&t�*<T9�b���ѲK��w塷�g�t16�*����[�����9�-���L�Z�*�J���0��%���֪��K�i�:�������2�pL�N�>�,o�	�[���&kY�qO�b*���| ��yxYz�ج)7ֲ	��A% �=�����	���5��Ĩޠ��[}<����NC3ʙL	!�,��e�
�W2�<Ub0x�J�Z@R�{��<������l^��-й���N������58ud���Ϳi�f���)�5i1 �����@�����yI�#HA6Β%���m�%�\��֣�S�|��SN���[�f�*)7�0^`ፈ��	A�U�	�BCw�m�F'P��e�s~����3���-
1g*��Y�ƪc#i�:œ���FY� �O��-����7F�R;$G7��N�n�6$�"r��������o�N-Vᑪ�|��]��D�Dr�~Wq������U���(0�<����5���� ]�V�+!�c�^�4{�R떢(WgV����.�c�������ξ��p�4��.�q���b�� �f��7=@�0��\-�Ɍ�"�`��� ����i�B'�������=ld?z9�����q��Kybf�xzc}9W�"md��'�d�9knYRe�u�1f�� �_�'�P��ծ@E���I����JOt�!+���?PD�(�X��Ni��֜�f�B��|���3}7��Bd�'��w�.x)�[X^F��b�͢����5кn��On����M"�-N$_L�
�`��Oܦ��W�K�v�^lii<��Z��H&���Ao���c��Ş'� ���(7�;�L��>��9�xQ���dl�	KAQ�ߘ����޽�E[�ɝ��5P�$V���r켆��R�-�Z�|�����\�&&\��LJ�:�S�j<�/�^ �ɩCv�.��r�bHCXs5zՎ�J�湚se{��_DU�r�L灡Ϥe�:O�?���6��;w+5^�dH�%�=�+e$�~"����H�QIVtỲ�v;�X\�'��C:�]�d&��&��O ƈ��v�����_YY�~x�pTd;�oe\��G^�m��p��;y�9\�	��^v���	0�u������Cx$'�{����3��#�LQ�������?��f���Q�_F+���Z� ��TKU.ل��d5��2yԓCʻç�����c���V>4�Ï4���xP��(ݖ����s��XA7d Ik l刟�ϻ9R����4�[/��}SY4Șz>Z�0�g5L�����`O�k���!��`��w�L &�g�'�0���0}����d�V�G�^'سĤ�|۔eۧ�,f��eSF�#V�/{U�l�_m2��Y˂�^e-'�����������i=�Ueέ�6�%����Z�����B��K���&��y�|~��T�����Ha� ��A5�
�ܟ[��Ze��D�Sm��'ل@�}�*��E ��|�0�un"+:O��mv�O��ڷsT!"ؔpR�����m���������]P���gܚ�W�b��i�i�(h1��KO\)�.������N���_Ԫ�������~
5F�P����a:���,����"�Fr��A��T�_ �k\�Ph�ۉ:[��Cd�z���:�L<���q2�Ty�K�_w>��J�_��ך��?��I��3#��kt�i���K�6�B�]��/�Q45t���S�h�e��l5�ٓ����꼠���HV7�n�A#]u;�j6��ڧKyYe����%�l��L)�[J�v���{a�a6`McV�Ԧ�f2�R����)!s�/�Uc�~it��C�|��Y� /x�{�Ҏgo�{��{l��a���%P"��t�sʍp|p� �7^ϭ�g��b��<:��~w�0Y�uTf��hߤ�uxʃ������&�߁:���@��d�߿���U*D���d�M4��օ�6�uh�@�(sLX=^P��Y_ƈ?�~�ncy��S���D�a������^:c�5\������i�܎�uZ�Y�<�9$�WL������QGa5��Re��⯊�'5�O	H��$W<v���ּ��v�|����Vا���Ec���#~��M�+#i��wVKl�"��	�tdL��5vǽVVIh��5Nn B�@9�]��;���A�'i�>#��Z�^�\32�(nQ1B|m�� t3#�h%@�t@P�f7�ݳ��e�|�k!1޲}3��R��둢��n�G�,�Y֌�v2�_!�i�\2t����]-���L�0�]�>S�.&Ɠ��x��U�$s���R6=�B�iB"�Ab!^�=b�W��X��{�D� 1��.ʖԉ<P�V=��o��W+�|'"���5���}\)�
�����x�o�f�L�Z�P`�	��D:��BJ|��7��,e;�.����F�%�&-f�\w���za; ��S&~�����(��}W�`T���3K Ki�����YFru�y��A�$�8�`������C���	�Yu�@�6��^مPƽX`��b��Q`2	(辥С@as���<�F]Hz�� �ݕoh�b��qЅ5FP�1V�X��`�V�a% �e��yx�?u#���"�{YgB����DSc��he�T�ZL�`���t5yׁ�9.o��U�qh��_�[�q(X!��-]R��1>M�ѕ<�����r]�q8�֋��d��o
��,}�+�U�Q��&�o�[y��Z��p�`����7W�p�&���|{�D�=R��O֋z��]�X��{�vh:���p]_0,��|���b��.�@`��g��CWk;���>4���c'�F��3%	� YP�r.����ǵU*Xl=�u(���k�KT��@R6��rd��簋pJH9�+`�"F'��^,��;�~��U�]\���h������l�����ҷ�o���a��|�=�Ők\���,V@�����0�#ɲ�)�/|8��bR����nhn���:��Tl�����A�R��ZߚXo|$xf��7""�s�L�>E� ���I�}`�_D�M0�f&XT ]��FMЃ�K���aQ�/����w=]�@r�qJ#'���o%s��ĉ_'�������\}����\Ƞ���b\��Z��{)��<q~� ����S�h�'t�ض!�lu@R�4
��ʘr�ڡ=���Z��x���6�w�s_�k,���Pl��>(�?5�;3E{]��u;�z�!��Qyݽ4��� �ϊM+���b�o��d�ꏬ&ķ�eQ��E�n�M��t@o��%�-��$�@k� ��ܡR�ˌ��Dn�@S�Ș�g��9��=�)z���Ux�/��B^k:��v�')��k*��f1V~�G�
X�Uj?�	:U|BJ�N)aWg��fQ�x�cA��&S.j�m�;�oC@g@��?�A>>ҮN5�/t'Z.ڀ0����tV��
���#m)_0��:��B��۪�H(1�!��4�J����Њ���e���:a�.��(�5��.��2�y�d�N^�#�"�2������P�ƙ�A����9�����eB-��@[oӮ�!�N4$��:�N?ײh�ZGe��	�(^g�T�����Ey�
/U��ƅ��o ,�c�H��V[��a�"���|�DG�W^��e���jb$�^D	Q6�:A��n�T�.k+��K�1�x�PQr�Q~j��hPס��6�p8x��#&D�_t1�,@��G;E��@Bz6�^�g���~.^�����4:�zk⦜9L�/�7p�~��;���Ĝa����g'�-Oh��w��V%��	o��n�\��7���ɕ#��LCb�s=��/â�~lP����sh���J�������)�ҶC��׋�3f
���+(���0��=*10ˌ�>T��=B��D�%ڬ��?x3�4)$�KĂ��5�	���n�U��}m�N����#��x\��/N�):0�l���]�;Fm�A-l8�M{؎ u v�P�'7�%Сgډ�;zc���n��p&�I� ��@��h�'z�p<E�|[x������>�:8$yO���C�ƇZ���\�Q��T��gz�		i��a���LeXsL��������ۗf���N1D滿�~�_@֥̅��tvUC��G�`��V3N@:+p, ��&�ReQ*�)��GJ�|�E����^k84	�m�0��}���ðtf2���w�@�f�D�S�*��s�'����b��z�@G��왡�|�˩��2$^�6�����s6�*���W���b�&9ڸ	�a:�l�����x��8|������w��]�})<�yd���z�(	��y\\㫳�����bG>���/7��	b��S��%��#�.��f�=A��k��}�U'�7���  ��Q!�qw_^C�������a��NvVgֳӓ�3�wF0R��m�$i�>�rj�_%�R�����`���&��w��]�vND{jcPv#)�
8��������>?.fK�+&��p��q�Z�w%���,~�$һ�ʩ�f��;;���f�1�t�9-eKkܾ a���]12�@������;c99�c��[h�d#�q�Q��l���t�خy�ֆ��D�5A�OT�>�}3�ph�3�~g���� fy�wm����t$�"� G�nvJ���/�'AJ�[l_0���b+]���I�����Lb.#\c��Z��b1��ܝE)x����c��o��cBr��\��*�o$�l�Hޢц�(�m2�������[��أ�~���o�N���C�����LǨƇSTx�u����<�Dg��ؕZ{�eB�e�����{
�������Fߌ�ӿ��������l����5��qƈ�9Ku�;ғ�e��A��i�7o��&�
2���蚇���{�
��]]�^�����4uD����� ����<����1,|@޴���,XI���4Bĸ�c��.�e&P�]�KO��+~mqd����9d>����wVx�g_a#�^���aN3�Pf�}�q�W�Wy�?\�3��@��l"���hC��T~V�k�Qs�h�}�[��֗N8�[�j(E���E��*��� k1Ag���>*K�Ԯ]�D|u���K@�s�<ޠG6��fE<
a!;�|ϭ�4�9���1����i�b�
��Î���b��8�W���)��W��)��v
u�t��IK"lU��������P���@0V2�}�ئ�c�ם�㱥���Y�5�j_�j3+N�	��)g�HQ��"s�>R���-:����E��+�z��^܀s_���� �T���u�����&��2�I��d�t��)I�.G�� �ơR�� mL�8���J	O9j�W�ݚ�أt#�}w������Wkҡq�����η�{	aZ&v�wZ�CJ*��@��:l�Vf����
�4p ��n�'��b%c�&�����Ƴ��ݻ���Q2~+����'�υ��w�=�i}-�hhI��WH� ���_�1 E���K~bW(Cx�(���~��g~����S'���ݩɎ�6R��K���B�P:3�
�����g�ѥ(<Xj^tNI��v�{������՝S��٨b>ka&`�3��
���!��
tXM������?T V"�8�]�fr�]%���ۃ$�NQ]���Z�.����0ۃ�k�����I�{a}�-�5.���_Qؓ	g�� |��;5}Ny�mS�oK��߯`�;�A_�E��7�w��ZI����# �����������EP~�::���}�!ya��;���'�8R�>�x4	y�xu��S�O�\pa�K�������'�N���5
�i�Er�W�N翜y��zh��0��Wr.��!|�=q����������AD��Htb��	�\��Ʈ�a5�{d�^(rVK0Ƥ(�$��	5��G�I�	�����Ac�G���� �1.��s��6�½��#2!!��nu1b�v�*�f�A[����TV�A��ھ5J��ʻ�{T ��2�8x��d��8��I޹A!��� ��6l7�}�-��չ��RIT�󐠇�M������F�}"Ժ�!Aj�KR~�Liܒs�� �C|E9t�qs6T;I^���
��������B�|#���g~s����I)m^_lf��S#�A����^��,_~���]ǿ��ܥ���r��!P'