`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rtv30VufWkxfO/pygHOGpgCh8BIQgDOxlRBzMr28YFEJnQ6Q8/m+IxhBmitZvyyC
Z5V24y1esbWQGWg1VSDbHwqOyNuoxAzOQpnEK2lSKLhiTk+CAGeN1RtPSODLxKEO
XJB7wgHhRlBKabZEOR6+2rMd/RtD/oM5J8zmFmmKIbo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43776)
6fz7jNohxlZSGRzLTzrW/27riU/82NSVp9bfUWqgA4KmTs/OWReHOoG5bIdJqHRd
rDYSElh//qxFf4xEOlYDOJK5sVzi8T5OhLPdKPLQG9aKOuaCWDUMNL2VyHCdi0QF
TDwQ3IOoKIedCEuI9hku6D0yKeqW+jHQawDAti57S/V2PavxErIN534n1ugQMQ/0
BTsNHJR5ST3CU9lHBk8iz4m/vcKVWIvVu1+O8YhdjGoWvE6cJQgTz1nRJMA1obqn
tvgMjnfvkBMOvSqMQIQgrQ11X8QF7zA84aT/nEg0h6na04aLgx7CLfaJ1OfY8nue
cub+pazpipmMGFG6ZyIKoiob9t7Cag83AmZ5AUtCK+Jo8lSsd5GRnBepronyETO4
xWVSNFEpm0Y4J/B2jKHpl+EsyW/cPqfh73HhGpGLfyHJhYG4oiK+XSsdJ2CRmy3O
YikhK1GxdQVDZv9MVYLFN9a2H/yF7OFa98AOSsptjFPl9PPcfQfq+5O/hkHbjGty
YcssIVB0h2OA0f5GZ5IROpmhxCFXWGSpW9A7j2D0tjyNiuUC3ua/1ta0S854aRKp
MfXVRE4K/eeq8wJPV8Gpd0p3InIglRTk/J767RUjQbGvU4aJeqFtlDyCtqOuU5vd
OjL4UwM4XwbAED/eb6shNvC/SdsYxrBZ5Slp/mT2e2c1L9YRFexiFCjdzgEyeQ1F
9M7Kk3zMcLlHEMbK3G67ySKQv8r58xQvnsNq9QQJwYgbdBl3VlAqlj1nKLr3bj58
2GjNsgZN0MKADpuoss8E8BHAdt2D5sXLw1zSBt3CqIGwrEtSD6afwQ7HfBvV1t7n
kU2s4bcSX7Rmmq5nSIs11pk6LusxoEy/ptWi4qCb+hI8Sy8tN39c8GqGI2we0CS8
a3tavEMgjbUQ8YxM24Wu5CVXGO+IMYhOqqxU+wUisrWPMLvzYdYneLNYP48ErLRb
NJapKy+y2sv66+1xUjCM7570tiikQtUxe61jN08l9LLdhxzP/zDeeec5szCr1mlK
ZiSeSWdE3Ugz3xBsY4JrZlbVtPU+16mnWC8SfObRtFVQVUSPLJFkZmemD1zNc8/f
9++vTmD0pVCzhc1+idslfeEw0o9eHzYWjY/LK+orOlmtCTStmhWqFzjPub3Gyul2
iT8AGgA0JGCDiAzXTDtdXkQbd7+QkdSwhm3HR/PYpb1uoj4++1GDDG7jjb/cBWe2
WX8OvTwhIXlOKB3Uc+LelWuQGkMMgyCoPmUfbO6bT4tlqB6cWgQFFkG9ybcMFVfA
iCN/RHPWYQFfyet5o3SmHnhopt6+zshX3lL/jsjUj3DpKg5dyo5CF+NMdhw3/OYS
OMRO2yQa2pkpQprYA5iuO5cs3z5xRNrAmZqfOF4mYwAqVQ5Sbz0NTWNhxu/UkI1I
8R5HY5rihXmiRTC2IfRT6qgZCeN1H2UyvIUeoothSFO6egIiS4do8JBNHGGnjdFp
LAKg0vDc00mLWbMz4aGwG8mC7wbFTcQQlKFjLJcBc2eN/WVbFa46bQKzCaG6bwmD
U5aG/OrRTBZ+Puh26zThJNJzMJ+ijOudXh3GYs4FaRrv7knnp1WvzwVL/74WQClV
3QI7kNHVBfviGoJpZqi7FnjuRXd7kbEXrq+wgl24DCnCRvZ/DIDCmMTYKGUhIuNK
oOEv8m+BlAyHx0Jtrl/NU6ADX2QxfpXjPKilSuMoFo8pj2n4vqX7lRVrlJt/OFXZ
HtImBCzg3qIIaVWxrasadHemARePlzimuOuWAGsyC3YrAjAmG8Gm4peHI8AD4zLe
vw9y2AmKzOByqvH/udB91HZ9Zn8V5TEXX6wOCXqCWTjNq6kzObTDcDc47XcjwHjF
mqnRi6Fiq59mXKACl6pa5LuDgEHt99w60FFrCSLE/m/sulq/rOaCcywU/2K0P3gh
/yRwuRPR0Nw0H5wyowpNrrqcOm4It8RBhp6C8O7yEd+lIZMrhWCCoZoBaLHSOlNJ
sXk3dJtXFoRrQ9b9isSRc5nS++yMwtMNsfLbKBr296DZjwP3DK+6l/j9LdsxSgWX
yVe8ZvgMRM/FI8UrzMjAwb9wnJUMbV8jnV23Qah81Dh2ZaD7sDOnjzWby39YxaFE
JR1p7R5FEyclJfvDoZ0SG7HLkRP5uLtyCQkTjr2ePtUoEbVlANp54yWQKl7EAlQ1
ySQoTfPxDSj3U/zTGaTZPH/TnbqujisWjgkWDxXmONmM938CVTxONdO4lRtd8NOO
e30MgfhZQxT6440CyBMdB6wN/9KysLocTs2LExfINf+agFqp5T9Lgsvm0fRxg4Jh
qJB3xRRsERiamctuX/Uebr1sGzly0N9c6sb9Dcpp9q/aG0HCrkmyYV7y0Nhhg6BR
6UyUP65w8snvFsEgu6Bj0C4I2FGKZyNNKx3jMGCG9J4oiewQ29u0tkxkFfKiLFc8
2+0h1BbNfUxfz05MWBRsUpG7md+LIQEwVu8xDSYxq+dIQ1bsiqJ9tMNp7HB2i1c7
p+ScXlxcb8o4CYpGcv2hEjYm7tQFgJbDbWOs+OL5B35tWHblP0sHOIey6f8T81K6
GGB2lNl8yTLV4sRzfsCBoqo/C2a03fIik1l3o2NZSwi8ZqkGzMyvgEBEKRjWwkFh
g/ZG3mpRoFs/SuU9A9nlMR2Wizlx+wsZAUGHdjQf3o9OqOTZmm+v+XW3VQP4Jfsj
JrEglKsnTrpTdeho4SyIz2j2QxS2GcgjigUbuu+KzxLQxMEymgu8ib4rpWNAIXn6
qWWTf0QsRDlGgJn4qw26Sa7xE9osSIP/5CuUAsnxM/DO2bKFdP0kSgRNf3zm6Ses
h7frNf52ghCur4Mkj7iBpipsCf28RFwqGReLeDEK+tHqiUqzJPmK1iQpU184klo6
UutMV9PBLAGnNuiC3SXYn59WlYN+73y8mseESIq9fS7tZWcsZ4fXFadnDouXR4r1
XAeThEwSxum6sTwN1+Yhcg+2GtQk8u8YzefWOL1LPXfRzNBPIgIyHoJlhs6MHSRj
jqxbpSsJY2g73fL26hXn5tupEphwv+2htMoOTJ0VPnx4ZJUHz5V1hLeB6V3BC0G5
yacz/kDTbfg5nHAMyRgvZYLBf4u3BJFhAVY6dD7ODcWu5aczGQJrmShfVw8CMIjz
oCrU8BcyJ3YSlYRd1vd/c10zEYhZI936dhGmQAqN5+XeZ8cDzfb9iv3g1LRuKaZ1
asqXLeqLU2g9lbA2cUPhA28yU+8/P9yGFmSyVT21GYoXTXXpJczk35PxNt0gubUn
IvAEVqCokWtP467MCO46dxJBiOHY/MEo5xIUd6EKrvIglmKO7iKdz/I0roHM/4VW
/DQL1LLrTBR9xVprthAzKGkkxKuI1MfLxau1MC2u0C/4SxaJS5R1ktMmcL9PR5FH
dlTAVqQYED6X3DpKlZ1/VMlNGL2cRcu+y+BpIXdI7TQS7QXtxFxwoc0KZVkkUZ3g
1msX+gl/JWJ75aj8NFRcgPSJIVAASJuVbuH1pmlHPy7OBDkm2uHRbu1VF1DNIY23
JwhhF5NK+n/c6O4IVyf2Wl/uwW1xK5uWSq+i3PEPesmgubOP1JUkEVaXufLvz6jm
sj8tgyjAX671mE/Q0pczzFUC8RiTjD3eiMvuQkYqiaRsGBbfOIzCDlWZXaj7TXLT
3ivpxzzb6ku7sZ4AgYTuzbP0nwiXvZ8+ECP8Or+Zie+iHTXa4EN0D9juCmyGsuM4
bCO03WhHkvgLqL6K/DPXh//Ke3ZuwsLD0NxwUju6TQA49179RWb2ZWlpjzBxEKsk
i0T4Jg9/xI2+2Rv2BjFOcYTda3/T6uLzQ9WW6XrcxymJ9wS/1/FnOxyxfmvcVgDL
VMJBDJMv1YrUj4wO2qUFlzqNe1FoY5oQ787193qJn+A5luQqhUG6wJDYDEe+FGF8
+ZHKiQudusmm8inGXxEAsZeHYNrVseVycZ2viVtU+DjL+4Pt0yZ2p9UqYamLAgRu
ALOH6PDLFK6gvWNTgKyuXxF6H3IP9gS4fET+YTMAouVsZM5lcKw1JXNf0Xs7GMD+
DVasQn9NFcIRv0/W209jat1s5qc/4nxw36x0ANlnIhsADd0QAwybIEtTl8DsrFcz
vobjAmh0OOK3vfEYavEu8uIlt24k5ANYPPc3qmFxESMm41dNrFNBJo9ZTbD/95vB
QMp862d5620g5MbBnGHF5FM566erg4fN4+BlHCzxQTwKgvgYFjHeLi7gYFazMN9f
ghTo2OkP+iep5r02lukhweRLDp6NwL76YMTD74tl3lTfhln827L1mf2U2EJiJ04o
axrl0fVaYIs4wT0q9TFCY7bfvxGd31JCSW6eEydNAc0ArXa0fl26ZboUhg85RP9D
BUBXbUjdr64NqEnICz+1ijy3rrXMBILKpOQ95xVbG8p3c+9RqQUafTwy+rXNYwoc
SqWGZlD5u2D5MhmxTWwx9abPFrcn0gFV948A5wSZv2xwy06RXD/ljMQmW9Tcq2KO
NRP7BkoB7dL+DZVQT1OgYt+/xTDDv3xXF4DyV9jXEYyNIVNwqL5PWlgFrbL8fnol
ZOkl23osvNoiWckhsCjJnEzWyT4NDGa997YnnZU/QjK8/pOUyQakqAmfumqAdMZT
FpX6DhHdHy76+zE8RPr29jpy2qh4bW98IBMGor0r9tcC6HSInKhkinsTb5tFdRXv
3w08B7q+Vv+DBn/I7tJYvOe035lPRh9HkjuUfNuxTo+nEcbE7Ujd/SPi53m0JxS9
0uf70Qk0IoEP4XjnfpHQVaX/HDpNI0jGPMP6CD1qggWVc5QRmE6X+W5QO63ex766
N210v8IY9xG7nUSXXQA4lNRk+McHeShp/byV8pDqRH8Hy9hZgVqWNQMuFxxBpst1
ezCnN72m9qXz1VgZN5Q/Cilo7WGj9NlTO4mScBdr+NiXCNi+cEOKbQO46mcCSk7q
BzJ4crDKJty90Ai2+YLUE4sinqVQOzzpKtofTrmN5wYr1DJ6EUSw9y/H6Ke2FjAc
TIBAKmRZWetSNSlBEiEXEQbC0MhV8h+9JNHS4lrvQnjy9gmC00S69m1bd8qhgxEh
26oaaQt9Wh3wLO8u8YKxd6xN0bCG3HAY9MIgqTw5AixwgrZBPO1+NEH2MfjX1+Y5
TfANPAuzDPVhiv8mDfixP2Bt5n5ZZILRAYV6/5rJPKxyZHYzUXzY1vaS0cmdD3eD
0XkSrdLpJnB2m0O8rAkEDH/b05MKH7dte5iFwLD3vV469X22bu4L2BhZ8nVbSzvC
R0lBZRY0IYjDonvHLkoODtFLxFOMqg5KG7i2EUhzZQIu0sNvWN5GgBWlV22jf5V9
NPGUCrbLQFKen1EYDJF1jNC5jiAvT49i3ytR4sz8e5faIDW6LORMctwb+mE/1ORP
5ehNFyyzX1uQnHEttjm7jOrlpmBQekuMDPhRRtYTrA6rxGwcREO4PkocBA/u/YyY
cWxSzJ5XKqUriA3nrm508Jdij6EHMvaLVpr8DMdon+8jDYYVoDneIhKa4frOVmbq
5BMorXQGS0Y7x4r7L5z/jmkqeTC9WAASYth9qo/CzvpOJSu2JC42/1Fq/4W5wF3u
Iom7HtE+UJo8cqWwnGU4GopLPoC1ZARSUkVVJbXDocT7ddWr89fi07x21nvOpiel
A3gPY0TS1lvXL8ZK5bYf1p/ezSA83n5BYEIoNp/lUZ8z+DTCc11NDpXrBPOW5FJa
7cZE+k6SouQ4MfyhOXndZcMwf99KyLZP3j93qXJ3IsfJB/vPntunb/2VoM/Di0iR
FlcF5Lv7dmHHIKmzkZVDI4MFqT7auDN38pNhUJIMmShfr/QHNDpo/D40FeCdpzfj
5wWs+b1V9HHveYia3vnDYIqnm/blNvbIOI4yiEzi0eVyCi9ncgYyhhjYtkstGSsH
rw+HcP5SGiciRACip1KeXSDFpkLCSqGSDFIQp6MRyP5cpKO9vrjwp00UNXTkw6QR
jOMW3QFasXM/WV5IbtqTLHBwVSFGMftm1pkDGGjIB5sOKvIFQcTUXQyBlWPkFx8L
IrN6PnIpZGkk5q/VCW0tB016PO1fvPxf2R8mJb8bJfXxSQD4bOZmLGYHTghchawY
akvOVXfS4hbMje1lnu/lc9NsFjNNrX4HEHW5QDsbL/E/IhIZcRQiv7h5RhHeF9Dg
r/M4O3SzZdSLxcP+7ix0D6a4PgGjs1ZhKgc6BezE2iHEf9oop/2cEPSL50FS8rky
0qaC55gKphNKrtDSMiKO4PQg4f62d18C6f8ljyMSqeVDmSzGWpZYyH/VUBd2jc3B
6VKSsz1boFLG90h7tGCws0cSVAHyXSO6FKyIj+M/msUcNdQGtI5/yLtv973bdktN
NnkBgmOrNvQ9tcLW3M3VQA1DRlbOPx67OdL3HiJLhIfC10BDaCiYDvIeLmOfocAy
zE8B5dNgDGa5Nr9Cdu4rME9tXZ2IA6A89sXFrSpIXg6I6W8C0TCQoogB3bEzntSM
J8R1W47F4jjgvmtCio9L8AFS0RRFyM/bgAjAzp3K5YOQhIw82E+nZGc1QxpVkXiL
ccwJBV1kRiLe5xK1YTz48i4DYQJcfAjkVKyn1OVJ0zsZRGRZos38RkB8w6iq7MrL
wPPNaHRZxS6XQ43//cPM/94N1y4JND5q0I88/MRwjhNlwjOfT650tnT2CCDxVN0v
PvdbfWNCbhBGwwavCsbtf32O+I3p9ZX9cZ6Ncj51lbmJHc6gp57ZppGtKGCMjhN0
N49JIlb3dUDqCwx5xRm4a8M9XesICwIgMSwEo52KgBvXlzQEQ1yrNncZz4V4uvMN
uOxOskOs6y7H9P1pz8HgaF7M5gsgg7RV+3WJKXYZ6f8ytW30318PjUnz9UyMiKDx
h9kQmWOFeD4Viro4S2aJN2kuM3/+lrNJqdnaP90uxViPi5Gc/lacdh1P7XKr+tcS
w/90lOu8fq/KmLEbS+JryyeHQSxYWQcfsVwXxREcYpnoKiSAHJwX8n+FlI8Vudxs
GfT75qDydMymPB9B8mXS0wqzol2RJDY2KuNawzgUCM3nN/9UH2bKed4GP/ZBWrJ5
zsRRtbhKCFesTE5OOg3HeQL2y4S9FWCmAUe+bdGOmgrAP0I7DfycxLlPa2M27Bco
jsC+UDnkBsAI6UjAmXZFSkKaCIv9RrQreNdYtGZptHJYpP9uHJwyfO130L/i2pty
dP+8zyhxivd7MaScSgj5Qwobel9qwyeYuDjbn/Rz3CCbpTmPAtmQw3QvqjbX9s3X
oucIzYXLAwt3pIpvRpZTQwF79ZBNRLgjP5Vnjx+cfXQaWQ6fBZx241kp/h/cEjgm
lptYe1DyquSIU34xDS1L4qasYMuKQlniiKXM8l6GmEUM+Ij/Sk+7aoztll2IxTXg
KBbsT2HLq305wmBtkEMlO0qvnQkPfEeettLQ9o2pNoLqkZMDM1Ppp8Ld+EhARGjZ
yrvoF+eQFrGEuZR7njy4usFkMh18JijYpAh930wDLaip2Cefv4Ew+EYYt0LtrONW
XvP7/63QzcIhPuXVQ7yCuQfxeJO4ReQsQob4giGaMtiUUnFyswscTA7gxJSKJrVD
4NyeDaHS3MuJCOxx0jZiaAxhMbb5IT1HhkrMrgFxIB1UMj1XFr5S5EkVt9gmqB8U
+Hqo1kw48Jg/yokRVztgas/w1DV5058FkYgvYatNJvsgjSOqiLOFpMVp7Rr1m+lr
Fv0FLNLfY5szLSB0KvIicTg5AjOYgpTeWqJ5VAzcYNoBDYtJEN7sgasxXj6V+bkv
OC65nRwH3FyDqIzB9cUh0gtLTFVWtEnkf/s9SrhEz1/n7dw8sD+0Xv72D7YzjYdI
aP7GJbayJWZqxXwxWixeOmD/4MyfNyBsKM0+ENZAEpky/C0Q6F7gP0+GfNW1Lafn
wfp5PfjTe9yxwjD9YDFTvLkhNSaFiped5JESxYXqF35T9bWcJ+zIn42h9r+wyWwo
qm6CFVCUJ1vrKsQZ6nYP2wZfU8ym90ayxCQeD+xfvJT42KxtjD7wVgo/My/chGr9
pkmwROADY3caUPLo+CZX1KDNj7y3l1lccMriT31QfjGVcIoKYy6yq67dcfk8MC/z
4F+MycyAc467yRuexEP7kCE5D/sbdvytVAJ83I4kw4/Mdo+4hTBnITmf+YZRHMRG
Emt4E7QaSJzx9bxyL+YHBPvxqinPSSrkIljXOY+eZbAf3rGhGB+pSBHTBHXK53NX
FqdbuVTfv/eTc3Becye2w419NUpCFcZtVQgFzdoH8MGzIEMfjErqxaG50djIiVK2
1g0E3XCif35NjdXQ39CwayGjNuw7LHrpbj47NuaEEgFM3hQoVBZ1n+2vxs6CXJ4z
x+D7LdA4aZYOT8YSKadVWkw0+CeanJfvtN3W3Mm58QqZ5D8EXZWbb6KFvVaAFr5K
DpIe78v4NZF9A4PmAVV4ktuhPunwnOZXIiGxabJlWMCgmyEmXSbKKnb+sxoborVn
r71aWdXJ4PIRiGuXqjm2d3JrI2PKJETaiLtTUrlXSZtL/DZfDw1lAGnlEF3EdhQM
iIztvtzqfXyKLPTRVyAbYs51FHxpblPmezMTRuqzZKVJNRIyFMGvOzSrLs3DyK4P
rJxOWacvY6DGZupVtLvvCv1vMVeMsRchcJYrocwF5nn7VVM7yan/Wa5h4AwqGrlt
CPiQiB+YZuzj6vkuM3DWZjK/7gHAQ36YZnVIR6rfZbFj0qKZlsTxFp2P6Itp6F/a
ZiJMhdW/QuWUrxso17vgm/KuNlQiChpzGHow17rxnAFVWU0DNYof6/lJcseD2iGA
LUgFT5Cd91vLry8kobjer+zIvmXGnd9zyKWORm2zjKJ6Domn5aKSs0P3X1K7t0zd
XMBtJzML1LcjTURMAKN+z1C/uKiCz4Cyt2OryYapo7cgLsCVEwzoDny8PPUt7Edq
/J0+2kcraFKFUIrIcz8QkQmzSK1zVFsyeGdVqKdH0jlmIMVjhPzo9XJXYgGUHaXU
Op23TdfDsioGYykoVWGZXz/p+EUiqotOjUKV0CYeYEh2mM112YIK83W7XArAEl4V
fSuFsPVjuQcsMvAdUjRAqhx6UG8UV9kMH5godFl7aifH51uikFRNC+SFX3fjr24I
LorMOv4rQakySZNe82hn7ituOTlmYMMxDgQWDl1oHm1Q7nsgVBkmoiwHPbBxAGEK
1IImJ2M/zK1b7TFFk9IggmYCN/ln3NARJser7RoAkFCE9SpCxtyAhbmzRBuxO/uR
KKYji7JLVzOpyIJFuZ3FeycQpelsi2lObSyj4zL0P+4zZjiPCWdgzayX8/8nmsNQ
VI9wHzVqaZaUAwKdCXqlpKugiD9UC47sb0LC1Uc458B+fysz/1ut7l4xRB6tkRgH
mciY+Z1cHyAmcEIJavCgNn7DcN7mUhB/1cNWOLqq2E7s5RKJlfgB6JCzvUgPzSqE
7lENbSnqz4izKQffDcwrQk5K/cCjc61Sbt5wDziL7SV7z+K+UxGFPkI+xGjPHodh
vMwB5lJSjZJyO/ra5r09IHLfpGuyMH9cPdgB03oRGKXAoWvohR2Kpk7O+jXjXH8j
kXOzqmij7TIbup4t1UzhnumAt9WormEaX0YO0ZMb34J9+sfClQLhcrZUb5R4fmbG
t6Ci2a3rSp0wkFA+65AjlNhybeNOyFIx3QVN6TnLUlOd7rAO5AK3Q0xY8D1603S5
R8Mjgclr5TNzl+DP3Fy6JBNqOsVE2+z3iFTIC6VNbKEUO3ddHXHNHxugVQAv3qQX
HysCglufURZOaN0Fhlj2DUeB1TM/pfJGgcY7xflEICEvHJsO64yNsXMNu8QO7aMi
yymjp5WkvkgPtkjVsyqcJBdflkLcyfGGSmPJsjN63o/s82eHqSJC3ZpS8jOJng6h
WG5rChM3W138Xj5qcenJUMtN29zjztfXMCcfnzjPqxB6p319yaeS7YtPcOoO2knK
sfMXnu+y0VmxoR+pMhUgZ2bGaKUjXPYy9lU5ttbHWP4rdAf/E5ES3xikT3+2OjfD
mohAi7BonG35xcRQqo34VhpMSIZJLDWXtMvtYP4TDM1kZw7t1DOchzzP+SxfpQS/
MsHU9zX/Nf6GAj+C7KWzBE3oelj7EiE5DJRi16mlOEmmJIxVMbvdiilKHA3CDsDc
XJsr36ARIzS3kAtyTDv2ySW3yaD8Tvp7eu7H1x2kBLoePF+JZuWiqLcUz77Mau5n
vFpx/O5g2fSsutOO4nAy7K3x6hsss7HZ4WhkivtAMw/s5Y7OqPuhyTT6gxpvFUvY
uunpD9n8W7m/3lFXWPI8239yn0EW0ECbN8jb9Ca75itXFiy1+XW8wlfmvGiJgZF6
6HIbx/Q/WxDWp6wZHEsWd7rHkMVU7GSsvjIDAYS+6FS2Ri7yM5VAJoghYqPuNXOx
y7AnwURfgQmjIHrSgtbSRsGQKQ+9CcSpL+rPcM4ik8JsYJJKxmwxVoWN4JiDxbpI
H2JmCiTYiDrLBDNjvMrbHymePrzMpvKYwNjG6tqDnWKoIlfqrZvayXtRYutyxnGy
A6QFFGLP48IPrWxFACLxpAMdgao8+uStc2zGHlDqW9FdnHGeKzzgmmFh1kMaag/f
0ZFx21jQdljl1UhlS5GAIUXiwN0JhuEmY194csWPx0WlZadcrRi51ibmMHuTCP6g
VGIIA7WSgVP6FktGGF9+aHsIaW8nxhQY0HYIMFRMG7kV/Tw8z1RfeqomfBe/TEQp
tx9gS6NXMUdjA+Y6gQj+IJXN1ge7Ee+a2q6LpkC9owBrSfQ/CsdIGgLRWiad31B5
YjjtmrnoPultGTc0SN7xLZD8fguj8BzniSPmcjJDfR7SEvUMEYEbAezhS7v/2CjJ
gaQEqrPGcstJBNWmrlHnnWN47s210AFnXvcAqD72SUFBYZyoBH8ZiBddf/hFRkH1
0TnOBS7gKqMgbgDMQgNezL8emMGWu9XP+00ceGW1Znisw8tl3bxemmSfdR+xWf/7
wmMFdsy3aa8EeFzaFm+QSfMihPI/AbOhdpWDfATxoxn1silBs6zswYwcLe/GExww
f5ZbRstXAZeRVsYRBT1xBIruTvyxLJBg/FA7tfK5XDj/ci0yZJsDKWaBTTJzHJ9b
OW1h7i0upwwEX4Rg+Y1sUpDUgF004IVdj/dNE3iliT2GqTSdWVLyqFhmI4DoBteX
c09QCDgXViJcuKN/SPmOjEhUVvARQPwZVpxUARGiqmvQc5gbas+CXSMuBuugswX4
2ywEbAaMwbRX/NuAHENJ/P6O9odFHBFm1ICazKswxWhOf3nYgQFEFbGO6YmnqY6J
x8chiPkRuES1hX7LBMuuGeKErpgf04mKVBaZ+BXO8nlgyGKPIsH54LoejhwL2PCH
dh9dw2Ga1zVhDIRJC+Pg7fp5ag0H06KkTgfv/UGVsnIar400zyAsDvnbiOAYth11
AQY4Fu87bnjrK/FEakBtbx5fI/nsPEQcOfkkmHxUq472CMTsKc1Q8xC5IJu3b6Y8
uxz7/9PjfVCMoOuS3V9UWSzKgdm9o0GjOhfLuPwADs+mLMBs2jh52+yKpmXJ9lDC
p5BBbsvsWkRpM0C411z4hYGrpsMYw1kON9elRFYRpEDndQNpGF0zIz5m0zsHX99T
+9obFUdH1Tz84dxqOmb0CY5mYyIgHLhb5g6mwKnR0Om/BDd0GKgckORj/LeeiFRk
89QNhBZNW02bdlym9AZUOroDDenEzpHDRh5dfIltm3WY0oCqPrpwHJ1LUluwic6v
1SqW7A5IrwRa0EOcNir0TRzeVv64rnl10B27Pb+pkp97R9NpW2cr+Vr2FOPTsIML
ZHBSGijXsRW5ykq2fxiGdKWbTorbNu7K9ZjDC47uA5YM35W36pmtTrKuxauR6XT8
7v5Ulz2i68O12DAhniSjIoBKc3Z7EATkSJFjqMw8C0agzlDmeNhT+g3QC5Jb0F7Z
DtLLRJxFmAU63RZnJI2+ARCRTADzeIigyi/S+rnftudSHnkFznzmbX46NmrZT0gP
Zn/wtjwKpYpwfQ9aIOaP8QShE+PlS5sDsJ6mr6NYZ8qeCqpRuZd8okJkHGpphYpM
af1sCwA2hCKi75Ocuw1jAiB75zkccddEXhTTlcyplBCNuIEgsu8t+f8iXpTQVEbF
Y0wW2Hm7fzCXdAOaCsQWoHJajg+xJ6Li0eKDCsiIG+FJGtZFDes3JWGA1syGSaJ5
xdhuky4z3jorY6AQ5d+m6m+bhZUvUMktGH+3StHlhpH9PjJ/dxQ4oWiIqKrzGekz
oQr81ZTiLhbYbGeZUuT7HuFvTQMvCxrY3R4W76t5wWcXqtY+AxLjutukx2t0B9xU
NTiYtFGeeyWAyWhFvaJ2aImSrKZLuZXxE9F8jkMFEPDpWL6UL2OnRMPjiAwLugGX
zJXEmNglk5nRDD/qxoIg+WaBuznaTrMRQ7jfTMP0d9Z015IgmVCrY083ogriIbI9
sHLZJygsJCYtRO2sYRoHuxFL1LJ8Q9MrK0whgLt+CB4ExD5BXEsScGLIu0Wh9Hyk
eTmTGZTASWf5Gp/mapvIQM35EtV2dkfKy/VH8oRWEqQlCA9WynbOOI4iK8jeVqNQ
edS0qeYQfnYob7E7MGjX0UJAms3SzLO4F5YjeWWyxfOqlL42fup6DJwoNCrAyCPL
JMaytv1pdUpLyuzAbJh+7F2YnQ/cuUyoZGxu+Z89Eya8J96UmO8AWHPskLvd7Qev
zTdxBvZbi33Bmvu/1QA+8X7Uo4JA4Zqo2VO38lm8vLqF3UEj7J0BcOrACT9YYlm3
jsdwmvyRrLjSndz/efLV2ZoD4spqx5ZSwhhOdrquArXFunxirqTKAUkFSoDxdeKL
almZ8KodO6P0wYu6UitUy3mpAXsMdl41CXI71keZKQW0d3KoR91dE1oW4ckJbFin
VNVWDbfGeffOJqE49hYY0yjqTvEObhqRrCfC9HMVQo9Xt8U0j3A0v/BlDNiZlNXY
JGnT8fiLUOpq+M5i8WKR8Q82qCi0BAoA4bmQz/51cUOcSdvepuBu1c3Rrh8WXXa0
Cx/KF9yxLz3EYgtJBo3Sc9hgfUoH3k2aErxdkMrjJjSGq1d+hOIsR15rz3jbYhjw
6athBoMsrwO/2Th239/YAtpiKhpsq1j1w3EghqMCUCbhNy3IlZoYZHQrTeRhlNKq
TYnlhmzdoHxAhLg/OdIUg3pS6VczGXJPzHUlLgc4e4SDZVY9A6jjYyZkp3yGfYki
GvPO+9iJZDO3qNCkaPm1YGZxugC8Yid9CPw4LztCwPMaK4kqgKmQbVWpb/ly8eYx
muSzSeQNiyNDNtDAnsmJjoS+a+3wKU4fjnU1Ty7SGVZNewB0ddTfG1b7Hq5XlHGY
uSeR51GoEK1O/c3+BO93rLvmhV7Ws+yFghe2ot/j2ByR9memiwALYEim3zmYG2BZ
TIfsGLqAQUFsMF7ZtXwm4x/IwjX4/QvXz2kTuGjAwrcwzjSunRm+IObpioe/nQjn
ipVgO4XUXA7UlLnaavS9MDy6kvaZ6R48OIMxluNZI818vK0ZAnf7kIn5YbQBaHrZ
FNmwufRNsfdY54iomOMG7AJuD8EKtNXZrchWJBpmwh/OfHJzbbg7ELL9Uoff2sLT
6A8dUlluxjfh18Uq4w35GFRnYN8vVKwONz2Hubr221/jo+Nq7IEgzpf7Hzxt/w+Y
DR6ZH8j4aASlbPIloELR1AcvumqzbFNoM9rH/4HoZGvJVjbhcjdvI6QVYsFVtCJs
JAKXFDiP7l3Wzr4QKxSoeXGR4dol+GeLReqFMTwoeppNhTiPSQSkjMHplX53JELN
6kpi45NCL2Vmi9a+MhNIVXqitReoP2udDfZqHPFemBvClaHhfQBA2oQHzz8wRK+L
DxeH17FLmOPU8nk+2dXdyqCo7AxM7wrhuBjaXCVI/FajKP1sHGc6e+gxwIKdriAI
T1lOs9YliFI8jgYOwpvgteQI78tBMKwrKYtZi4Uav1PtbaJrJDfV3TznHZEirErR
rHw5BvBr9jgNl/NeqDhQ8H8xJPRNd0QHcbMuLaz/pyLloZ+EGIhlTp4f+KBgfjM8
iY3vQQT2V4VXTz5k7yJVvWghg+4TiV/KRjd3jIGZZNDy7yGiab9FlvYmzT7PkdiL
pvQzXXbQFeUURMxeZKjefTREmx2g4Ss9osLO4CcJY9dcBDHr4qHyIBtVlVEmaS5f
IYzo8l3uw4j2XeBkpzNnsW1Ew9THRZoY8UzxKx9C2TmjLBmqBr68/G74yQzlAQzD
7G+jyA5acIaw/AqpoaannMk1/kDAMJkXx5R+0JF8mPn8l1GNDwaaIBGL3HMIBIhO
kFpDVfqQXTj6yWWX3qfzRXJBy1fJU/T19VLIUW/oNdOilwbP4zeTcajMgTKz4dOM
tmPiuEwvoJYdoA+FsLgJtvDQ5dhZQaDQUBC70Hi6Qqc8Xv/m7eouTRe/7qX8FKVt
LIf0XsCrQ4qnHqYYpZRX94Y91Uo4UZmCVntVycNMk/r9IPi357BpXMWgtvfZTIot
N5Kw1/w3X+b5QIli5NWTMFGUHBfObtpDN8ALtLq1mVR3f/laNUhFqsRBsmNQAhM2
S5vTBnrjl0fr0HfkrJxUniO3rHA6p8sKoWIiEsNFnho2mo+efHNToVgtni/hTdBD
Iv8B3A6RdCj/l4Q7rq1xQ9RW7jxW8GoLmsxahADp4Ze+KlRu2rpwh5XCp9DJsEf/
+aE2lVPWOGEicu811CmwkTHN37Fr7i5vI4T5DLeQQTPPzuL/Yu2pl0Y92o1bt7ch
FOIbhgsyCTu7b3UrOx98L14D1WXr6k21lg9/YSBTZYA15a3iaU5hIapkPFB3no3Q
G3kS/wYm1PPQBqJaiCQRa0kuY6HunI9bqRezBVqPqBEjqGUp0kbmWZCv8J5A0xa0
6fjtlQV078LTcB4LTfu+KgVzb+lzKLP2YpNH+CeoQhVaeuoEjlz1/8dUkXrHt2sU
QJCO8r3HqoGVYNi75BKCJzGcKdAIduXFPYdl8ID2x/LgyTg2/jEOv8MfF2wQIb6I
UuPkg+t8+CGbYs4MZB2W9WJZr5B2uFrRXBMGDjM2RZNB4I1owMQRJhH3IzsZobdr
F+gqVgVWw/LLepSkxFlR8XMnOtkPE3syoaBujmlAAftD0M80gaK/inF/ocA0Ug5V
Wd9CP+3VEq4WDma+ttkhQxz9Me+riMIXzwJkveaT36AJCiI6rjuGAYW/JSjHpSHr
PbKr97WPGvWUEhuwOwzVCROjfWaWp9tQCEGUAJfB6jC9LWMPpHJ2kUHrHpuDD1Bl
Uojm4dJBvV/AV1gQDFmgjITSikiy7jwbvEu0HXmjyU2HI/Y5ovzkaEdum0t5r7yB
m2wEr97ZP9aw9nY40LopoIA3ZyVOUyHFcX1HMEusG+enIDhaF+qNYbv4ug4sOCtL
k1sKrXpscZq6UwWwNMuAkT4YfmfuWQtmYD+jpyZE6qcjHzutfY/6WnwjfbR0pj9u
3ii+ep7UlxKH4BBIYB/Fo8rLviQGLaDZ+DXdeQFvFXXYGTMo6s6RUAXmWYMp8kqR
o3Yl4vhTm7BU+Msjqfz+dfp6fAafUM1slQp8+K0zQk2J24zFyItaHLuQTygwqzF6
ugDlz2nv0dXNnnkMLDkgrwEePTx/dcp9cYcP+HHL4vtxAxczEQ7nfkfGznuAIMmo
qbxuLdTRbV47JznZ2frCj4XDStxXOmvpECx128Lz+aNmybC9mJhjJoVK/t4cQX0f
aYVLnecvJf2fTDXHrOBRrik7MIaXS9CpdUjca4RXe5x7MnVYxt1c36oQ0BXn7Lbv
NGqg4+nroiL/JSZf4d2m+2Y28O9mvGIXnFeVf30zIjEOZP7BeHIZeDssoAJkCbLK
ill/k5iGEmYXemAhZPXE1Vu7YwXAZS3sI3urBEavKzLdwyJY0LnTXvbLDHWHBySe
IECS3uchbuH7Zq4bLvn3oPsg3dAS0e9r27QX3icbhwvO2jFchjYZv3D3eOGFcOpT
dDaNOTXGuh4zYUtNK3vSCftuspBRFqlYhKNAatiZADYfUGrvjKvays1sUSfd5qCh
eddE47Pf0a8vLAIo6WSwsHafulm/uRQaObL9s/A/eo5QWnYW3KMJLe/9tL5BJxji
85Kvo6h0UFiSMtT085FrhqBIRBft95TYIvXXf/R8lq3clZ6fnGUsYgTZ0XkFendP
n9fdjOYn5qnseazvZ+qO2nDIxWepPk3pd4FvGfDeEoakJZ4kpPbJur6Rm7J7MN7e
I4reL50reb7PffnnRz+mF9dEB6BmxIODFjdMx4R3VjOhwhKbi9xEzdDOQed/zm/R
QcZiQeZLk8b9QWRXWUkKcYiPnEr6NH2KfFPmr6AfJclOAed2NUvYB7JShZWK4hSn
me7fCWQHke3utZhBWU0IOa9vKC9gcn5UcWgY5covBRAyVjYLYmzEh0+IxjtHGmB5
C1fUseODdfcdWA4hiGBObKNZSUxLiQo3H4Ev29nAN/EtyMqOA2Tgx+M4juHQXFoe
Smxajk63Amz6oKxjesuFjjBxzCMPEGYUp/FQyvH4mQfjc1R7sSe18bZNOOe/lMGh
ZP/upi/cQfpSlBneFqF5T3rtXTFNHn/qHk45NGPCnM3lbjXOb2HcklgZWCpAzyGn
UMKJ0fQLWtwuourzoKWueH4KGfFknh1aq2xD6crvFsfvwIqvQ5BY3NYtU3iW89W5
sVn+tODEtm5dtOSGP24ymK3Ebazzbd+yIdgBNlHvV7sS6/oFhOZUfEQeE4B9lIvc
RdzXFym4k40hac3Hsna2GHFoA+pU2yhGmRn7/tjJ0MPiL+3oyFAwQ3emdmWj8Aq8
emsOkXCt1JxIKrAmOyzOKz3fhVJxhgD+epGH1xcK7UrE5fJT6d3mQOp9RFyowDgt
ok39NhmYh3OQCJHWTHE5GUFWMCX3169iXr5zA85UmnyxOSCQKewgYY79H0d0CX05
EmoRuvZSy6/RhaOlFoku0HoH1IIBzsE80kPzIjAljyJusCNk5vloupSj2IVeK0L5
hmEZ8tPU+VXiQ6xYgiC2GnPkImwszLihpX0HWn0ZR50u0fv0YFD+wNK5vz8fVNkB
1o+ExceAqwC4PNziqBXlQsPCgZJeGVzjQ96qSxU7ttWhmnKVl4j10ZvatHskEuM8
JgJluvGj6BlhtDBVwGj66Z4G2Wc4XrGFl/dqgMPumwKm9MgwAVTiOKqirYiO0Tsh
QY2opo00PgLtCKfS/ykEICuieB96wAnPJWMZHADnhGo6IPbZBgXVZrXHQ6082Cd3
vGHRLsK6Un8+SXC4BH3Cl0ZP35SbdjAemVI1dg/VVYJWV5NRUajiItd/a6ETHGnN
Wx6vDaqcb9usW+rjmyntDidCC2caeRHVN1HBKU6YiEalR6OpICcCj50BbcfJtqys
ZtcYyuItGBIeRAqHHltx6G3Gh0+GyB2cSvKE+aVXPnctBIbJQCjYkon71fQFdb8v
J2ND3w0ZoCNQCNI7QEOjf7j3A7nDQwNDbN3bJoQdQuwJJW0EIxIMHhSyh/3UEHAA
ir95y/sIXItssW5DBILVtO65byQVOVds3yordnQwo4aQDRlAL1ePNvzdxf9usIxA
jV2l0lU+afRd+3CfJjyUPTGQPCD0nkaldkEnpPhMRgOeOGV2A03PXVhlByBgOdno
CIjGkMg8Fng4e8li/DOhcZBO4lyfnCoVHD+Re0qHYNp7BRHvxgCSdU2bpyk6xGOv
pW0HgfV2y84Vz9J8mUfzcqByiqzJ2iTWtLWXf+9l95JTxjDOoa30uaO5vkNkAnu2
RycjXwMkeEKHQKFu4mrLSyKa8zmCexrEEHC4qJUlv88cNRFRrOYHuNruRwMIjMVb
M1GRBcMA7NyJjQN2QbCtaqm+s34dSPYlIYIYLmmlTvNW6tyba8LjqB9PharpwCW+
R7AiBK6RMOXJuerZXTgeFLEne6js3a4ULecwyhygtN7Egca0kJ6gbvrFRy6aIPsQ
ySZreccO8gE6WQtvxUfQSZhbz2lVzuAtH/JIXcX3qJP9IEx7Fp+Kxvi6oAP/a5Zj
+5ujzRbji3Tb+ZgdbEiWfx5KDRwleEIVdRU0bw1Aozu3hGsxUI4aALYuwbMeMlKw
7Iwae5jwHnVv00lOUdjne8gxFuiwRUwPrKtuE04nKd28MORlQNvzcaf5pEg8MXOH
/lS1/0128WcHmZlMFVNxiuiOv7r1z671BUSmxtK2ApNWJ74W9audy8Z5WHI0Umns
VH6Ike22fQQvvTRqkl/8SDS63OmWhXdfc/FXyHLT1VXy8D9PjRvrhLR9cXB6wsdr
s2v3GUqoPUZ9RFdyAL1qI4TNpAK4wJ6uIn8UCSAJazRK9x/wP1xrA2yD2hwpEa9S
QvpGK2eXlGQ22YZIo0FiJJfASrlH+H6ln2JBZaVtzm8nAcmC1xXqIzk9WAUl4/91
qotQBrmvrv6jzI+3MXnKbFtdh5wSlTdsWF4n60EKSP/Mn5QeXVCpz+eERDPuAY4f
LpbDPG862VtyCqAIPG9XsT035X4MqSeON7cR4M0cCtCgzK4mCnDacbwedVF6sn8E
TQTcxuSHsHo+TnPkSEx8mA0I0bQ3B7+1UjnNTWbnVa048AedjASxOzdO5JeQ7KSu
08JBO0pISB5axuM0M2u5lwr0TqtVxJgQfbzVf6eETcE3/YuiOGYxlsvVRf+xtjL5
Ju1ArjqGa51aUkSQ3C7RvKexYf4lroIYVTwynE85ku9VyfWA7DB7Ka0jzbGJvWzY
qKHIY9prTnC0fG7M9LUW2u0ceMJ8qhNxH4cKJ3qvKSZzsQw9N7wB3QoHbQqrZWe1
BPv9tKCvMVFAJW+poNI3gCBjeGuJccJjQ3yDV/d9vJKgaM4FXhokZ8qNcUD9UInN
jdg28dn7e83JHqmm1aZ2c7B5JRx6qF8FpRQQsUT8GmSWJTC5CdypF/l6t3HwDZ98
GRKBEdY/0EWd4zMmoLT6nnw41RvRYocv4jv43Ex+Ub0J+Jo2r6ZXchCYLMn41jLw
jgMTKWNQYuHBSsJuveVGkweWy8RIrjFM1JGcRvCOtwZY+4XRq9Co39hNkzi+FndK
mnsO0Tm1FgnctmTX257y3VdMWr/XeUZpgs9WrRTFiQhf1wNzwBkSwpG6XTvRoWaj
tVSszIMH33Jm4R0CmgiwaOxs83hgpiXMKOqLUsWFILcrvF+1d8m+gIH1Fq5NhClk
sYBqWHVnyzhBeawRKEdQWtU6EdfaWbdkd6GF0gFgF4ZRScoE0ZKLzISSHcEQ6WYl
jt4z8uwuqWcxJRUx1dDEFgznBU4reMhcZgi+RBzr6hNarecvKt/ZXtryW4e2andW
F8MF4ICqbvBA7EouKHijkZA7lNpIMYujvf/3TmV+/MQrMxjmtVo33h+0yKYUbuAl
5dksZp1n0odOj5Ooji6Yc/I9KQe711ew9tZR8/lxWYv55LDHyDcBiPocT+IiPOYd
KkoV/Y/ODWgmL/QrAcv6uASj9m/Am8mwHkpDxa4aFQkc/m/sc5GIxBXGE/I+xKQ8
pKrEr4yXmi8q77r1OEpU8j7pLNsYMTt3CL1ypnrt7/SZ3IjAYN2Nd+aIUoAtFzxI
6O+ESGmMJhP3Tl1Zgy9nBYYMEvjjljxsx5XaRsZWfdtQn3BtC2i//q0/kZj+y9w7
C/8Lq3JoDX5SWP8PteEJL47h2rre7LXJjMp2HPd+/d38/tfFHEEgjLGt/Tdt4a0K
sB7Ngu6VdJ378kkrLeT89sGku1o3gIu7rVx/LwkbUZV6Tvs74kf1CEljVJcO9re7
Rf90AZM6cnTGjMNn0zke+zZLMdrT+P44vXjrQ1g+HRnkGX09zEwjFBnLBJq8o+Pn
FQcr4Unx1+53nWKqhAzLO3lCkTvG6Io2FO/o2gQltNbBjkxpWOwDDn+Qq8AdNtta
R6MPT+LPUuE0TXsXrBQXaSlfokyBc29LL0QGapTEpGvanoR7Kbi9nv0kZk7SQDit
E/J1zGAdha4coFMTn6ByHojyIvNAqETaoF9YRvdg28cdTpiUqQi2g02B1RjGj7lC
qoqyjg2JzZGwijcNDjO6mNvhvjbwZ6l5jyr7cWoHSS1OkNmMWz8yamxFN59zOxG4
qrIRZnjJX/ClC3B3CFilxSnoSHl/2zDKuE2ikn38sqcoPX7el9jPjgt68xz4Ydqf
2X7x7czCPe8pn+fhNI+msoXJtfHoufyJAyMSC4oc7hIUwoGeXGNSkbhRQPa6KBPL
qA4EqpNMxz65GM3Myr+lNM0DPn+rf/IK3cF6DVLKTs55bO2pfrncveB8FNvorIwY
APfsL+JbALHpSRhok9o3f1jjyJgCUB6/JvYjqvfWHqK3SDjFzaRADY33Bb6IHGh0
FhV79Ig2fVpz83wqwwC5PPtvQebFXvxvHTopcKRoaNwwhmpCU4DEmTLQQb7n7unL
uEHgMRv6AokMLVzihsaWpfOwlj+EHsrNo8MlwKhieJgvNJRLzv4yBZO/S7Bv6enc
b6fFr1EhrDHlhgxUrWM+o5z1w0lHRXAlj3zSWAhrURk2XWv4pE6h5M9DuIa686Xs
hWN5ZY2FfJ6wUfUSOJy7pMrp0xOaEiL3OeCUkenywGM0xvIXwoVuEO74ELsxz5zR
UOLDe9NwWFVAn/s33XaVhy2a2Vz5fa9OyNUHDFsOiZHFiQzc786zVErrUwbs2KlX
WhPUJHjWSN3HLhTlAupag6wLxawuimuhrTIKxjGBXWWD9XJdz6waPX4ytcq8TlTx
ERp2kT08+ZEoRoYhvDrRV117q4JPAG8anVzGnKM9WGfXCmZmuw4UVccIRhyyELih
aVe7bZuAxpDi63nU+lgNwwr6jy4F7EyKdDI1CLexnn56DxLWJxSuqzKiyNVcSIt4
4D2sdl+Cv3gnMRVQxs0p6jjFAe4MbQwYaqbvQxYZm/lOqUP2VwbYEFDprHowMeNH
WyJthMdIWQy623oGnTdsIHiLpF4XpHk9Q3jaUpSR/fDnZFKRjnCMwXFa0KU4Zrv8
kX7hhGMZrfk5esVJ24FfHz/Rk2V6kJLUQA1Rm7lm/0cvWlDOLmC/tG6ZIPsD/9DT
o+PEZ26THbRW2tHUHTbjp1G9O2ju85dA5hrszIr1Hi4wHkCZzc00iW6oy9IaGW8u
d0z6RFHsJ97dSMiPjTOcGkA+WKrbdl+QQcIAzU0wU6MTdKckV+GGdvGKsA/H8m5s
oSk+Wa3nwqMvPYthJf8taOHLJIK4XpgWYcDsR+okWwI1Q2jEsRRcdcOHvLFZRosa
xNuZQzwKYl7fbNXnQQzVQ1BWFk7AZ/j69au+UdirYm2VkCQmG3WdcLZUddGKjwrJ
CHr1eceo4GFAwLQZePGzPuseYEeAohDw0/KHfz59YgJkCSnwlXNuVRuTic2O5fH4
KwHyBRVZFtlpnEN4V1zsH1SJ2U5cI4kSd27p80cXyxByhzIPbr2RQD1whZb1qCvJ
DOIEbA1K/Q5MwzOS/Afk49SwIzgGtELY1szMd7zeNk6dZ8VgjiNlJ1hHoqVvPC+8
qczvyNA16dY3iPK76aSjZBe5vV2H6ZxbkNbW5owa2p1242NIaUHyt3kxNWah2QMW
mwXrsqyiU9II1mrM1CL1E6SnHmjCbIwPbqfAnmT5UQeugs3Oy1EZY1LuqIEKyyBQ
JYpmXELAYVhbtBaCNqRgJxl1QvGZFzw8LP01dI00fwFg087HniavMOAHVFonIL5F
ywjsq33Q5S0/2nhAWpMQG0Bs2MAM3FEQ2GNWFyVDxwiB5rjOoBEbyoQdPgYylLAX
BVEXhQq5yS94AspcLLJZhOEv+xEjGIMCl4FTXWUHeJKH6R6+sWmja3jKhu0uFLBe
QVjwM6KoBy2/dGpLrjoybWxnkTKiDoqc9TIQJxz7ZN7jKc7xgQeXOunhUc9syLr3
mqMWrGpmV3PX5XfUfc0iFMWdBW9R45GvQWra4bryFDdkkTLTT1G0kzONsPYQI1mC
P3kY9m/E6G6MpFxk8DTuEIfWVnx9DDRjl6rD3str1jEO15mr54qptWa3Zt6L/c+K
aSJmMtb3MTdGsbyfH4atgdShWw+KS9Oy8/G2+4syudi9kwcAZ29lpfFdUgPJLDcG
3Kq2Wrz9E0WN8h1ZTW91O4gOO26tRlrgOEPF7HLa7OaKh4mT/+0RpsxHdwM/5sFq
9oC2I7YuT8TfGdjak5m8xS3hF5lq/gnsWkEF3RncsYtPSiE4NvcUHRmHQTA29iQz
7CTwKBq2Igzk1mxZ80yYz8hK06f9T+WA8KTsi/lWorbiME85Vpz8htW0YNAyV14C
700mvTFwyEOPXUjQqlxyxVR0n2zlsv9W8r2oco7H0SGs89dZqc50Dg0qNUTK94vz
QCyvz36nmh/Ju/kwy6X+HNl15i1zdxmfqa2SKYVjuBNVK3rCKQWYrt8xeShqfSOQ
ZG0POdBEwTW/HSuGLFR5looT4S8M61c4+ckNgYQjpMOzbwY6RqTEUA+h0TidP86T
4ShqLP8xNoc0nTbwz64dyFXbjov8hhlBqh5sd7zpbKT+I26DWyIzMm81/OCR6QnH
f4BsM4djqrsp3koyX50+GGck8MgGZWPjT7CvLVgaSZXICoVzNEgC+BCHcrLGJ56w
M6r+7F6UkBaWkGg9v/TyQqa646OwD3HJbci621HDwXX0/7kIiHa8fg40Dh/JPC5S
xTPdjRZncPs7W04W0KEm9VAGN/U32r07d7T3ME58ItxI70XvdPFY//ncAlAZ2BMX
IPkVpK95gkVK6QeKy4F3rvL+yKFToDoyApqTNtpya502ev+QK1mjLsI3x1ta/F+d
eexsIm2+A5GGCXoTd9I4XSQkvntd6HvXCinM9V3FdTvsLKDABVIY/85QPVJHrCl2
fNIRWueXB80cwpmNSNmHkbV1WfQkQUnmb320xUTukulT1c8BEPSj24HxQoOu6BT1
iEbbGvFc4TBoglS2xTuXVhSrlULHlZWt34/s461qcFqNSa3xeNmv4bp8tl6okaeL
emgIfS/w6xXlrfWgoXJp2oRgPGcPUagcrWqteR8HASkIjqa8A8XafKpbDdUiltoA
ibGqDStWb5XKXTMC/UkAPnt+1UvPNLKno6KL4GZGywC7h/7Y2SLMKLRfutYIl9Hw
PxZMgKiGdw3lNKwiYC8lUwu6YC033ktLrGWuoRhklCpCsJ2BD88C+OEfjM9PPCE0
2qZZK0KL420cGHJgfU94iCTAfP6mzgQ+GjKjlnq1IB1YLNu6GCpmK986bTGki8bG
5iYRXzlDNKQUgc3faavFlhOX+WiRjVkO9gU/uBHtfPM+ibbxFAXzUKY7zNT+/AhQ
TFua+ccccPHDeTfStyTMfikpVzuLZA6XsHbLBJbyQ53zDrPTzdRjkJHLOyfYZ0ez
EcLFP1HFM46Bm6vS+KNtkmYNzT3FOJiSbeMRJBmnwLQsCVjiulRw8389PUHz2BqT
sR81I8NI7Yh3AFIM9dWghbW2UhnjAHBZ+p/giaBojScuWdWpoaThqJjPnyy9aIEQ
nu7CABQ/ll3qoX4VdRtIkIyMt9X6k3TlxXBWfMv2tzayr6wV5mcALlgZ9emFvMbD
rKkCaqrMvX3r8v99j72umgKiYndMX1KyaFpzevaEZj63VZVA0DnvvdnYqhfLXKpu
jIDmHilG4/cgdEJfet6TJIxlsdxyBkmGxH61MDYNfdaeqv0bqwg8tqf4zh7gKmcV
gEPaWpvlkfaCKZIwLDklsk9NFwZgd7w2pdM+7AHWfX0lFidxfSvp6Airtg2QDsnP
cGSI/+wSUm4EDPv/dSFyHZl2bvBTa+Xhy7go/iaAGrB3nLe/1syVtyviNqPPu+JK
T7nucTLs7E8mTLDZHoE9cidwRiYMlNOrMagPNphli5CUu6hX45NPVDNSJ9HbCKOJ
oKRgdwK7SAUNSY6b8gn1+ZAwencQIIdyl82IzDYwxgTvddSt6BykjRXEo+1/lhJB
jBmrm1xzqdTI+o4ujHfDAgjmwFof+cQIx8cKmAyFSAhRJcQC4ulVj3DptW72BHxx
KHY54n14HG7Ei1wXdrbkB7EqHvNH9ulHl+vB69Un29ObVqROLnwHodQ9+x+OoeEq
PCSCdB0gQEuJpP9x1r1DZTyzD7TiqTbvWRZ/FydDqGQ+Gd94W5GnW6e6TR7jNRIp
RBqPDDGqIlqwXCTRySzZDroAVWBrnYO+Vg7nvTl/1IGzexMChWkGzXAN5Qe+v1Tz
j9odD9dcCjzbXUZ7JK2O+RiCPARYzODPmTzgi9heLnsyMuzOI0Xis/r1vrDf/YEL
xEH61xar6AbB5d7TXmbC2UycXHj1x135eAneNUL/yvBZyI/QcmBt6pAOrv4paeTy
jeTL3gqg5nRuJTWIgL+RvTsOKEw/VdUMZymn3+7dbXM6W+b1gGwMc5jjOIdnZPLK
KnTekeIMfkLXtprWbw6eBGZr53mipsh16eJVlr1bCtyrpK0kSYrD6Ly2WD46Iiss
rra0GoQ5na/yHXSvMQZXQJMdDPTpy12q6v8sa1z0BGCzXpxQk64vR18SH7RNKixF
uhHi1aLqp+wsMHeULhpmp05KXP78JszMFpBK0PI9PzFsuUGYPdHJPKUGuMGdlcny
UBBdlfOEoMRioRZL2K3d48v4fw4xXQp4SHbUN6ygCBbHkdmEfhVtXXsui72kRVk3
wcTGHSav3lUXMDUvQmvjXDeoPOJtoIYoZvuTieT+hTETseh6OtOWgJ/mXW2jk2tY
ujKY8noWeYqf0K3Pra+Ub99hx9omb2K78U9pSxKMBZK6BODKYZVbM9/HcaU4YeOp
JqYNHW3rxv4SsqkcYldDajWbCSzKUUvjsf9XptJago0UV83J9wC37CjoXCVOn9SI
ABJIleqUbjUQzgylcUO6K5nt+TW/5XmLOKK13dXs8KvN04VzovIUSl5uXM0AB/UO
CBp9COex4u7VcyWX3vazDktQt1Svt/ORh6jACT4NdQZ/2svSulEISsUlGxh4zVN/
ANMxefRyBH18GMn5UWqdnv5/AdU81ZLcjpTGLZ6S/3y/KMNMtSMVUbif/aFuInm2
WctonDLNOM3wvDlgKu2vPkCH0ncxQVzcQcRtHvqnn+BZZi5S3EFSr8R/JD8JhSHG
9G4fv1Ldl68aqzF8twJuGwgbm3SwA+jnvCqmMFh6b95Rmrg1DQfJJUailJJflP4A
UDsbRI0nN3zhAAHSn01ca+jD4Mnog7G2pcCHExnqRg7n7AkSUD1P8lhYG4c5cnFg
x7xmlcKSJn6qXAxn3Qy8CvxUk6UOhqW57XYtvOtM411zDdLMQj7J2yOZQsXzTMx8
tkx6srYNLh5kvYFsHZfFRl+sOfp6HAF91CImYcRZZ1FddvVniu6AVur5c4I4v+ci
o3i2stwMeTk64zgz5LOC0XAU1kZyoaokNAIHF5nzCI4a8FP6/vY/jA3nUCq8WXXQ
JEqQF5eldLuNUXhNP2bJicuaodcrWgc8oz4udUrQSKE+UiUFqUmr8UpSBupFHKH/
VdLwr1Bt4HbdUstTzVny/EBFjBIhoc/d8NIPOnJppJFbhpnCK/v7aGIZPLwiaJyi
vwCheND/AvQSSeD3cn5JSdmrlMS631W3HK5NdIEZVdXzp4WZe35zSG85j63+hULr
bt4t3wlwQO8rTO/7LhMzIJpX2i6MsBaHN1xjeOmWc+jAgxchEksZlJDhS605cW2W
sBXzJPp8pZf8/DNStK1f/4ZuXV6+ovlklFWy8WYX4wZiDjbXsdCa+12lPSTzGi2N
epncy605IFsowm0ZB0/RYF6rMATCvKMRxsOUZlpdUr07BEJfpNfIFxOZBXNcNBm+
fd1wgVkV5taLFzDfr5uF6S0KflVZDNnR7p5uop+ioVSD1QOkzvc6xqitrRnqdo7M
fOExqNXIHb/rGZvHNItA3l2Uu3rlmPjk0DdMyWsjGoHWzpG+9HnTTojmbMLgdeTz
6p/Dc1/7YVf4k8jrYa4SAQz0ghgY78pM6nEuT9TaGeaxoLP/fSq6a4OPendByhIM
IVR2X71kEhu2HJgQjjtZ4RjY9PrbwfJ77rkwWC46Z/7NsfEMknpfZQo5vYZ3Tarn
TfufFKSGDkUPvLuSK/OkMiT7g6QXWtF+Bml9GMheeRne4kgectYpJCg/q53WvHiK
5QNM+s6TuOxIPayLMHetAz/vY4mhzzq+NzDfvU/4wOWcUFjnl1B3Z09zHngzLlxO
LiM6FKzbP3VShJJtYK+UBNg8JGfaioBRktPgE5rJxtvEUDKjO12fGCUAsfQlG3vV
ZXPNoRmVi5B2Z5eNWjQSfvP1ChQ1k3qlfgKzCzRwYrCux52SYlsSN7Xq+F9gfw1p
EV27nK0A1r3gNYOq40e6XNxsSE88WnIJRgGGX0XR1yJYizik2Cx3t4XYokeyp1lf
3S9tmvaL6EaWJ4ceBiSDr+kjzklCc40htm4m1e74ks8hKPkq7RSoKplB/xyvYqoL
rKlsmSLIKzEcRvsRuJcnQFF47TZzF3PfMGJZzGDSsYCihcNj48QpOLiRXh0gBC16
KcfsHR0sTTGnzsfkn7b0oipusd93JydLPt5ZpZsxJUN5qm4MDTGPbCrC03HsEtSs
fMsflKZV0wBQ5RzhVKciviFj8U2bc4FbzjSsDxw5c5HSXejySewm5Dzd5yHzEQYK
5lmXkKdaoU359j9xxrWKpls9JoKUycSdzDKf2XrPrs91I6/kP51xY3y4u3e1gmP5
i9hPs81RaJ6wy8M2HyYhT/Rd6BmbTHM6AyWB9CTETpZFvzy65E8ldLwQa5jY1eSV
SRDQx42mWe4llrGXmrshk7AjmkgAPthJSX24xjHPSdSshUm8OZgFnWL1hyqMnpn5
ldS3wAik8To+AGwo3xAkz147UwAjZApos8/oY3QsPsaKmWp9ZPO3VaS7luP42VUL
Grbvn+W07sToAutRxZG8s7HaQ4u9/cm/5L8ViJ7gbpiIRZSCI5jjgLqiZMcbYHWD
Efki0bln67S3U01IFscCPQu7ro8fDTCZbYvnj5iMz4pZzBc/wM7UfReBoQPHqWBI
70TGQKMCMiak2yxbhCFLGFW08P9l/Q4l3iAjPjrgUNMGfjwFWdl5cjlAi949aTSn
awthiXsFe28Q6edauno0buTt3MThAV7xqD1QSXLOGqLi2iQNqTsPhCZHtREeecKq
eHVuqfTZ581yI0AUNL6c94Y45intXi+ZzFmVYwxcf6+T3sO0Q20R1PneYET1eAr1
g+PDAiaybNFZnC4v8qfASDCcPvyWlpBrF/yp/UQZMU5fMneKXVaPKlcfgtU2R7he
lgzzEfq0ySpbYgdvVZl6ZbcIpYWuFlN5M1YlrwtxjqwktBCO1WiGmW6ytmngAJk7
8MqmhE9GCYxljohlD6ShbWCviaOWAr0OHO9SkMk6oXs7y/UgdgsWsM2BKBgdgpcn
9kYZzMrBsPHkRyyWNS9hfp8vMDl1N1vtRQRvETp5pTHDNC+wv0CPBmwFuCurS8HB
5hHet9KptI7A12aOKuSYN0UfHnpLVFrJJOMX+Q9qVApOMg8m7Cm76oRKwQvsihHi
mrYkaHXkhfRXLT+CGjwn7+cr7tUyYQ7Mb5jHtF10X42UxTRZ7IgDieZx56oW3emZ
YD2POo+oUplbL+98ZTsSaIkPOvQYxBb96VoGZtHRz3j2KVNz3Rm+svbtw5McCBWA
MCtqhJl7Ront8m+4UjKRczleiNwOmUx0SZqmoHrgZjh9tfZ45AflJHY0sg/IBdH4
SohAh7F8UdSS5X+k2XwwyxExl44P4cKCymz7Odtm+xTdt982RBN95oy+GdJJ3kZC
TT033tPp46KSR/vrUr8ioyV7QSgrIUcvNQz1T4C7aGkN9RAy8VFXE44+X/aiKOmB
4mjj3lS6glCuovGxN7WvJQIP6KAA0AXrtbdHTPnE5Y8vj0LHtFluPAHYMc72Kyks
AESHFY4Jhp5IRNWylrr6uFYk0sb/gGeBOeVEeykT2lPcMZj7MRti9E31hZItt7Vq
9VNPwT1luQmyzbrrdphsp0KenuQjdT3tB2hSphXBtZf2YZGbwzXM9kyoFLpOiXTV
Xc3ATFP/7NcF5WJxG+51KZh7Skz37juUvrZDE0MeQDBwM31N6QLv/0c++1QF6QAn
pkmBQj//EioagWjgm1X3SuNBPS5zCW5RODKHNf+r+SBVQ9FbviDClp58dx+NVy4d
EiXYjE4KIPns3GNRxhGscjFioPNAgxvm4/JZousyqycW+zBvYqW6RLB6hafTMIBs
UD25Yor6dqqOdPV4ngQcl7Kpwnuj2U41J/v5so4W3JiYLId+5vxgAp/hz+XRB3AD
stmBaHyYxgUTkfmT1l1b/FvG2Tj8VBTSJ9xIz+ad52PDRGhgmUS0Jo0qE0/cV9qI
mUwwTxrOou6YJfwE2H2qvacW11Ul0BxRZksQDxuLXLCkyXYEq9R088rtz3ksu5ab
HnzR1EYei5Ne/XTCZsQ2AjJ2zLHGu4R86N3ajHETgbvjG+jpuLwW9gks474wsGkJ
sr0AasBRLVa806goUSCpYVhhjSGDIjFL+8zYxWYbpKnqn14awtc0i85hCD1ddfnj
9o9c2Zx0PZ/ReDZXaG5LyiOIHH2W60+2TMPNxxklfHDDsSloIgiCdYVAYCVV1fNA
eZxtVC/ytm9WcHz6S1DZUF6PzKogU+bBpO1AxqNZ9E8b/wpznWNuf6XZwQO/Y8Qx
T5muq0UiexjA+Vmzy2VbGQJJYbp3r4KTPFpbDSeqL1N4tgAS6tWvPkHTb9IQPTUW
xP3tWTy81ersTPC4md8K7xzViUnt5KonTpTYnonmvPbETAejFka5qZ/3mK1uk9/P
vvVosvpPMVDqJeyN+g5SMzArx6iXXp6MIwjFpyzgrQlYmOZoyBmWZldCXi2P5s2B
YM3Z4Mgw5zAxw2h5YfB1U5577/ATfD/ySG0hm+Xi7DKoru46KhqNpa1RxmgkMlwq
8vhIlecqHypsE/2zPuIUWz7xvwyzoNP/mcma2y7aSqHrzZ8QpPUrZADZ6IueP0un
j1QOsUyT/L6wU2JxOeorx+LWEiJSkVXFvuvMLEVSvdMbWum1MzE5l18oYDY9t00U
0zH6XY15++J5hkoD6BE0uy2tXpr5e6+gfl8KEzVNcmICJkvFylF4xFXvySWdq3BJ
ZBhNEVSZ21U0Ey6pmnxn2K0Bvtau9xMRteVYsVDCUeWrVvYWKeerx3KbTmFSpgUz
YDfxH05uWvFu2+Ckfpl1a3L5sZI18xSC8SsyRfuV0KJvfQJL6GOPGJ1YO3OqTFom
dhT3rOK0g3et3Nb7U6im0DlzLBP6W6/hHe2vUMwBdwDqHFo5DtmiKRXDQ1CLYoEO
EwMnci+eUymxm8FUUe+FutLLiY//BRH+Q8CZ+/pjNYhScVTCWQ6w0Uuz6yEGFox4
3zuwKeLRoILVT1ku8PwH9UzpsTZmquZ/xLBDLjLqtj6u4PeNjhnk1ALay0ycf0nM
I77di+1/F97BR205trViNgieezG9bbKAEZbhd0sralC7ghwggPR3GCKt3IYTBUni
LdBfdWd/+Z1eOtnjXUwk6nHNi+ZVbH+c/i6wAG3sWEqd+VI9ysgf+vZf0/yrWhqU
wK1lleyQjDEbAI6wDpbO6mmI8/v2TaEi4AEEJGftt1u9LccD8A6COqO9fgm1EfRr
av6EJVDFHSgzzPcLLiKlU9FPInoUkpWnQUq1U29L0ffC3/4HJp3E95TmkWzuk6hQ
9ElKb3jnuUUYhGa/NocnHA5jUWd28cr9n0C1AqzgygQZat5mOjMdI54wyXWO1D3h
i/6I99CZRPpTq3e2g5L7jB/YXlg1+kz9//AyU5CnrxAZhyK1Eb1oMFskYi4OXz+Z
yHlg2dADuHnvJzex4wUuZjWOMcmbIPVqXcVvYyBTBLSLUZqhUkzyZ0XUh90G4W9d
GpCxrOl7x0n9PfFAOk8DSXjyG8lbcZFgp9CGwGc3raYJ4XD8JdAvlU2UlfREN6SQ
mIl7tzw6dGvCSMv+jYjXmLilqVKqBlp3yi7WnC7k9mtzTqR3tIoH55oYENqt/NxR
DRaM2e3wla9Y6DhrLEdh9TibhgJNs4IOz6L564OLW7IvNyxI0H2wxWluprcFdjVT
CFOt/XHDNuikIGJhII1PIqkkavPRvMBUkkcmdPW3ftCxY4zgL8MupxjoScmyI3AC
8wfRQBnu+A1IvpgNCmJLupUVm4QgA80sSdS9XgwEY52Ecgh2nGLdrNm7md2DivwV
Ya+BK1pKa1H9sO/MxbA26PuV9N90tDWsLhkRmc2yFkHA9on0EQQmNbbPSmHwJnGN
Ecj4AkulGL59RTGj9oUOkG9YBxjYY3Hg8d8qW9YviJ7OLqMkjhdwj/5odoeE1lIw
WVcHLOcPA+DI3q9j/kOTTvVXVgjI2bB9mbvzwQ+72wf9/XFzuSFySpbm5mJJT/WC
r5rJGaE9cSvlX/3KxSoIKWMesDNcDWoqWGEUENdK1M771MbYVzgHY8fWxV9pkxPl
yCim1eL6hjcoEDCM4YsVddL//99jD3m4CO0Eb5Rlh073jAdVAbpPGWqZmK6+2VUX
CR1bo8M+nTnZItruCwxcA5npYMkGIELlwcC3Ji4t8N1lq1DAMjXFhrSXC0km9zix
QqGLLp5HgzlQDoiY9dMoSaZbK8IetmukJITyp+i3NUlrvv1pvgwGspEcuXPv6lGO
iMnBF5rl0c0ILiA9spblDKUhJUNmJYsfRWBVhCisUXwQ+dIW+ypRYeB9HNAl0X3E
w2kIgzqaYjCjc8hniwh3+FFQsRm3FpkLaWbJs8hyVN4za9VzUJKbvKb7tovRv53k
iSAs5S78YiylXvUiCmOGBFk5s+fsA+W5bC/AtgTYlcrlxmkAZcgJenCVVfCJ/ND7
40rJsnG3s198DAvm76UWX4Cz85fqsHXVsJ1OK/Ahczle5+sVLcy4GQxKuqIKAZng
aiWpnWNvNPOqSW8ibfc5+PmrvnCDFLY1eU+pIzijG0rXrF+J8HEo/9EQddEbZm6x
9crPMatyWuI+n0C95jMq8xfxju/9oOoGWHrmh+Y43WZ/QJDgWV4GIyD4jsyulX0y
LGQjNAB56tIVKOfLppEKJcIVc+fpGpltwo8bMzE498+Prf8dDo0QZaHZ/n4UNCeH
dw/eBIbtgdFJ56lcb7dyQkO2kvh1YvMnYwa9qPTzm4jBHJ1JG0HNUfixTBLOoGx2
jKNYXUCHOVvKtRkEPQTW+xyYElkXwu7GF+JnOMON4jQ1pH3vN3fTDZjlNDLElrke
/NHwU3MTvdwUWlAqtBFEEGril8wC3N5LbrTdefEf8PF4RqzdwF/srvahWl4aRdbY
Huu1PY/FJ8IhkH530WnR0TQrtol+7WtECrx7WIGGu99jyAShv7raEQ2moXXRAMN6
vBy0/XX9x47s/5cys4y9Y8+5IK+rTJwZxhIeOwUUkfVbNRYvb8/X/DdhsZQ6SpdB
4VeMD87TjaaAVSBiDhpEq2JBhFguQIbH0ob7TOqcCtKeKC0twLB/wfcgNM8Ilr4A
/NGeFRelDGMVzvukno34qVNXT4twYbTTo0RL4iHfJe7WXQTijqru7/iqMCY6xfKS
CbWDlIY5/8+TbiHQuoZvZnCGCsNb3TICX7phwhAZ4QWr2RbhOGQpiQXVY0gemiKJ
RI5y5y2+6uEyrOga2eX2cby7H8fw66zgM+jG3CPUvTTtb1xsRWxZVALF9N/klpVT
YhOmdAi1y5GgxX+3wdgx2o6G46Q1see0FxodOPYJgzSAH+C0c4P0d+gTmxnhiP3A
O731RdU/5wAG4yviH/AF+NyqI1AItAoMX4RfdcU7WHf9tQOM8ndTbnU1vstcVyRG
BYgy5awP/2pAFkFXigcE53bAgtUUPuq6XZcjNx/hQTkCJzR75dZwy/YBNuwyXz9O
atcJ1TCL7kJaRVwTd3ojnjCtEdJMOIL5xiG8v+QAf+/hRcC+sWnsIlRGw30UJuNn
JxHLz+wl+siwsicDvqgh/49tfQdldKzlnMeAA1Xz8hBJT4xhJPhFkgJ3K6RlFI/5
a1w8rGwdiI1xTUFPfyqxQ6kdg+8rJVRQA1HXdcJ7VtLtENvJXzA0VuiEV8Qduhz0
h2jwFaypF3hf4bnYIU+B8iBN6NFB48wpIvcEXQjvxdaxGUhFgPa4G/R/0fxhjcRs
PNmAe0OSfvr3QIBKzMGI74rEca8V/JA5DMMrktYZ08Po4IHybeso96theLanOX8W
r8JvbTq18O9YBqczOHd3BUQD+wH/U6XFSNV61a4++RwEm4Rv7sMIoejzJMBtvy6V
FZfCxYwrPnDqCO2SSpc6LgxrKERprF4Ej1BcGcrOsTVwaSOyHpf+mOWdTNQOem2d
raXaHPsa1yB+JOd16VTLXY92zqhanWP9pDktO5iQwjzUea/j+2tHxBoqM1iNEPZL
kGMLvevDhFlcZP6TRTmOygn2BLEvuST7XxqUYPYYB8Jv5DO75eLreoPTl1xQchEC
LZfk7ktl0nWNILl/vkPUtkUaSIlkXxDC26ESF3Q/OhGWreldxsmtEI2bld+XeLfG
JgMZVM+EtQ19TkJ3UKRe+IoQ1oY5xEwVkfX+pFaYzS4EgM52fjJTkUf3XhL4f6yC
OuuWwvW5tuZhvEmUt/BvRI48/K2xPwrvomx6oURf++ozpkoKDmGeys0+SX21PXkS
OacSZy9pCnZHTe0tAKqE4BgRa7EkfBH0j3aI0Fa33zKCobGmmTWarFFBwcFCkynG
WOuUFG7u/d3bLVZN8ptlkmb1BUDW0TBABWtYHbi8fqFlj3c7O7guz1Uvjfgj2HwA
p0UbisVbP9XFPOog1jV9GK9R+Nc85sMk33XdIKMQoVRXJ4Q5NtSIK7TGeTOCVufr
1B09ufSMjshpD+Ybyv3y5fd4cbwLyz2B+BDEAwBB0/EDCHvCLuNQRAkjVPAXUXFM
oGT/rjTPUrT/ofpvTPt7r33TdtDXV+NGtpdRhApO8iJTcOztGarPHe+rMNekcfrd
WRK1IlpJ5e1HRvzB8PVg3dh7JTGQKLEdztpu9gO2xNt4Rega7FB9bf/3ss3ZzjFb
Th7cwtwRzyfmWd03ukB4zGQrIVY6WnmJVx9X/0pMwOkaRq59kDP3fUZdgMHG+fSQ
Grs5t3/eydC+4Naq05nnusWZBnJYT6vPHGLD3c/fujXac2XyKNO2Rydek98Xy8oD
wkgwdsm0NzolCLctF/zYPXHkDPMooeaU/rLMnpo314YjcPerrBo8qn81LeQWZVI7
dYxQfZCbq8JRzDwAeax/5L2uKdBhhz8K+8S/4608kUw7DilZ300jMWu5XXx4RV9q
dHNQSay3H/lkQtS434EGaIYQFaNVXpZQpP6sTIvBI3MCDpP4YJpEN8FBgb1aUZFR
bb8EP/+lGm1U2kyzgkBvXt07hS9pCjax3/qrVsQCsSCJcMyzaxe5fGHQXbSkynE4
w3dmXtrdC/kycXbBoFxhG1HsOdAaklmMALY6WGzD/u4vRR62CyiK4sDgiseXr5av
WLKcUpH0xKK4NBvNDKPCYh0iTnnLUt7b2Old/2cXEM1TCrA5vlVP489/AHRzFgPD
Rr15NptSd9MQjwnEOldrzkRVRXZ/w2gcXh1goclz6IsyNXdg3VXBWLrLsVIjOEGJ
/pHv6LMZiqRy9TCo4fvlcMKf+aVbgoKy3K05OD0r8taGkJPRKp9KlIsoI7Aa1E9U
nNj8+9c8kt14WrHzuD+VwiGYaXh+SiLNHRaqtAvtJCGwwf5jdatLvQlebAHcn+6b
TlJTqAyLxl9ugK/UGv2R7qZONAL7rfdHeeu6RazUUCo1Nci9BrUSlKlLoujzWFBY
+RmUS8nVRgIUvxwVrh/eZaczPsfnA9HspP+wKwqLyoearCvBbXlGCY1WD3Pj5IfS
0LBRlvznMraqe47xCXPt0yX+As1apBG0CRZxfRHzok2iHGNcZ1k5elffzQNwgItD
ZQATNSmDveEMCscp9cuiOkJsGMc9hqAB1FqEUiNeRhis94X61fjwWA7SqWeRpcTB
yVDtx3ZuY8wLPr8LVus0gJJURMM9rEsTC2zs/9Z8P9IHwxvIJX7+f1mBXocMbhZL
0+mM2pqp6eJVra9B9kVzMW1TVagTVr6ExN0rATJYXuXAtHUkdeESaYP/+Y0EA2J0
0rBUDA3iyYzEHHVfzlreD7w1qT+m0ghVFA7Foe/Vx2aum+JTaaDo/wV8mdZpFdIi
dY3E5StcpKiYqmA+Yu3gapsHYkznytmwM+UuJgKy5lNSbdnhj0f8kwXNyKU301ho
27xY9F/uRcogV7FimURqzW5GEMtKr3myJ7/HH1/wQ5sVZH24xBL9wWJiZEEk64KS
pgIEGkPNiQRpvn6mO+LpBlPvebF1P5H0L3JE8iC3Zx5rgE4+jjWofhch18u2JdLw
OPrabCZ9M6jpJRqOp5k4dAdGmZDYEgfCjoBXAM+JL9NKrNeJo60bmk+u6jCDbv1F
gVJvQ90E9FwKCB3BisOb4+mzjasw4u7Z4ED2vqO6nyx/b5suZtDYpcCSJu05qSR7
ArMp6gXAsd6wJIx2Yxf48qXqA9i7CZz9nH1YrftTNSxu9lFbsFkIxYfuEIP9n6pC
XXPo25/m/9r+gToPET5o1szCxhJMTPA6FULo+GBWj9iLynJuF9kssxYzCo8zSEPA
Gi5LfqGittJ8fJIWqM00ZDzCcLK0Vu/n2JzLy+HQ1hhPmA6tVV77jHVXLFXOQ/jD
/HCnJY6KtBPegFYqv5noAqmnSAEKeXlxaU6ahR/MZvrAHGgbd8PLOJA1IeSYWA6P
/2rL6y6shiUln2ZInnLPyIL1RZDTJ7iFPfN6qp2vtXQYNtpFpfKJOVc+CaUryEIk
XSxBuv+bCyRYHQkcsFL9fMJJG78QBXadcjhDGOIfWX89GE/cw7XvYK/TRFMdrZQ4
bnWFzI3R1kE97wDOpINaMiqPyMzdTRUZ31JjeuKSC42in7EzFG1S8tL4XHr1jTbj
VrF7MCk79YXiUk3459wxvbcnxLP3apKREUzT7WG+qUEIs4iHrealwzF4TOnpFm8U
eTJdtrV62p9zL7iDlZ72NbbaYYYCS0M6rPIWiDTJYq21TBggFsUzfzV4moyZ8xHW
wJx0wx/kJcRCjZk6zvsZ4Px0V7WZQZc/UMt0Isa6a23hTQ6Mlt7pgJ2m4CpJ39jD
rPEMEcLAu461g2lI5RxUsi8LFVq1GpwZQ01AXrl0lqGH2LQVi1y7hc7akb73EeWY
t2SeLNjcoS5sLFuCqxEGB1oPk7SqjtAi7jFtXT9aFVgb5RHPwtAnHPVBGYLwyuUx
+sPUENGAspaHv3YLcSAs3j0FvltmQXMAsD0LUlefXzR239uSHzx8A3VEhIgLwqpY
Qm3i1L1rOfVSsBOmWCQnHRk9EEeowPxEqqBYsNamErPqh/1uUaVqyHsdVmcSl5r2
QOhlU95QMEQ5wU+2y3J0AVbz13UzxI9EoAq+WG+Ms0UyAwhnXhJEboscdhGxPA5a
6IAbpJRxu/fYkBIpRH7LpJVyWKh9GTyHSq4awAUiafqoLmGAu5dFTA0TZXRSDL+K
1/JRziwQ9ER4hTtROB9tE3Hsm2RMx4dkGOhjf7rtdiCJemaP4qxfpzXsKBoqjage
QVt+JPmn4gbBS7XkMWHXMxnHj5fQzgFX5CsRIdKCMdpXHxGsBIvoXFdC9AGgdYU4
+9w83C6/CeKlD7Td4dN+6ZeQc2awY6UlxgSYub9LoXyUTBrbsyMIX4bUwk7aXZ7x
WfgHsnkrR624Ws43Q9CJWvXxBPmRR0paMb2jWJ8d6AOITFxWV0mKU8a8FFFwc2x9
PnF4sLnUGt3M4XpcAJRJgOomqSOBfpWhOs6iQANJJUOUJ19YKpT+xO5D44KQRQ5x
loKK86eX2CaDAWR5V4bcU5Y1aMaKSzq9S6cT6utdwV4JzO1r0PBGLO5qFmWFUcaZ
7P2uKgD6ure/vy1lTBnxC4qTVQgXB2gGwyQMaD98PEDWsdCQ542H8Q1jyS0OpH1Y
LNbt3+oXkGo4m9+OCHWuvKkHxGEOZttlX3duJWJh2r0pXDx4u3MK9NT9MpEZ1HPu
DbnT34WHBGj7ePLWjsjzKEv932jXzyqR0ct9Snu2N1MZ6xayq19C1FJ+hqBRCmAi
+Hq8pZArH1gQJ5KS87RdWu46AJKVXUwHTO77JBop9up2d9oiPuUn/bCkqUBeYFt/
12SjP8cA/zHcXoCPWPme3gYo7DOitkeHR8xnNjQFGifbIo9OdHUAuv091TpexwXt
Zr3ax3OHav98/tk5TxkluNAk2dMXSoPOJjmIgOIJ2FI4r0ZmKnds8WARE7ZNEF07
gckETyEyGLcI3Q6fwVLdA0lE3ky86NwtwH3YThaoaC88XPDBcCQkmJXruNWT8V37
ubTXunC3eYHRI5eRKxNcRSQWYBhGSHEqLYnI2LkKrzGAPR+igGA+S/IhOSGo4/Z+
mhwmdcSvbf0cHkNGJlfK+HbQFF296OAJoNSUA8JXAuM7bIuTCiJIkJLnyifelAXL
BgTiUTz+jem/epPrZ6u1/NNYX8UCmwkvTEEmlgiLQYaZDyBmrVHWlKzwZPVRqXTP
riRK3Mt9ihmSyFuuhNedCQkSZahBCHrPduX3ArwztUu2xz+7FfQcAwfN0YzbICMI
JC8A69z7HB6urMpY54XMvdmTVxPMmLTyxrQ01OEtXZDwF5VWn4soY9A8DO345ZXu
hR9hs6iK94Ryp5NqT9Q+Y43oKQrp1HqbQ3pI0BevNd+b7/CmX+gY9I0DFmyrWWeo
hqPT0eAtH+qMk4q/rq3f0+Iq/P72tQsDEPhLwuGNLx04pDsbC01KWC6SORXmpNEq
1Rl/gSXYMfJB0wUpHmLUE+SZkno9IKJtqR7MXqvJubOWbkRKw9hHu7n3xL8BKl7r
QCth7a/E7O0+C4h/+VN2sxIdhXyQISKMdK7qvZiSRFOTkeG1BU37idh1NhsdmL8v
gdJBRNBVx2Qg4mMSiMyyd16VXg40qXO5Teb5hH1jAyp5ehGs7mDAvFQdRcbiJMwo
DC0bQalApaFDAgwUtvcjIm/p/uZaGBnoGFc7zEAMwKksOgEUSPxWTaCLFjU0HNQs
6Ph+RFYu3aJYB48HkQPBBbTwk4rFtI0SaIymvfDug1ReaTeYTzJ3vpb+oxyQtYkU
hnldVjOUkU6Men6hr7R3cxxbtHHjdUrJtlIXqtzjuUa/oT8wVfdmOPoiXmXVPCvs
/L3gFgNZouS/rJPrWNcM9lq44TWm3dpOP+yCTNhIwg5B2TmS9qtLZhHShCG8H2v0
QmwvCA0+Jl4PI64PYZ5T2ma8AFxMxMKUSAoQBFewFnBl0RRC8cIS/qWrLU70Qw2S
SndjYgSFk+ktLO0xQkWxbNlOYChvjc3i9S/74hzhQp/6azbuWy2HIoNuQPbDRbyC
wLB6LiEW7uSzCFXhV/ViYu1VORROArycnRVtHOUJeM/lAjV9lnX5FggK7fH0C8lP
IJapEWA3a3ZFu56xtJvLeYyd1q931US73XvyOY0xZRxGJQm6AmJ6z7JTiiTWHuD/
u+Yig710vzCTorJK6vGk9mZnDBbyYR4gPRVXg6QtAAndSwU3/61dt7Aqs6nYVFVZ
5Wa6vz2m2WR93TvM6ma8dXshVrO2MnDYjI53/Eah7DRjrU7TXJzeArLSRYXUdcBK
VpI8bB7JGR0UVo9YAQbXDhsVwEQEhSw13jO3mt8Nh/0l9cPGPMaCtw34cFfXDmNF
QSNBWDOsF6+vznvd0qS+/fA2mPGExyDsk1tMzOBtQfXi3aTxoZjfZGGWDQGnQef0
tvOBP0R6Pwv7r5izlnOYyiZjfXvF4b1Ti1wsgmC7kJRGyVUs2F5sGZFhDlxx6pmD
z3AVt26GojCUlDXL7FlEd0knOiZMZQ2UWV/oeJJpH85MvYooXwnfI4tOvi/esd9c
tN0Jtc7rFQZRaQfRAUW/14L7y+NM9hwHc+ym3+iDEp1i4w3IuXJcE9+NdE/asoRP
YNqCxS33en/hr69KI4mq+B2x5gquvj84A/sGyyYhfFqQPum4lpcnb5OZUwG8fZsj
woWk/IEAHMhGkY6j2kU/XtSb2HrqnJhJvO08UJ2ksgYNtp4ulvmC+mimogdTUdrQ
ZXQPgcsYZ2YgTdFMB3jSXCfhDy2oD8HeMDjHz+5DEkQBtFmZTRCsWzPwG9A2n3+N
BnOv2JtA4hyR9oskIsXKNsgzPXIixJQn3yLY6aUt2u8CYcF5dO9812Be+jmJZVYN
ybJIYy/qytimX+hOwnhPXsHQ38/rX23JYt+3MWlvI/BnIWl54ZAGId4vesOZuPMw
M6bMR0oyNoK0ddosVJMH+s3LKyRwqCdA3ogvAMBL+CUpKOvhacsXxJFYkKQmQ79Q
eaQsknLgPiFIykZb06W9rcyY9DBG+cfISMWJRvJaT4oK2nmxW4PBODQ2uPyiMg+O
S42PfBBntfhuoQrWUQ0DpPmCYhO6VpPLFSw3GEYJqCgHCBDKE4ZDx3WqI6QedX0F
0VLZV11fyjKAzTKkXiKpCEFY5vAEn479ssXUb/q75HD9TEMhI4YaRro/wpzvkjJL
sqFhMBYk6KBIrD9ytX/VBCeBulF6jScsRUmS8x/vja6lDeCurWSRNDjSRQtoXzO7
aFFmqsmQJYmjxucd85+ltDsy0ev6qOtTA/BXYxRZUsiZb4RP1Ezu1kKPAuI13NJc
rsU3UKJTHt2UTyiIZXaasnB9QpEu2BPyr6sDEsBdXWNeuaMmYU3bqi1spqwNAQ5S
wit92SHZZXURkjNoIIlu22Os5pZy1FJs5Htb9Dntnq2Sm/gIxfr5yrdYsW66OC0c
7wFKa/3esWpHMkiw5CzUhkZb/CY71g51X921NAHlFb8GwcJtB1QDQGJOwRSu/rFc
ZBnRkgcuKiJLrCoE3+p/AUorx+d4aTfG/PonvatJRqHwY5AtL/GkKgJOSn09Bpqz
ogczoe5Kg7X8YHGCRxuKoUk+iJMzK1tiLnRI99VLeI8GwF7I/o4IcUa54dAwC0ke
sg+ODabAJRY14AM+K52e2I51kdxVuB1mKF7laLQ2yK06EUjXCJ5sl6fh4N9xVFLd
MP0+f8sEYhzefQFRRkrMweh9aceiemHn8qNAN3m7l1aOpg1Rdua80XTqq8M1aaEu
lpvoWWmB1XSn6oMkAGKMrXApFnbHttYdBwCW8oD5QiEcSOktYcQkrISvGHst20GB
tyS0P+IV9X/uIhvxz2iqOWJ+20fAK6B7hOVLDwoJkIHqyDLBN0KWK1TbsEPzMGeK
shV7+ddO2HZvM1CmNZbG2KFJOZQtuCq5KVL6d6U0kvbZ168UTf3IgEk8GI4mZn2r
ZrICZRZn0u9PFaLoP21LigsQwvlzJPjvq6MxQfcUmocz63UfkasRY43iYwgig23E
bn1OmjCniqZu1RzAVyGPck70Jm5gQEvJxlF+fDSbs3j4hRnvuNnC8hMgM+oeRnAb
hEL/s74ywcUjvtK0ZiPN0eflg/g03lEvTKjf/pTPmtyD+l7mocJ3PuzEtWGp0ceX
0FPwKAKtiiPpwIs61kOlIKeaKpPliLZx+41R4mOkBtcHFwewQQzxbsJS6OSf39ap
D4Yvzd60p7SQ63Wz6NGOQzL8CxZD8FY8UgzHA0PRdTYXcPD8TvhHYdWUo6IEbGTP
QEpF+BAln9rkeeOAD6mzChVEbtQ5QvWO2YebTiva1bsQTEK0CNmSy0eAiyQo1YFy
BWGAQjKWG46kKaLGiKlbrxinvV4NeE/Z639FyUb2h1g8XOw3XbYPkgV4k7nl+4DK
cp21ttm1oJZaBXMFF4y4xPoCuLzLYGy30StUn1qtcF7mI2GHNdiDzKQeehupoxiY
GOQcWAT2MObbKIiIruViC56mBdXos5DRs6PwE+/plZ4GvnCGFYs9LamfNOkZO/A3
OZPYGpIxdfbG8vMzHXXHeC7ewfm/vRjrMbgAeo7c5pHySWHQ9yULK+PTkKK5KJMz
jNOFdx0zNq1fTwf0zvvyQS4lWmUt9moLs3AjoO73KikhBVv0PG1s6UFvtIdBEgT6
+6AhI4v4gQldkSIla9k58FRiYWEIYFz2xun7MTrTRA7w6UU6YZI/pcOSfmgufKCv
sYxIcom1YwFm2YOikYDXT4JYJIyfWWRCNjvL1KOxxpESdFWYHLa5GCRsA7wxZWJa
khACqp8oHI1aQqP8Wo/XDJCduaEFQNhJ2sWZxYhWOqtGw/i5akxR6KUNzm0zT5C+
QQDgmDZJGadKa+QxzFhlga2q9eiibrGm5uQBKL9+qVWLIKDWgzE9ad0y2Ipk/xAY
/Dz78vQcLlJr6UpObMPwGJCeXOW2O/EQrWx1CY5+A/VW7C7JwgeIa9nviAlpcmvZ
yiVl4B+XHE2NY7PHipgpLaDNNOWttKlDMF9RTpcvdmG2t2oJcwAHV9PlzsyZq6rD
bnDX6mWFjVEEVvOAJSYZbf6ckDE/c/9/ZrmhSfMoBigL0g+l6cJFhHntHQjp6FHp
aWMKUwsuYmECgDMEzAzMcBiHchQiwQUkWngaTDtR3xedP8yDRFbME/utx/Zb0m3N
AGhobCJ+dN/0/Rg3CMshVnbWYJbqiRHGKzMSZvbLTsJx7oZgUjakGpjQf4/B244+
ow6h1ragP6T3ZTrXGz4tX5BDNKJuFfXcetxJp+tN5VRAEb7mbrBdxwYjC4I8uK0y
kaAnEuRDmimhUh78XwmHZmS/Mg3yTrNpoYP7yxjcFMwtASEBQTo7zVMP0OqxTm++
Fy8GNTlrc4eCK4wzXV66QfYSwapz8S5U2IbCNjYTQ0bDlDWhnTCBQISaOslkv0pQ
nNvJOszT+KFvEHHAS9XRoSBZ1D+ieU3w/Q3B99RskIax+K3mFavXgB1Tj/as6X21
7x82poHBNHTVIJUcNUMPWENUyD1BuPudlTxLfYXBys7GLFPXMIpVAwj6o2gVQLdK
ojApi8GcATP1grj2k95oY33ytZRsOKfPUWsgSBgLu5k1ceUfL6DoXkjvKpufeDh6
s/3S3Ode43Ht4w7veAgNvfHFAOgGvPg3H/k+E4hE6bqQrVgkP2VKwwyQFK1DFXmI
31FRsJafjjgkYU/R6tkq5C6r/q7e2RzGFYfyPxF6hEg+xLeAAH4ZR1HFWOwUP4sY
vRD2KH9mqVr++AT2p2JPrSHZ+Whr8p5zYpd1vfrAY/KaCsO/wTspXiwd3qXLlF+E
Psye2RZgawMIUQcjJewDXZS/+4+oC3lGKlqki46G93pSkbFsnSPgc799v1TPzaRg
qRxdziw20SF3kvGbqRuTCKfkuz5+fNYti0YnnJtIuk0vfd89GOnYNBgdAXJ/kZ+V
v+0YFBx5GYFHwj5PfdO4fJ2e3zddWPh5yuTgbSbMkUmY0jd/PG4LpK7rN3NIAorv
l4ULOVGLwwXzT/kEcnN9eTUE4AztzOiGNw1G7Amh1DDJkAWqbjcm5DLoQ8jtnDtL
ynHnIC25YEHxagX4f6EewBOyz2lmS21yUM21TTviGb+X/Y+xC/sSQMyCpSxeepaP
dKDJe0IyAfEcZ22Xd9H/Ec/SA9dRtb1hbai07Mcrf3zwla+Emp0QDTUqfRZ5N8T9
mwsDo2iv+ga3bvs+QaRoyLQ+CTSpJMUesiCzoEmbJfF0kThK1aHuv62T+2wUe+be
QKyfmUIy5BXrGl+wHOHIJenhvbGQDRQM20TYK3qwTQGJIyOL0HaBAga/YFZKzalw
YyrbQBRn8f82040oWkcjvz9+frFvIvt6iWZrQLiJ0cy/SreFe/C3nRRxnnIblxzD
zsZopArpJRzYmkKlS7x9K1Z7NPHTBkswJpNY2jork4e2iEAQ7Iqyl8eCUO6MWswQ
v3TEFyoYWlmtjHGiqICcVTCIdeVLSLC0vMXMYzV5pgh7exf+U0VnjMw4INOQtpzN
MnBmyY41kW5jFNo9OZISj1vqw5DfDGDmLm774TEy7XnXh78Yn9cOHqey2i/Nm6K9
TVgFiZGfbLQPr64cs6sLLRIlnilFGLYH7WnLBkR7UQxZh5HVKmxRD4EaGe7fE1ic
R3mKfuU4Rsdh152y1NIcbg3MF4/fdnV+78oL/IBL3m6hG7i/as+iksurlsPTZsGQ
t4Z3UWT+sBt1duCU3kvmwNl/UvE4XsHRilTF6bzN/42pH0vWkZrR0ZZKqV+lEFr+
9VTF9Wg+pymXLcgE8OVEKuQccNwID/Hy7tiEZBH6Whra77+rEsfYcohcCw3dIuMn
mN7cCzwKT0WDmtk4VSfsPZicKOYGElx0074miIksnqZ8Hbrc5/jEmedZwX+iD0ab
ezzb7CNZsiZKbTOui6Ux0owZx6nNupiTPez6QQU0T0inH+HldeFTlcpWJnmQ7d+s
pgfD8VNMYbn94rZ0hTZ+xb0tmJD7GhJHnvSkGUtSelk9XfIxTtBaPam4+7qps3zM
YWSjXKjjIGObGtcc9fotaFNw8gZXKxyynQFGXNiyYIVj4Q04bQ1P8rlAcoiNeQi4
ZWdlYkwHIcWZdgno4FePDKa7fgZxS9Sv7RwGY1wQLe4Ea2+6dog+8OyJcSxgQ3MQ
Y7phBUWh6VwJkZ7H3i4+2uRd0frFwXcjOhVeawW01W/wYYed2uGGPzEPTUyPbdfy
LnQVTWs3LNHCzt4emME5zrz5SRMezRoRJRtI/1ZVrswfXoyDPsA8nc1dYrw4VFHO
l5SKqfctMA4RFEV/oc5t9Kr+qQa0NeQbNDfyDjRe0IHIZX4bcfY77jyAf7T/oQJx
1IfSC2Sf0Sei9W5hEbJjJ2JZ6SwET/STvJUBRT36DKdJ0JTO0x9XwcygzoyfcZL9
Ksc4cfBT8Pe/n5KFzzT74HeeBaCeFF3kfRCDs77SFL+LWc2hvD0ZWsoG2XWmizbF
jhv/BJdYMr+Wkmi/PSo/QGV2iBSN8gTrsLSieBxVuVWMuRBer3CpTyX4+l0Q6Bys
da8UNFznz0crcgYEyCfWORwE9UviBc+EudvtD+IBBpW0WeRotk2zPlzWBhr/unMA
9Rum1DymO0XRozb0vuyLz/UYIvkQ2S/xWSLrhho6jj7bRaTY4aIL52CWti4UTpv6
gKX1yCSTwS7INcxyjrVgIzXOdXrvct5av1hSDPoCrautxNttdbZSf5ndMbXZoNOR
fCAAc9CEyZDLNDkbpZf63o2hDUu519aK5jmb1hy3q+mxFb2DXIR3+fP+OIkW48C9
gteh3k0ouzFa2Ivb1cnqqLINPnzTUfmiAiXoyympT7SmU7eUACzEtzOk4K10N6d3
DDODEvbzlJGToYmiRXhLcrFXx1B5peCL46VVtiqzHnav/NLZwP6PmjTyo/rQCDnm
VLjCVdVzf4jxt/hjhflSTV/kKx488enRdtOVD4giJAauSBvzQDzYluk8jOUo59yS
fgKk2opmq6eO114OthvTrY5vpqd4qbqfrvVlI0VAeT5GhkfGXnoy3QZZfJMQ4l9o
vo31wLD0nfSlPPaMN7fqTiDFoTIeRmO1aiB/QAT4GQvWzKkiDpYu2HShgaxq2i86
kEs4XbNtOwrq+dYTiAaz3hQCd1QyRHGzkdJ+KUeTsJ/ifuiCYPGiDm0lT/FuE3zH
MIRg0Yc4inUx2DqJRqfsEMTbNAzVKAan6BTJpl1nBGup25HozjxWjzk6wgkakLD/
u5GiQBPZ2ptkQ09kO6HAlBgqPaghSzQ5axlWwe4F1D9esmP9pHkpRPfTFaVcHZq6
WAyTpmtW3O+/HyCfPpEe6A68VXskHGV34NXcFhMJ/9veNkSPNO9ja9nOfbRUFxaF
0oVAlreCDf8bTHQlYG45zP38FIWXp2OJlX832GEebO8+KR4mFujDR3Ig/73WYmEj
Enh0Ayaay0TO7CQioNRcrbzwzKEXIZPITmW86vTz5h0Owma5fGX3hY36sYjCIhvB
4jOhAqqUppSb1e/UBogxVEZzW21ZdW3vICpbkBL5BLeexV6CzNR3i4ZtI4QhpTgk
68n3GiRi6UjHGYCfHc3YzvId+QJ1Q+7i537ERz5fCVD5FFJLsav11noNDLjCU7Wm
7lEMp59xl/0vczp9R+ZKEYGAeznn9UoGp2tj7homo6tBhj4ol5LT1OOqfABvdIZo
jI+uXLHIeKPgigA/VlBN0HrU5cY6abXOXww2onV9amCLAjGKcMx9nJ5AuonrgOBS
fcMbw768B+NdE0LVFoElI4hNnMqt+5gl6FpQgj3EdcFiXsiWJM9d56wDx1SWz0NW
2r88NWr7AOJgcANtat2qWqlwQLBx9v78LjnY31XEBaBgmCZkFVSKFjasQzwEe4qk
r+msKuleOZkqDxI4asmeJ5zeEYMpSo8jWKaek1A/Xz1UW3txgOfZh8lbToCKOs0D
EcJTSTsiCsEeMqTRlH0e21yIgBfsMb2tVdif2mpW7dy00VXLJeN44fWK7RgMQGwq
4xGImB1wJ4S9jaOxtGuy0cFZkI/Cxp9rm9HqNJBi9LViaDc+ac1YG8froqy8et54
tkRNnQlArREx0SBnC5W/5WLgq2YUC9N2iuONDfv9c7FMoao3/FyvL8qfLwn/2qKE
iuMMwdB1GZ3v10BhEKwtY69/q21cj5gLFMvnWnjOftN1wekQei9f8hDs2qLOs0ZW
bJNlvxOxftPRRSgE0x47JK/Bqq/OteOn6VWynuMZx82rFpCLoTiWROLd5rmQ2d29
KCJW47GC/dsXwoEPxKvdAaF5MZyZOegkyHdzYPbCnfFHh81aYRnBYOk6xINk/PBf
5+vUGhkA753Mf2ZDXjQW6Oi0lIf5cWUVJPJd1hhdZ9xXjmFZlI1Y5AaIij6F3taC
syiiz/mizIyW5f5HZINVPBwFi4Er057LGc5K2obgLpmzg5XngwabszV6COIaE/4J
Iv735g4J8ezcRzvxAfEtbiSSF1wSdv4iuWuqdAmhs0xxjzixqisGCjMP4UBoIy47
aP88rWd+e1ksXnwznqaZb1QhCGyE9ViYrqeeAeeqNE58vw5wAYerJ+JT+S92zHOO
CvGMIJxR+FrEUMzTAPqo7HIi7l9uEK1UzckiFWMJih++pdGRmAmggbgqcftgh/YD
h1pLWPkPhZLtqmHX1kDgsURpmxERwxZgP17KNe4SPoa45O/XVEWioODX5ThuzJEf
ixDU+MXzWK9wRBMQA/wVshzuPXloswPC71xOXXKy1yrsSnwQt46tNlKDc+ldGRoz
eQhgl+6yVwwD7gBMQ1N5I8bMRxYi1nL8ZeaIyG6D7844MNKOOGm6IePB2v0Fju5h
F7EwQiJvjQ44uWrZ+3DyBEq9B2RIUad3LVc92wh9OYLKdZ4Ynd8Pfer/y//ZN86f
QS4pLpk5u94yJtvA5vBf5ukYgjbkDF66IsPes3tVMAwP/1n4slxyIgxTegYh8jZ0
eXJU/PHzZDbnHLtUrYsDChHeUcwdUNvTsifMpXFLYe8zh9sr6F6ZnFopspO2H/Nj
OlZ612y+b+X1f9k43am/MdF3AP4ARbhxr1pKEjoFD2rwcXpUHSUGjpnT2hs9nID2
XNyuHvOTFZyJZvFvDaXqpggn5h3crBAeIdx5TfwxAxSvNUP9t2Aub2RfrFcrWWum
L4Rmmho67Tm8Ki/iC1dOWRFEKezntqIZ+CjGOQFW2XWrFVo9sh8eX1y8wz6TpqKj
AHekShO/bw8JrZxA8TfUe4VPfKuk+pNv29OI8eTehUJ/8ZZcpIVOhq3W8dTNmn8Q
QrQNJ7N1vrf/lKgD3ftAuFdtgxUY2KZ6+xDf/eZusRbt+b4ZmObL1e8w0s3uodIp
/5meBwsflu/dnyOuNAuraOQPQDrfJ9mVFwf6TOa5jynFDG1wRZPeOpMqGfz6WqUn
7wu+5cUdpPxaPy5Ba0sWbRizEBwcMFJ6vQDMH5smk//v783mvquEsvwWkF9vtkjs
DoKjVttzmhYHDbMf1FytMAedXDLWPvJv0Q90bnJ0fIM1o3rS10Id0MJBXUrWqt0z
eg6L+2VbDUjl8HNFX2U2K8cBdkOipNUlfP1fWnc5H2dAr8jBEhRxcM8MzfkYxvoz
tHb+JqEgRXkBQsPRWgFyQfz6SqVKlpAVpm0fIGFFV5QTBK+zIGMhnafQSD1mcUUn
e8g4YpEPYV9UIXgU04vEibhrdrR6ZGokgd3u2+5y+yghM8AlTs4/s1xi7042PjeE
n+m4M+m2r7LmkSkLl1PX6acpdNI6jJ3eyo/jEJFy3UVmmuVFlTW6kHH/zlNX0T7I
D5i94KwIDq/86VdFPsDLTl73fUJomqioWLQXvfAOkN0x/1FN9P9kSeFvRoRtxe9H
PsAnl7RYOpH5g4lkqyzwekvOz4y/v8sss5T8JtM4dGyVh4LSQYgYUNhMN4V6PZ8I
u71zMK5NEuQlFI1pTa1oAanh4HsgtWnXP560Z5znBzYbtn4GUpmzojfTN7W0x2B6
J9QrlyU+xlNk9scjF0uOoap/y9qkvC+Xywc8K8wNWStvjFD5rrQ3E13hpu+y0yFf
oYK83uk5eFPBtrJY2ObFw2s93RZ77IJOdTMn042WIIvbZBiepgTJCRkpnPT6QSIf
pPlG8RhhoW5BF6cH4IDv/lAk9miXooJvwNhnzpTYyomLuRNZAbZL0kEhHW93ixqL
oZSKeMfZqptIeqPvS4VfSASHfL4Wrp8BifQ2G9oprKFD8ITMull2JLhvBgIxMJuS
BlLslxy7DYYFVd1uvf1DZe01fh6YbZSxXaIRAO51d8xqIwHe3xeyMksJ+ShKKJ/K
Bb1AkLQ/oVupRNsQFBaqGBZ0P5YtvSrbvYWKG7BDfPUoFLwU+W6wgMNnbwPqd83n
U8O0VqdZduMlHSyWzB8Ow8MM+0GWdRGYVpjMYjTmaHFXJL0uNW4BYUICT+jv51oi
6Ce34dHZaokZj5ET6Gqf85KWRu/cLmMRQVhPgY3w0shvMIMA/EviaWlG9mgKHVsE
x3DbVF8pVRVBijqA+MidToblX8hSmWaVQvrYf3ezBglXWRdFj0dMxepoiAO3HWZZ
4i5FGYbYYoL9yEzZ+LDmzkBTsqCEw3g+QwLAs//R+Mq+Yg378cjNgT6RtydaABdO
xWuNOLOh5r26zLzEh6WnRlMCVFfbMA7V0H4QpQBgZzGIcS7u/j0cLi7AzNWFDx9F
4Bt7eColDrEfWpv940J+d4Nmp1gWolyBPKrs5xOl4cVhFJ4VwHs/842wIS/IHLn1
QgAhwPBq87PyjDoZ5y0QhSbYkI/QVxxej4HPy7ovBoji7J7qr7bYmMTDDYzUsy0R
uyyy1kS0UDpjhpk+8dVYmyXsHoJlibTz2XsEA4a9pUS+VWZUJWHBe1t8TNj72dn0
nDDegm1ddaPP2a3bneZAUvWjRE+DQfcuHv6Yp51jdKwhEuSGOBkq/2HmjKXzaG+j
scDfq6O+sdd/i6Xi4TdVD0PWTqbZjnmAt7CAriRUafaWOfBsiJK2v6HAHBQ8uyiS
ZFYjhpEv+m46q3aOwrfwl7VORaKYvucQS4is2y9gOmWBd7WKlG5NKYv7l3tyVgjT
Kkql04rSwVREbJ58EP7BFc625N1DE2XAO74kN3efjjdCnamX/fW3nSF7zepQFzcP
5qGojnultHnTHBjnqhF6xxpl8fQcoTgjiekaCYE4gvJ+aPfX8ZjUVaA57V4DSPbC
TiwEq+LzhB8Y+6lfgwOMD9OGSBANWzYTgHI9AEr48RXpk0Lov0/tDkjowtjd6jaP
hhV7e+vInDF/RImvKXb6bAQ2wAgoD7zAwBx36ygP7w725UWPF1hGSO5I5VeKD30U
0ECFqNbTbEBEwD3G+eiN/QrfcNQj5NL07CaIB/ocUvdtONc8TZAVy832X6XZlVVl
MUGHNqt+SNU+jAn7G7bYWzdPLgZRjQzeYgOFJQ48TiJEhQ61KPkHTnfWS2taihIz
2zl9YlZNZX9qejJ04Mbi5BNoIq9vDXN8XzUqDTLsCL2yXG7i4ChZtzZ1LU5sl33m
QA259yXr0sWhmXteffxP7S2XzIM+WSEYYiwv+MYQfDAzmHIalin1Mj/97ihWHYdr
SoZiYkIaFsl8JNplaJagqv7nRoLGUyzxoO/dMOPpUpTAup+xMGmXtSQHJRy6GkVX
FEI9UKx4PKVRP0VQhsbRF9+seUsOhS9MQkkqIZsm/J9c5atio9GYJqVIT8nxXmux
DcUPzVvKZuK97nR8Vl0U4aIEwOtqdYaMWsA4pB8WM8GePtCEM/zYe091R6ZLl7/0
yUfOu966vO7wS4Nk+32sZutAQkDv4Zta0vRQ0HNKZx0qZo8ZgjoFxEBDe5zQhlIm
2pi/95/Bpl/LxBw+Y3zEqtKXDnMf4D2sKUnmiDI415+D+jhbrRfF3Ehk9HAQGFXU
qStVfpbstYf3N0lFAtuZO/7+v0b/HY7hhPSS+VbP0rn3RRl3o8C0ni2s8i6A7UlV
OtgL/gP0NK8FaUoULbxMem0G5yC0W5elHjKWmZQb6hOKFJBtIlYHiasnr9E4Rsi2
3H8UGgmF0fenZZki8+8thSBbuH2XkqPt/ZBVizzyQtn9Db5ZOwk16OsvkJPrMCxU
WlKT8IgaU4tJaCYGtjN15PA4R+QrriVSw8R1VHZZQ8KWfmYfvLQBwlo8dvqNttwM
8iYY2FbcN/aTrLzY52fBiIUvM1knzTTiSEeTsu/hJe0F1cx91I3JHTRvVuOxZUc+
c5OR6WWSl5bORlo17lZd4WSq5CpJF3N+Yobi+CjxPDKz3ZonN/CJj2PaOBqcJwAQ
LWOOyQ4uaGhWugNwYM3buK6ZpelbGFrdwnw3QeX9lPkFHkpalJibkniSA/RXBlbs
euKZtv3afZF6u6AVIk1CqNhOkoGzyCGbdJs0MLqKoRNeF5+uVFEFvo1TXIVO41cT
ELARAK5CSs8d5gl2Umr4aRIfEs+SH/oedUrTeJEcNYy/S7+7mtgXhSwULrJjv2fT
vLeqMHpHomUUhWAOhq3ah16YJiUaXDx04FKDyMSU5UQYZT21qJKn9gZlrNpLjYoU
LCyUyJ5rkXoG1ASiwjlXNOBwbLVbNpeuO9F/Ip7as6n4eCk+vJvJsYKibMjJbdi2
brY2q6BpcbSIDjNxytdG/e1C898U4lKQZGM9RlLBKu0VkAix/QUpH5bC5DVLntkR
8ZbmYDYNhAdQIUs4VzIdugUweCbar5RMEZRCeEO1Ef30Tl6JCHSA/Y3bTIumjaPm
DRPJSOW3zw+I2Ab6ClvPS+a9fZv1OqUXxElayZSg9ZmXaV349ccfodj0zTmEzNCw
0Ecvfw/wvchRHcYZVy6HDZdgWwYqO5xrXg5L6NNBciMitmrwvo+60+aA3yMhYk96
+FX6/XvAK6qCH4Gkkp5Ui8cCKsu3rPEfLWp3UR2oOBm2ALzUFJ1kgruhm2+ZShg1
BoSHK7iS70/zjOvcsmfrz2nB+ooo0/JDpiKbic5DJOte9S7mtGgtSrlptrZji/yn
cqU2jzrYBB+4yn461ofWsf5AEa0hEPiit/Nl2tiy5GwDF+CSwav6R6i8PPXs4zUl
y7CpQoDUDpbRSc6d0kIhRulxnZfcYNCZgPX7bM7yeUDnqBpWsytcHEE5OvXCHowe
ZLZJDU2ApQwgesJVyGXgZUKHtPd+PlK4ymHmoQ6G0h144ZRAAT4rTtOgo6X+R2tV
Dlta1shBwAV94fMXgAJCxSuNFMxNOxB91j6xNA5qxhP70J9NayVtlitgOSBMtLiV
QtGe8puC0h8cUHRbKjadp9d1XfnCMsa8RttdhVqmYNrYn0CC/xaFNYtwp1KMQNTB
x/BfXRBELjREfzy8QfB0C2EJgBCZH9ooTCdYX89TGECblnaUL7/PjCcXS+OWOpJv
jpmdMEV6PsqlIV5JS1QQp+fZe5PiwigM7FdDUjQg9tvuBUmFa8P1wFYlXIx5TmOP
PAtH8jMishtLGeKl8SsKePyDPBj/QTaPUWLMz+wUPRepdTaOc6wA7ZhY/p4+2Q1i
kllw6iBQ5s+vzeEatzzM2+s7nZRpUJMxROUyUT8N9O95sIL1ZkwtD36d2N7F93RP
xbDqyAz7xnlWATjTttg4V3bUuza0aZSHJQnmBCdDbWb+Lxh87P943D8hsgIJnl/I
wf+QTS9R/24ZeW94CpZCmEDfu9AiH6imEtxuFXy9gSNVQ/9UU7MLYON3vJUNBcOM
TDZ2aJ1jyri1pGfN8CwIAtttXWfr6YA+m5LIZgrOJUmmnfxduoJY1eCV9lHrgX7f
80FtuZu1BlPSm7RwgYjFVYQUTJTS7Gb5VAbs8o6yn0GMWQwDnx9UTKWM5p5eWCDN
R8FjcULvU/Ep15b+IqbCo0AUkBF5pMc3WLWat/6s2vO1JW/0pVWbJa6YrMO2e4b4
+gjqls5wPLjPjRoTe4Nife8fmIkrKf6TOOWjpxKVnJau6Lx7JeBGkJvDjoMHCA/m
+U4z0hUuYPGvcFcDpRpfQFUbqYnNkK5wWJAniokL/YnSt6410tzcFE1nzPaLvnSa
jCZk58TIakyGUvd/cRz4U3yF+iTFexFdVG/YekrtJ9k+bNKI7pjDuZzdpJ/uik3b
tvka1xGYqcpsoVkl5M+EBQE1LRkrOkp2+j2UzgzltL/SOalGviXz5LilCtJAzwfM
mA+0Krf5N9Ay3xtbXlNURTxz03UcowOm1XroubsV1g3TMGmolRs/Hg7oxqHj4EvG
P79RARXKC91fNDvQgKaUy7DgngVe5mnoYDwSpbpXWcUZ5OlwsYOvws7rNP+MZVkH
3dhU+uqLf7Wohf2qOr0Hs52OYCiTCCrpmB0/gzmuXC6K/vuRBFIOTLuNylz0y65r
AMXED6EQ0NE135kNOTgHeF9KEkSrwqhgY4QlWP1nlUo5VU5hW/IM/N5sU6QXyQzO
MGPJEwQnb0k8Xb2o/9OiMC01fjNw/il02KPv1D/v/cWNZIn8hjZlkzJahToH88le
86k4iPB8h1gJvI/or7t8E6PKoxciJV0ApDOdxv+P/1L71J86xUNL6/N2RFf5LKMK
3kc0zw5hswf8jxOLavcR5BR+7SYAvoWaMHcDZBoGc8LimJ6cZjjUsRMKX7XdslXE
0KEvnQOu2wp9UbgjSd0nXydc/XbQ37YqEhMcOWjwB4sNei05Kk6QK3+biSk2Yvw7
KOdx7WhjQq8Bm6z8F5OT/IdNwJA9XKFSQcFQ0V3O7WBrZ3OrmwP0sltL1V8Z/B8q
JbZfMWIVMoeRrmDCquU/OdDgKWpmaflfcK0zxSeaYL0xlORay7uhoQEHZuwz0gC6
rQI+YdHD/5dMqNCaumumFWLMCX3xpXudKcqv7g1OfRkGLjzCZYZccxCfW8IAfrdI
/Fpvbyf2N5RgaXc8g7psbSSuOqeoYyDCQb0gI0bqwb+nevuM9YK7w33VbgpH1vkG
zfFPpQwO9DFYADBX/3RsOL0ohZYdoDnAWag6HCrRgcqy1gGqMKJld7F+qBCUW/92
D/GPL3N8rPlbaVQ7XyJHosVLxL10yOnez+zTSfg9cjkreCYLznpwPdMNNU3aWaEU
iuHGCkr350myU/CYdoD8nRaLgbkqHhubaq50CQemcRQNJETZQXxRYUhqPekNBfSL
wra3lifaipV2VVVgDCoMRCduezu8nvAxFT85EJs2eElyH2SoG51nIMUylUK9918A
Zyzfn8j1G9Dq1GylXM4qqEN1o99IPRmAIpEW7T7FX+VIDZYiz+92AXWqqlJfHz7i
VowLLTjaT2y9RKyLPxPERD+pBrvjeAc6BtSmaFrJ99uiYiNUmQ20ZrTUvnrQcItC
DsVKR0xv2V6JOYMEIwyIn0WnwrRw1V8NlSlgCRG00HxXK1PyDO5mu4jcNAme/RgY
LZsP/50pRbAzSmVyoiW/NLYlC+91Qwx93scUQHhBcXdmigWh28DFKmzm7GpXl4wJ
9zFXiec4CkV4ApwJHeiRR70vfrkyYzyIS8sns4lneqNeTOy99kkHo4Kv1VGKa6Kb
BjGtSE3S2rMVR2D61LzY/M1/z6/WgR8a1fL1VXtcLHTJQSdc7FXh9XqAKNaVb9WD
7s7YZx+Xl5U7mCMi99t57v6HXII7/rNiO87SWXUA7KkJy3c3IKc/efVI2bsjcL39
YCooi3gtdz6iFXsje1SzLphCY2bmiZSnDX1aRJC9Aa+mdZfZ87VxorTml0F/tPGv
BgTt0TfPoKBvfTWbX+lAi79E9IO5ZUgVvi1AL1gyIpEkBx9SiO4m6N/LOSrFTjjs
9ikvr3txhNLuhzv7d8Q1ua6ffuEIl/TArzuRxgyxsEMAr/v8WC0UU+iQ5mHF1N7B
JPyE3G/DEm4K5Amniutqt6NhRCcAUE5daIwf2oG8yMTufVP/JuRwgXfsFmgn/BMH
NIf3rDfMTI7sVOpzhrC1w/lLPT43yFBp8RNAIGjLFqlD27acmcZbLzqwqs5YTBI+
eJGzc5ptYneoOS1rZQCkASUlQrBs3//iZ/LDyGkzkxFRDgUDO+3jLuBDkmYVgVgV
4DsCAQN6B+1E5Jnx2qUygfwxK0ZdB1mp/O+Rc2x/Z7yQ2w56Np+l3VqfqrqJEssX
67UBxiu/ODLWBuIqfBJQuUr9ALBCneXEHYAPZi28NskPjbCyaMNTOZBF8RQnwFnh
90C9KAfiBv7ELWeFbYCVtjmvlH0K+5NeXa2Qv1fy4UDGx4TQc8t1wR3gOXPB60n4
Udg86ZZSogOxhZnHTGW7KzPa2Go0UnUeIyaQCuXv2KcC7gges9yokz5l8AsJo3zm
1Yue7bzHvJe35MY0slztsxOTs1T93KraaItU93FD3D09GEuBzZiO0fI36nX9WpRS
u7eK4ebm54b4vVfMugu+P+e38AOZWuCM5FKhvsxH780SBn/JHIprgeUN88Xqjhx4
mm7p6ngdwgMA1RqNO1PO3hWig3A6lGIbUY5pHKr0jpbsv3b0FrcRIL4lQ0qvQFXn
FidfE0V3fIYeOg49VtwAEYX9R5sUR/uNtd76ldErEIqp0kTNsLGRi93fwFXcsBD9
CdehpTSH/DX0JdbbnUXOtTcpWjBYmCG2WrWnawzZ+RCa5CViGH0ybFFigWgvz+DK
eX978bZXizAnPF8223N/jLTLCEEAjdSnbFbqX57Y2InS+sPq4UA2XMe/tMbQXzOA
ax544Drqw7v6Za0nhTmjczOdlijCYd91NZtkrap9k+PVf+DyLIwyf+cOuUXBYFY5
/T0I7kq53uygFEJEvMaV74pYIKoUcYEyI76DMyZqmzsWKroDVumwMBK76NxPEKbJ
HOJmi6FeFdqieUbltiPX5U1z1wsYYJoLv5CTgRENvW7jwDjsMcui/68dBJessEu+
iiIze8gaCEQLqNRszfzSYsg//vq1jDlMzVvM/AiAc97f6LBXyKFedKefilNE5+zu
DyVnGVJsOyU4/ObF43Tmiq4q8ncxOsRVV683NZoMbb82rA/OkR0SbkWL8IWqFDqZ
4t1pXxFmO/evFylyRll2F4dH0PCV1Ze7ATeSYvCG09cEFTBC1WXcN7qwvxs6swis
pnBbsRDhAnz/W4YAO0GdGRsBDoDyIU1XEhsNWZb5mCktR/4WhdR4bOLTfBLObhTm
AeE7BZrdCuxdu5geyvSRu0b8kxKkXkdbkSuJsOxWE5lUvL/Uwtp6i6+4iO5+3b8f
UHvxbXIDKCzcDxleb0ObEPyaiSkAOwdnCIdu5V7IOoMrYAL1j1yZpbSlq8IM/B0h
a5kEuLYW38ngi+yP1JPLxVCXD8dGl6Hoxzv7vBsvrFzO9DRxdt29Xs1MmN2/VoXF
gD6U7EPoh4pvHx32HlhGgaACSxyTIjhnmwDryLDLsjjFa4Bm8S62D6OFJmlyP5g3
HjXlC0z4WDzNEJdgTwt0Ud4wLNDpaausNQgA2tqzvZjImUcSqH6PeYlC/ib0AkGC
4Oil/wUgxb68d/vN+UYoz19ZH1hzCSUVlgsKinj6mchOK9xru+EvDQBMlyTezX/E
pood5pluddiGUIbc2p1xQVWBcXeTJi/NlkAAWvujsxCVHVkD7K339QrRiCz7xIBw
eXprL9JHRugs/eW9PBCS4spduBFwS24GAYYOABTlBslx2ozUd3MFIrzdlyBqiJe1
n7ZqZ1ub/w+hCAP1geaENAvvL0D03rNrwV3aVOmSzuK6ETaCUfbvRxpUOMVj04Ye
kAkW0lF3bm7NOgAjVNQqAJ61cdjuUJzCjrTRpZUt2pEcdNflcX2lLE1k4QOOkibn
kpRYhGJHwxh8VD2hboKZOWHnYqRS/8ajRmTYLk/XxoWm6ZGGPEgNq0u/Yg6ruMYX
L2Em676cxw3fRioCNQdJd657n594HcUdQO1/ssE4LrXRfsZlB/urrQQxljwMiXTz
wSvs/BjBy/2x+5vmZ3Ewa3WJcF1z1zX2/hjMIqn/acAnhH9+FhsiSmGSPn/Onc+o
qFP72CQ65sSezxCI8Df5ysZJb+jyrDyCbnQZQ79wnBj88mE6TuOmpP7evnTIgnoW
DEQxGZl6y3aobGXJ82rrarJFxTd1oCeoCSzirnbAVh4IP5ludDl6VBW4aC9VEH2B
3rrAoeyvYJVouIPjePa9MVLdRwvNI3G72lNH8fowq96AknYE3DcxctpJebVZtSud
34hF12X6hU8DdVG615U0exS01s4lwn6B8HSTnpvl4mNuOWdUwsTlGsCCehruLnYa
KtGl0QvUOZNyBZxqSgZzwNt1pSzr0Q4EYyrfExbJ78H0IRRotfOeUD04b8h1rv6O
M+Q6V6Uak1RpEBmPa1JiJWDooAwmnRbDRX6BmV13ATsUfKS3LXBYSq+kmkvo0mxC
wTr0KDdY2saFVxPnrnKBbyoreXwOrc8OdSkR/MhtFi3ctqWq5ijezSDpFp7Oo8K3
nVzOvLAGQXcVygxVHDwzEll3pr7kA4xoeA06Q9raRRKkf6HFB0gJN6PXByfAlChQ
FApDerBbrF2Nr4cu7vmb3CNqRFJ6GeKF0TMGGXr6nRjMiZw7ScEhLv3CAgyaO1gl
SA6Vdf03loVdRLRYuDgczxjGbYe4op9EDGxoGNmGCYe+FNfTuHzYm1oR1WPnb4F1
6mvQRNeQgrmY9dtUqyWBb6XjtoloSFchzmFgrnBMF4kSKqqBnZVb+KWDxo/7hhKA
qV0JClFPq1ibeXo2aRdlJlRYvspqXuB5knvCNFr6RHB35sOg8tc8i8unHK5MuYCN
ujyM8vipYH+Y8aU1AyFQkv9VE87lfQ3nq1O0/awNYCujDTX+Y5I53QyefcipI3du
QT2rIb5UVI1jhnAhBexj5iWtMThe0oH+zoE6Q6gO7QtumcKSPR1asbwaaxAFKvYm
KMtw5U4Bo6HNNpMNw1OgNEogUnEWZ+NVfEFCA9zolJpqBDYMXBVK7e8kWhRcbsiL
WsbcXa2agbGp4xImDJ4hjG5uAGi7hLciWK69mySGM/cEUZfSNiiJ5xARixBNPsr7
rDGfWKUJ+Sicl1HgQe49ewY2Gt3HAtqU0nL1/h/JQNww1HFNLIuBrsQ+ch2XR69h
A3WbSZqIXhVox+AF2577KS7voaEKljEoZefF4m8XKudpcYCNaSTUyxGgXCU16vy+
AB0Rz2EdZ76pOsodSc26KwnLkUauRBv73MG5WzPKmJ7STwBUgRG+Hq7BDMK73w2I
5axtrBZ1nSyNix48SYA8ANsKJCDd1CewaINy2CJj3SqyS3vcDRxoU2oOz2uzg6Qu
0ooYLxqER1BLV/bQ8dT3Y53qNvOmDD6xdCMlnJhWT4GvzjAW6VF42WrwOP8Q49fx
xpoC3YX7ruwEIlBSitTedWsacpVgyGcgnB++/aL/mDhQYOBaoJLkJ9lwxaHgo+NM
jxgPQFTB3eecAM8mVNwEQzx5kyhkbMxWkEpCx4fLcXRVKI378OJh7xCApPPCmhxD
jRIjkpHq93YEEpGPDjI2kCmuXChCvNjYbxlreLjSrk1gWWeT1LLvHwxJAaXShbS1
T3JVhKZJ/cmRBGt6pVcHSBQVj4Y+7dHLOWYQ3/4NH9AYTIfH9Y6BhNROs2I2hIPC
FqfLds3ftsRgVGNvz2ShG9CubEjWET6SQVug2O145ShOjuCjc1+zZD+XmyNqJPqx
D39lxRt1H7U3Xapkbb5nsJzb8VM2O49xCMVi6JWAFgsE30/vRlgKl2wKMFcwGYGr
0xhEqaXVnA5AbFISHbZUig4P+VX5ns3PfDqXYa8w0M5gdaDI6rO7tIUSkb7NKqzZ
HntRycHPiLxZhPGY40BgZTbF2ONYdfyaL6reLJqW6PSU34ArZ5TFMTuowmUW28dO
4tYcmud3VWDRRtw6xOX26BmQBUUO1vI+git3+7vXuQ2cF0DFMHtjGn0lHVaZkKrj
Tg+Coivmlzpi4dcnpII7IUp2K+MBAAoqQkWWlqGHcyU1kIqAeRtu/D/GFejmXNGU
lT8JEib7nSUsZOmNifOFMBhLt0/IWHKHRGMadJBQ1KXkQcYnrH4CFqczq67sh1aL
DKfAkPv2osdE8gKnTlTDaU8PuKsUEzF8Yca412SBchkQAX7ojIcWCfs9iUGqAYGk
8EAxUfDavdumMTfoHJDNuvN1zLy+w7LL6nq5A1YbzSfLZw3lAKV81d3EAUVpqGVa
bbhLY/T5IjUgSmDguWevBmJA87dGr9HIZELbiVfLM0FMq1+0kTcZ64rlNmpRFH/2
bw5fB3JnCrc2OLqMAmVI6IwywxuNGQmBmg9QL78obgPQyIWvs51bbUHl7A57HfCW
qSdi+j5iMPjDJnAro4JcG2DSLhq/7jbmCZJqEq41FWraauJRAX3ocIIRjk3kTXaU
e24QuN9CTDfkYHA+sIqywqKGhYRtsNd/yNJY7Prs3hml30OU8o9F06kAQWaRnVWP
qudaO2K2l1iLxL7LrHV+yWHZ+/zIx+KNGPUm+T7YM/vajpolFPOdI4BOFl/ZQZll
/CIECEomIAsKeMbJBIW7ZqQlUC9ytt1N8Y8QTIvHoICDnkxinbTaVynjakaixRxH
YTnUyyVQ78cL4abIanejtNsSAB9OyIILdPiYXAFq9P3AUsT4wRxvby1BGaQz6BcZ
nDFaJEmvxXrGjilqCwc8UASF3f8/Kd0+idcMU9fi72QY0CoepAjj44SNujSW2hCC
LF5tmanl8/y5lZ59Ge4aWAynADaaUu9F00R+W1RowVE3Mbjy2Qaqrlg/9LoNI0qB
EMALwYLIfqq1kF+OGXZ4+4FcUa12YiqmCzp597a1X0OSEilZRkrJdM83i33HLmkM
l6Djtdhl1xB9pXTDK4XuX7Iegk69QaZD4EOZ55A28v9lDSa3wGvyhW8hezinL+7/
qc8sgBkJ9qGkynfnU4SeXIhqCJGa7DT1aT7N2WARtkNqM4QudbwVQuCa+Q3Y/qd2
np3xrH1RWC4PIJwgtkYDfpie2gN/V77cHq7u/y0JmC8zG2Vat/VH7mgyQzFHv7Ye
uyiKGDvtVJBZJ8VMzAVIfsT4SwEBxqakWQR3ubLTxmKEXQak1+p+u7VyBQtpTpPS
W2KARUyVvVgj9yeOblUhXTdtejjr1fNgf0Of0OZNtIwRRThmAS5eFOOpJtprz2Zh
SzRFT3Oa5/1xlUvCHp+C0hB2KFPVXgdVx3yjTNmtCL7FEVc/CgS9eDNNroqvHyoQ
KnLXnzwBHa0WNjCrLHIcCMA0A8GZSN8lHcA53uV+pLFlSVIImM0JMqM62txasM4a
aVPI/0rhUBvVVGMjQNSqw69RReashlh8Ev8ieh/iAASULkZFqlfb2zMg6vXItIpA
RXCbXDs1BzECN7Wdbp1s/SiDpObDx43QM5dwWXj6t5ZN4i5/UxR+0jhz1soG4C3P
XSozk6DjkeR2/0oxliZBlPdO1T6I7a6Mer7MRLt+wlF/8sfHfhYGEG45RjLKwklY
7Z9MKWlxknYW0h8QP1HbtgmF197TPGamP+UiC7XQGqBFdAlT+GkKTJQIViQez1Jj
Lm83sEoKFPmdOztC7h3hwvQHIOsqkOB7wOWWY4QmxWmkgLiWtHwlGTfyVMVmwcxm
lnYtZqEx8XRl/EzD1Gyq4uAXvuMy9nMMT6W2zmwPUBjDb1FF3enEJCTEW/GZHwXs
Fl+VBsXkcxbmOSCdrbRlwg0h5td1uf3jzOq15Dj55kqxCLJGxgNu9KePzS+iNUFs
J+pOzIWXESSQWdArHUDO4Y2iCzxN6rCfgStMRyV8nwPzLkGUTCniA5QavOAwfLmh
9ya1KcK0ruaaFkwlPQWRyTj51Rtv7pt4qPXxch6WDLKvYvFf1fd+j7Md7bZd9U4M
998etszR9mETcqq9l70JTmEYs4S44eVd1Y08hFRgoG8rYPTqLlY0WwZpGjtgJRAn
3KkVN0adV+SlOoFG3z4+np/HHotQQT1dePsiu8qItekYn13aoJIPOPAFe+49ML4o
4QP7Tl6UwN5wZrKggs4a6eGzv/a+MJ+A2lkqNMDf9+71hmwo60FTtcCNOM7Wo3ei
M83cX2aO83zEAln+EdhFKnxkn5lX/cfc8912LBpK+LUYQDcKt34/5Vb6/NeY9Qq8
PcHuYKFdUCeF8nUkWaT1oy5arWPfzB7rl/KSosWZAacJNKpXwhLkqH3YEqYlNAIx
`pragma protect end_protected
