`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lRwzq78V1FpDoTVD6WPYcNnhRTdHU3E5crAGGZJz/gIpRn75xqJmfL3gf8SdYrVb
YUXy1GKnQ2WwadA4EPBRSKSIvwvVO/nrSua9Zu/5B6CKrogMxi2w5BaHQq53N68Y
j/RcEjIPbeC4KefP5gYOcjDnJRRGnWL6HJLkxWjEfb0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50096)
2PETBU4j98mIolUf6KYLPDEuzZCCwpmoj33i5pEUSQtVpcpAKXwJiZ9ihGAJMDCr
zRcNQ5ieRf+yqSOO8of1fcG6lqcBUbcGAgPVvo4SI/8vPqtLfbHMqED8MogC4Dfi
kEFxpW/2JhD5xricXWMxb7D/IArRah4A7oAJlw/wbaQK2+XLFHP02bfq+/uAf96o
9pxkVckJP2mVg3X8FrJWpGG0DQNLSajrLK7h+tP6QrihfbIq2Af4pakjtfmvlnK4
dcFoXNmw04g8onnJUsCQ+B5iJz0GCeG6QICaL+qIR7Zq69wnpLwYxfj2zh2/uIAE
4jJZvkn/cVdWCi4NxboaqHonu8nAe9Lixv7eXvXI1Rw4czm/AuvPA8s6JPWq3u5U
8T0kIRVg+yfuvpWtWQpBoZ5MY6uc7nbG848oxedx/F+Wy2bPF4uoYCJ4Vfwm3uEw
G8caKwKJAW8FUHe4uI4RhvqsoQ5cT6yqJY6om1Rnmq4R/JR0twGt9cC771su5RY/
N4X7WKDhfD0pk/7NmzRP4ZBT0CQO/M8pq9YUw3I+/rZukxTQ8VgVY8NV1TMt/mc3
QO6KzXH9fcYkMOBJY3/FqmZJRyEIIlqkYwRtfV45ANxnoMNYQLX5YVf0Aw3g1HoP
yBBIgBmhcdevBvDABD+IMerI/7fI66VL9dZBa/i5hE37GutWYP4IT/4cAMr3yVer
/gz4AW45Hw9V9akr2tgN2Ev4M/CsHJwLwO/gYr3+ewC1UNwiSEcMbFr3sYkia1++
rsj0jSXhdkfxTpTITKm+9I1A7kaBL+jeGE2n2Ix+xlyXxGuxtPc9SU5MhSKi4mYn
tgCPIxehqfeaw71qk36wJ+P4ngA5zN2gjW+aGwF/uTr1t3h5CTpVplMPko9lKP4y
CEjhIyAQth1zCjI5pSia+/HEXKlTPrv5Zx3S9YlgTYMkK1xQYHxWiVRjG4527v1p
l+cedS8YKje/TCutMqBCJ/Hwc6JE+0COlT4iLZQ9txLB9qsje0GOoPcfeG/+vFJ1
+vN6OVY8U+OooQg4VuTRHURreZhmdYy93jQHo3RJHjMUaiyi8WCTn4Msy8sLQ6yb
z+d7TCZI9aXu5IAu37e9G5hNvuNbOBKe7UvzdNQRp9NBFmi5XjWZZS8QSO4aCy3A
iaKQY3b2/LAW13xMpAJM+PWHnklq07rZ7qLD5IBg+4OnYtXxHvUjLnb1aCRvMqka
uTYixnhgMjZi4UzYPPBoPut2dIeovrYGoJSLIhn/7motAOhnaSkN7bQPblg4pNVE
5T+qasfTJVr68hDGlSKRhDzH3hJON1TqZxD6CXuJ9XHPTr/ZANLwTguaL3sb/eML
xs7feKT3tyCouFEY2aW7N8KTfJmJenB8SrMCoQPyLKFIkI1HaXwsWyPHY6LK57sJ
C8A5Q2L/75eLNi7aqJPqsHUp2U96hbUA5M+Mu2TRTYYXdJphL4rOB2+/fUF31zxV
AdJBf16ROakm8UnP6DKuDvnE2lAnCpG6xUKVabtQR6HWtGhyyrZp11JGjaCqpLEO
LKm7ENlKdjo/y5nvYUyfG/E/YnJ4UPlGTdeY77UmVJ1aUx8hPZBlisa0BsW6IcNM
1wd6a9t34FoooBuMSLdROi+jWOTuzKyoTwkiLkcATa1lfWsU89hx7FZrvlsjDymD
7A/Dn/wuBZzq7dZgmteuMINdmoii2X2d0Ew6fTsAF6wKAk/s6ltByxh6gAksmxzZ
rbu3d5bn85pgyP0+BbwYw+9ni60B+n9HmulfU0IHh6VrvKEIohOHgIyoWe4vrf6B
GhxwJrASy+zNOMQeqOyzcoT0jEECSkIH+0Vks6AsMrYA/MtOj3LgVQI9PhCn+en0
HR5cuvFnXsTENqBS9ZjARWB140DsQ7wqyP/lLlTpCx+mOuveg8DqpNxHy8f/wW+f
lVhtcyvuOd4kpqdIXHVUJqzJZ1QprGDSABuQZeC0uNwPFE18F+F3+KOcvgz9U2IW
UIgMCaJZO9Qhwa372Mm01kEY6k92yIZO1Y5qTtiukMKIqikmxuZUNppiLWSrCd9C
1GXyKZUZkzInQY/Ap/jPJYvfR3DMAzhotpax8TIo0SwvluyatpGm6oDiLU786m4C
6HTjFCthlb5KL1nl3lOG0kSfU61Eru5gJXbCTx4Yx0zTGCmj1NCu/0Vdzkb+Av6p
w6l4NhgqyeVANpMFNLnlY/+UOkiYksKhIIhy+T9suhFERb27dAbLbUnp3txVmDs6
t3ivhRphIzQlZL0ebw34GOpn1tAt2rbXk63z27S3WmWqTDZleqLB/yk8NmosYm34
8SI86z6wyQSyxlxt/3p66eRTUb/cdmYuLy5a0isYYptV97NHi3Su+yISM3HlV1FP
lUJkyXwJAnKkDuzBVJrP/cJHezRaPbLZsSfW+wa4EVqXVnygCEAfvDUge7dde6Ti
4UEZq4RmV1NbnLNwUk4CPd9Lg2+Wm0i38OQ9LT5QBKTjPO9vXql6Y4Gwta5JUmy+
68c1/LIQxzGPrsIh2ZoUu9xbVu4+z15XT1YM3vkL3nsGf0Apx2KN12TagUyUm8hz
SFOUBmcDv+cNousIXyJLD0a4yf2j/SX3Qzd0OUOKIdepfaKBsoJ64zVswjL8+LbI
aMztT3EXIaStpezAEXOioVCEd+2xVEEA8+4vAfe8z+qluCUpsnw/q9tgSw0sqS1Y
JhoUKWS2hvR96fdcvUeA9YNzOkS2kjbmNrTJgI+89zBwvrpZWCMk6wReE1ndOazC
GBSril2LoOzZWleQNsdROe6hliOlVYrhERdS7GWct8AtdGWEHaIJNB6R6VjSCKCQ
qdg6pirAtUDOHrGeFhwuQMyAEctFyrohAx6Pxt3Mms6kTzHw2g9OJfIOE3Lt9fKL
UeWTxGLdlh7l1sPEGs/2EirnqwMpn2NTCelbgelkm6OJG7os5wcZODtyt9BdYH5S
hvhoTZZnWjfFYQOm0wPmY7YSLTKj9LkZSWsoHyOq4GQCf4MYk0vskDnKf+DNUiR8
cMY9BURvHDz8qYPWRu3BOqpTN+hYEP3myDbaBL8MbjWC5lY2IP6Rvq+ZhMAGcEhX
VBpoP7v5tc6krNmRetjRXHdZMK1k5wuxHBXhGgcVyZys32h+H4d24yECC+FneBR+
iD4VjFquY9MftxZqtrG85uJhcrSKzk7RfDhLyRjeJEjqBix788GZkyN7Bdt5v3/L
Jky+sAZYxQaEeKYSVv5dwjG+niuu2f9tPzW8Un4MvqYp1+/lHWtd6VnvaQxBjy36
i3BAmvwobjSmTrSKGu9TLFNvoM5OLsL6WgfuFurc/f8BD1J9yzaM+kN66GH+bgSL
do3EdhyOZLGlJn5iwyshKGFb/ked1HMZqw9VhfbNia9oYDu9neHL3ekopSzRvM16
ziUtkIFD172pOqkPQSsYQ98hNXISD0g7tLVrdsO9Tq0B2PfRNoQgM8qfxWRnqMWG
GMjT5ZVNM7cea0DKqJXjXBaylMqKFfNIfqrQ09rHY/2KjRfOkQ5Q+kmukoKO93i6
r5FoA5JtfJJK2Pf5jDBX0MhI4hM2KBt/69RHoYPBO+AkFut+8L/oy3WylWKR26EX
X9Hj9uezEPZNTYcjV5YUk2eEKcYbBuWMAzWzx6X40XQL/jvlShnniHVLZfPU52ox
oSKZRsgmFszQWd54ja7GHvHAKWUw2gdLrUGXfAfkpVmGE2vKfjRbltrilsXPI2m1
ouKAP/qQ14X30Kiyui4wa507JY1pBzfVQ7jtHTJayRJkYZilAWWmMMrJBq7/+pwR
c2LrYbUvi7YY95PFbBHdbDrVotz1YuO49lPYD818KK2OEgYO86BIP4bINbsNYBrs
SNwxH8rpUAYjdLhhMLX57GrzMOpNZzGOcULLu8jVixj+/hVignE1a6cdiuSJDhmC
/L5wnfrn6ZiKUZrqsfID6AlcNqnm07LHKdIjj4keLxto3MFq7LDD0i68z8fQCJnc
7j8GH2Z6D/uVo3HHQO8nFE0ZsUSSCrIQPkYh5q3GZKH5cwTBGIRwvufmx9EtVWB/
j/zZRRDHJGi/SMXuwJ8V6xU2eH6o/uy8wNVhU6lwJ/EuxLdCxqumetqtzFHUXt47
MHHXvP9o4MuH92ov3AS0ETHZGo1Ib4eaDAOQTNkqclW87cHfn92YfXsF2xsfUfZH
S2m+HUEh7oZy5KVFcsC+M81pUdXX56A7d/KYtfOU6CrqZYEVKEYcODWu2+/t6NGc
j5MnbOoQ8XjiobbW2Fg6uAvEStTnJ3iJo+EDZsW+UQ0FYL8WoEt5VsklqSZrOwfQ
A334Fg9kdCC56BCBhPUSXE1p8VfPvkUtVWH1dlmLVFR/LPlHtQtp1lknPCd3f8OT
F5gVhz2NXGJ697Ezso+3+4pkD04wijRfrhKya4YKZY55KYSSKTL6OROPdy+nKBgh
u38OxNwUcz47eF0W2pA6qinNM0gLCpgZk79zxVm8dD/cF4M+893fUNKkwvbmU/Ow
7FKxDrvFVLPrDmD0k54Zxb0FJc5ZF54KbDy39in6AOGoH4EEtZ1WdBeU8LiXhODw
RdoyMjcJ8Lsp9yIvtvvq0qzXegWCUH7ZD0ImjBuTrZcwnvBCSjVJ5WpvsBfetKBz
iC4rzvYiYQ5CSjTVnn1nJ+q4LvR6QWYR9HOsRaFhfOMT+jfyk7CJvyFugU2BokPs
ZmTPknOl9o5BOiDkhv4YUyivji+eFiStX1ZtsaEMgArXlkAXJUFzdmKLwW/vzIhq
scSmu5ItPu3mvMav7fB4F10Pasd0YQ1yhezS5rpksA5gxUdyq77bTwPwuaG3ENYO
nYdnzKKkRkA7udF9oHqWklsV0gdHczZBLJOuSVsjYfrsW/5yQ/H4snFemoeooNkn
a+cR6aeJvB+vjNULcDkI3tuKsKxHrSugqWRk6uy6xMVXLSLPw+3oxKauHuvr7zw2
zjrYp1PsVvLHOsgi1DOLPWLDmfm1CtwXEUPNHIanOlAT565peF6FjinzH+LdlFSC
+dutU3Kg6jCDAydodKnjOpokTc3vLmNMQd0q/s5RDikhhSGPFTMtHpKdMAZMS4UP
YVDBais3Mpes2pov+nP9lYxnlt0aOJOabHWdYD1AvXCppc01/8kih81Vxe7jKWbX
VILe2wfX0FINRPIm7Q1NJhxydNjjUF+LBjZFGOAQ3MsGS11B0aEblWmwJRtkknEn
oYnyBYAUME4RXWrAYw6GFm7FYTCEUJxSGuABnLuhf6cURJLHPYG7KtX4XexlIBYa
aWJSMm8Ag4obx2P8ogdL35YCqTlz/H9rSJNrkmpdytCRx29Nf//P2NHOYKQ/DFYH
xHTN2prE8wWNG5ezrLsvsMQWQ/CEbfE1KZBpuAOLk6lbuXINjBypEk4vIl2K8gYd
1CW+8eZ//b+5saI4+e2TvwfkHKdXoBW7ELp+soPeKGQKK8XpND8N+YFNXSkCQUFS
cs1uuhPMlAOq75TKA+S8yKYtenYmP78PPyYVBef99d9EfZjsLgHFaedjRAYRIT64
Xyhx4B2F3KWviYICUfeoqy/VoZJ3zDaicBsJaZpBt7dudD5/juUYGbiDz1f5E2Sf
re0+O2w8dHx0XzUXwlhhmLi7462m4vc9VzlbP4+MCFsnVWlia7UZ8B5Tcb/95oWE
aaJcaC6jS2SnkX/DlVkpsA4oqSNXEhvTbNbv2Re4axONYIgjCUFA5QrA7Pxt049Z
uwsYwQTzHZEQtGm6tnPeaa1tXAFgNX8moxvk1AoxcGyICGHl532YCVQvtPzzfEbf
LSAGq/4Y+/1zMHulY93NnqTMWnEwKsmTt0tohIdjsHk66fK+ADpVDeemCHzfP+RJ
QMW+NA6hU7NaZPJ5Ig/2yQgmzhT/jw5mRe3pacqqZLAwlemfsC/bJSFvTiBw1W7E
cVUQ10cBXy676jBKApyii0wUEe1glKJ03Q0SWyWGhLQxhPkrOoL6P0hsMjUJKHZO
pC3zsP2+5BeTYyMlNf65r8g/gBbVprfExRF7/Lutc5yrwJh5XshrSDb6gsR04c4+
5GncKhTngsf28EsSAczUbXyAzbWfPHeZ+qudT6UAXNASRusdWgN2492or6QLIyk3
1jlliV0c20FUgia4w0AQius/vITgkFv8cE7m9eSC6AT45Taeu7P/fjIfQAJx/Rcn
16HNgEd5ZVipnqBoCDCW1b0F2IkTiCOP9Z6rY3pFNBsec6VjtEAFLmwE4ydBnnNH
dRlkcQzdIM0MthQUxeJybxP16GgcCsMhQhmcMne6Mfa8CLZIo4IBQ+y5Gv4j3luG
HhTwmCYtJYezWozXJgia03g4P/M0/8aDri0Ls6y8ovTHNpSvswPPqE1GqgMaQFR+
Mlt8TnGCN5PkiP6WVZ/cBITpnpWEpMv8LnakhBYNGiEbaEdwronTkBcEvv4A3BhA
FUhGPKlJMCKQQVLBW0IV3cmCZU5ykXTPYLDw+rbebwUbP9qBhA+uqC+iJ7TUMed6
II0dzVucELP0EwBgTnfNeM54BjWsLZIKrhK5g3jlhpXgXMlrJNwNmZjOpAlIFfgh
S2UsWn7zDcRz8ESNL87kD1lqyy8mGnFzrIZR21/r+krLyIdolocQRfE+9Qmibcq+
0wxkjNIiT87I6lqYDUMllqjpl5mKZ6w1dt5VE7R3zjRe5Sj8gGPZz4ZTJJxx3bJN
Es/3IdqqH+M3cCp2zKJoV5slReiHyIRKdApotb8MDVqfXD/FIGTgNlk825Rn6H18
6EwdEKaH5w5A9AP6Vk8517liXuWmHqc0y633xXqfusj6hCabD0qcsPkM28yxL4Tp
w/0xbYN0m4SqA1C9dGVJPpvD5T698QFKKrB0KClXvoqtm37S3VYyDH4P9TGOs0LE
1fQZuEWbakVrGwcTnMrUazX/hPAzKypF4MT5WZtDPDTnE/Z+M6rhv6pf9FpfRtxD
9TIz3En9jEQpHfWkBKZpGbwUFqKudJh4TL81vICjl5/LTvSCLoQS/Q+u8qffXHW6
UUE2/Df7MjSXTYnknWk7mvJ+jqLl8V8Ia6FhxxkfmZcHyOsfIY2s2D3fu2NeYIua
tH1wEd0gULT6uK4ZAqCuggW+HLvsJXJGZGzk9LwcvXcdWugk39r5zm98fVpLukaX
WThI7ys3WEpAn/zSLYibEeEbwAc5NhjbP92vYo4mw4q8O5UEyETvd+RyrUk47hM8
K2wZTsb0yED3aPOqDox9Z+/46NhS+EjeXQGv2f143ewAOzN1/zcm9foIKJjY322R
ijxIz2PDJpudZbtQJTTNovSpWJ22vhQ32AcHkkouLwlfMQ1X61ciCN/AfUhiYE65
HKTSE1lrjyf+7XtBd6ZPe4IEFNpFCt5CRxOfsV6VpJA4+1YFAc/pxXBC/zn0J+vF
KM2BBe35+q4KL9df4womZdRz+Rh3FA8OEUFKvE1A9wnBdGnZBMQNHkVjVoGjB1Hw
/YzS88d1D5qBBq+FMtpnEVPgA8po9I2OOW21XdkAFw8BwuLIDMBRpszMyg72xi36
qSfnmJOSKsAFPWzSVeYfnjxLFXHOUz0/MndGZ+QdRy+ocJFpQAQbcsLyoi1L0zXx
xZ0JcGJKByofaOWlpSJkW8bY2iAASIJxTV+YFC/l46lTvs6oUeP8DRYCNzqHMEwM
X2YBO+J2/JWH9p6lNzR8PEgQZWaNu7lsW4v6JOFj/4ati7E1znW1+D6qIzTF025V
Q2/3323UscWK6VMNoi5xX07krTh0GGrb2ZROzhmm9aIcF9YTks/ECl3XiTKsFpmy
hb6qKZgdwwPEEpaBzJOY06pFLsiCyGbv1ivfj4NiZteHTT1S/yQV1v6JOmRgyXks
Xu8Tmj0O5AUaFEmDm0yhLos8jlhHvyqdhBIjoTitIE4T/Jrrg4GeBUpuOyirpxt2
UM3Cu7m3rtDVjqfXDE/g2OjAIgSAvAK4KLhcr78FJtpfXZDa8HkLeLSlhC2Ndqb0
aYqkWohaxd5Kt4oVidKDyz5cqmG8J5njkNmPoC+P0B8V9qvYilEQcyoedFiEqk2D
cbU2/iNsP5pJ/M3cGGjAK8FzGRJK9EXfO4eWm49O2/MsrlLngYTf856CTaDet98D
vMQj1nt/l/hj1pOPfxgsiJMVeUx4sLNZQ/uQhb/Zn+Ubba/6XweWwLEbXmmk13ej
/l5wa97m7rNUgMn6kR+YJNRQND8mDrhEi2YR15QPwUmnvn979OrxtjVya6u9wnU7
nWYZ4rW3sMWbEFWZW2Q2axv9XN1TdmAhGUvbZt7Zhoub37hJSzH6u0+iDch5ZmMn
XQNcDvB7Ql3xSK3I52PLSnEcMWwhDCjZDhyufUZESJr42Dk/FshePNaJ9iXG3WDy
yaXmIoF6OADIyWadP5eBueEetEYSQ/EAqIQwgwqMLNx7WiUiyosrvAKynvLlwjIa
gJFQTf9INHa5zMTiehRX/kgfXpHtii7cyAFK0ObXw0n2EmKWMsoCEZoikagHqgJG
nfZM5mSWIBRFbsNZCgnr862/CsZpWyTz7Pj1kL/9C7S+bm7OUuezyh7ZMtroqzCe
ZA7hztYlj7H+akRlF+NW/ZigwKbW6qfi3Kdn6qgcS1wJuwiw1P//DYWg8vd9iEOX
PuHZ48drO3q4DDsyOYzDecRlN7FPmS2VFkDRmeo44K2ZSycW4pQ0S8lfbf2nxiWg
uF2c3AHfBuNwyeQRQobAFdpvTq2MpEjvnZqAj3Hhj0c4yd6tdcTQ5gGUZ/XoH0Yr
8JRrR8Y9IEQQG65nvWXKfU2zpovv9bs9yOk5ynOh02V98oIYWhhNLcWqW2w+UvXM
YfocBICaJdxqr6n1NTV7L0ByS/d0BiSm9fSDbtwIunan8rUAF6IuwxlwCoh6A4GE
j1yfmk1iNr6QxPAZygJDKvxTUF1EfazoDIZ7H+AVh50IgeuGRIg70gMDgPPJswvN
wJPnQosnJHW5FP7eHeOK9vdO8S3sQ9jVS0t964eGOkADCC6hOg6m3PBgZI0EbXhk
b08gpwoGPI5lSoeqQIyiPuPlL3mo5QrXzfmTBQ4NOzdR0doDvgJmPDVWRDSG+wpT
urtRGL1VdhgrmPmN9RmNscN5BMUFhnvqBDmMtQYFHsBykfOODeZO4osW42ZmwjAY
iN76VHCOXAU28gIoA/sKXo3jCNQ7SYKHjKi74xM0rHxF49PjzyukutRvX+f0ja2E
Y4ampUsX6+jEAH1cR92V8Gy7UtE/bzhD0AoUs89xMmJ6gs3g+KNFcvA7BGJuATQP
2QzHHZb1plwufMdr0rGqBC6tZ0G9OsI8H/CaRzd7ktVRoHNbCZl25NYuKDmnTNdJ
KkK+8bLttPG8rJwjLNGnMwqKx49kDNmnqSH4Fpwwnt0RhcxTAijJqZUWgsS8Ly4x
b9GnnR0R6nnEFJHHWWS5Jadpas8HZpoYiweoQ7ZEC+FK28pQ/TzYhN8Sq2LRXzvC
5BVS+X2G1BI7kiCBkyUkIFBFVctgtLPyB8At3m2R1tcVI13+74bXNcLcHzorGCxb
8zZDBS8hpmOwBox9dDnecrwBXKmtsyJFZ7tyL/C1eomT0z0iCMi6PEou1m2Ri/Ra
57/BnepvmQygQDGRkRjk4vSz4tNr6zhNuSK7/yMbXeqpdsbBI3rKNTySg2Ul7RUT
CA+5BvO1g7GMnIDa1AX2XQTyBGreeiwh2G+J3JFWP7H9Ew4umOFQOBVqYZ9dA0ok
QuL8/uey7IJvkuY+OFvx2DwAdPsTJuxDJUvPwldqf8j8FYw6l36vH3KER9jk6mim
RnHOn1vQ/GsvUB4yQdLdFNjGDTeK11h7r5DRZsMrGEqgIjTgjY1eRY0t6ubuvVsQ
z6IfokhEwMiZ4yvSKH8PEC68K9qSFzV3JAHA1ULe8gW8gdQJOEntWxxbpMkBI/VP
R1/ivj7UHRLIB5tlLYyJ39vAOBcxqkQq0em/giCMOuXUQVRL6a1ar7SyuwdX5jU1
K4Dp2/KDWRN7eRoEwkR6mBNXiC099YCzqOlJIxNOg0ZJf3wi1UQJf8VjO8tVLvF8
qDmUaGPIn8vFjMVPCkoGa/uwu4ULd55SVI2VAiFddmalxGYFHnBtdng6h7agxaaT
1xGQ1Xm2Z55H1/x5/vi6pfzS5hztxLAHX9zMWBzJozA7zfS8vWvSfvLs8SWdpUJH
2r6p5lnBV8gzFaMq0nUC+osQwqUHUV94Cs+C1sLY5Md6p0ml1nf7YCeL7uHJQ7vS
Ool5o2xlBS8kdluyDY4QXSs3aY2Y+EGTZHb5WXgzAplMvKiNHtDNB/sxBJdphrLJ
i/FsXRCTfrhtbUyZbZGQQZtxmgDAbtNnHHxJG+NYydfKtOM1d6ha1DQ+u3S7ChFb
3qN8G6NOD/Ck2dSVi8J88AFQMnFgCyvNu6IjLf7MATKIEsyF+QZF1vei8GN5w0UZ
6FWKBhghsodicqR8ylEv3mY2IZjz31sKCI6k4S7HQ0isI/np0hRMJHYslU+LDUP2
L3ELDrKeL+eNwYMPOs1FVrVWOv7GxiOrX9noCYjVmTtzgZqjaLpd3LIF5rQzoKZo
u1We8FPIR62C9XMR+ivco7F69Pst6jvfhDBr8iwof5os99ShDyPzSP2fgjz0if6n
C6RXBJtnmWmet0HrtDMNDctqGG8Mnm7tIPDiZsnPgMghxtg2LiNkXJV0ltpJEQFh
ddYShx1RMKA4qZOrnToIzfWDxGoBDg/2JM94GurlrquUtl7obe7t1ZrIUNecvLef
JL4SFFyG+Uw0yyjUmaqxv93jsJri394ViY979vjZxrwgzJ951NbCRjC1iVaFHlWW
iGQZzdl2xOevvmwM5EZArUynysCnlV/jE7QLeja6PAsVjN4I4FceOtGawIMrfdF+
fs84Blp84mwkJPANjMUppfgihmO3RPea3EfeB6vz2LVyeW8dW8+2CoPHdTFctJPY
xS7FheFXIuek60+0qJlWh7lZsBmkBqwBPMh7pLPYvRGY0nB8RPvY1BcPXmOi/RLN
T5p5EHC7awSVXp2e9gfBqXgHoT27IxGgN7rapz0wQWlAFTqUiabI0E1nLY3C6Keg
JoTrgMJJ1lnKdKO+nqkwHqRljSE8ppTdS/vRMpyFhc8vOew8ZIEz6WyXlIua6r7J
XPKuJwIpxH3DreBE8O77cNuj5kl8jrtYX3mirTeBQR2Ijs/vASnv5H7PzVFRpofD
lT1K0IFHjgxQNyV860JZE7+1I8ZQDkh1pUr+BmJ6cq5tzJmqtLV94n9myehur/Z3
HFPST3C5kXp+kp0NDLe46pan6UJdGcedoBc0Y8k99QAp9WR1JfbifvOIau3aIl8a
5VbUwVF19GRHz/d0DOC7uePb/DGWdTGd1cRvPAPePi9VoWMLnThXkkWsccgUiZKs
tGMG4LF/6ffQgN5fUlPyiUsHS1sU55DfgP8EsOYIWsweJOLQb0SPx/TOav/tfW/x
9hCEV0Y0FfNTyUFbAZjxZxGtWgBaP/QIWpUDPxO51opGyUhxRwYBNf2VQZzb2A+C
umKrff8U7q0yes7k7GOOeO+GeWxh3m7mO+b6Vg0YoamEyI1QcxkILoM4keOjg2LB
vAwtb/+FR9bP9k8TxGHqRUYtWe3E2CWvvid6fksy/2g8VeQ6K8FM1+ecDGZlqqTq
K5mtnPvWe/s49vb6Sjkn0+sDBvi1rU5C0uhAntJ8BQ3CSYE3VI5t5LALJc3RPC2O
1FhUAcHLg4HLEn83wL/pfqXFJzmtl8SH88HkwzyAuJUMHUUpjdZ3wc2CM4FfCYDP
DWwfHFd7uf0LqjqYaCTyGxtkBjulIoGrkZ+e2gMRwDba7wNPjjKHZo54UmNJ0TqQ
cNNDIzuCJGKCreaTtoup8Dodf0fpWLv96k3ku2hGSzRFH1aFgm39gBOFpgYL8PrM
4KPi6mZZNH5qbQnLTtL/rz9n7G42ntbqM0I5+GNKzF2TPe/Iqgb6+bQR6wG9qcV7
g66+Ra+IbwpIHintQzCMURiplR6ns37s+nwkBlyD8r5+A6P8xFKRHNUg4MDkXpmG
WQBhLEzi8Fddp4X8G945PZ/jUl58ymiiDhajmRqW0H7EJioBXBUlzCpOQdx1moHW
OoVQvk7EjrDIZcS1AlssaHr2dZ2oWRBHxOFCQVAoo/KTP9MK/AFlDGR0ctjJzyDO
J8P/+hn1maufQuwWOI/Itm91RnUwiACvsrD2ff7LrZPYRVLrl+E7+EFjrrXwFJ5N
yRYNM/JMREwp/ilp7jna6We03YD7dR9sdomVbNNPWUcazCMRoINlo1xl76WiXW1z
7LUtFgowFvqNfdbJtFrJAZp5HgdDu04Il3agG3+txOtr6u4vUUboD4gP2jO0UXWn
bJ+8LcHG7HLwvThQhpU41oCBLlNyNV0M6rsDgmkLiR0pRwiQCyVWOrz4Of3qJfQW
PzONXg+VgcPz4ntnC6JM3iMsiBXPnXrT+I2+FP7+LWk8g6+PEesk3pdNpw3uuMOW
NaqS8TGYSJ3U4/QXsniJ9wUFT13DoFvXJ1CpezBIYXmwHlViRmu/qbGr7lTuqWKc
zOUUMsMLIuTE2/r+g0VtgtGE2ntcsdhdOAvhdwIEuglqSxYQwdg+QoYO28uZn6qR
waB1oKaeSmuc3T0KAD+Qc0sOkASYA6nxfMn0237/CzDi9R8oIslmFfX5TXd+kGA6
ljmJlnr5agE+APi/dOL833buvwFxGfmVKoera+fIkqSy+TaDwwjRskNbgG2gVdpZ
h2QOHCesmXyobJUGUMxg1lUJkhmM27LmqPB5mEwO65sUasFb8xBso2OSJzJ/W7cE
FBOpO40ASicAUuDvxSM5WdzkV7pGNNkhF9BHQDUUzi4TlAj+HFDRWkBqoPcyfuOx
VCMnwR0Jl/rTIa1KXxHh+hdLv1KpAMYXb+zLUeLws6apOtEwGrMwnPu4hN065vnS
10qcRIgdiI8KJ6MbaBfK0fDjug1dUQnekhF9zf9JIsmtGUSXJMcxknTgWFDuNjzG
2WOmBdW14XFGLigYN+ruHyFv9zKsoYztZqFcA+QVYhNlZVRd/bTxxEwbdYe+qDmW
EnUIpBC+LFojrzx3FIrT8XONQcy+8EdZ6dV33t8C9HZaMtXSVqwxAvH1BtjsAiOa
+pOEz3GKtWb7N5KN3NQSdliDZkCbhANgK8cqSqCneu5Jznb4StmnKrpXe7qu+p4x
l+ZaQkRmFdjiVzHhOjb98b0NomyI5fpkJNKuqHw9grd3NOOia7youz9fNz2Bfafm
KSSA26f3vB9mtCKKeA4qzjcbUqncQDlz+QWuJ3YNSzkKx6DxDKFMAOPxlky0eQ0w
r2pS6ogr0E5p1ubYqzuWOeFS7Y9XD3VVXEJeLEqIP5ZHqG+0WTMXemwRwSQcESGv
P0k+f24/9bDUUxZB7/zYp4iDOuWsU4/HZHiRSpnq8oIZkgG48wqqvpP3qwC1MrBh
uUdFH7kPtQRtpk9ogr393DW/JniEwIwTo/r0yYs94amxxTHT0NvApzdT9VxlnIIy
cLHAS5Nnq6ktNzYwbhUHCUj0KGZjgWEinTjMiEGYDdAGQmADcPWXuqK/vU413unf
M2Mg9CQGwEjv+neIM82rljjQmjvr8pSKQ5n7hWtgsx+ylFggmUGzZ2yaD/USkQsj
uIHahL9eZj1E9Nnn+6nfuZ1asbHmcb3Z624QGBnxC6C9S12ff4gyjYFNN2ChfYnt
ve1hfF211+dIMJBCWrenRylP2IhiS3VBPtLNTafgEIzvoi8yiRaLsiUn1GDmEVbz
StC2abDGRMqsYyTSQkBXzIoNwIYH0ooPYkWyRu8EO1dVzuWqJf88eC8CUnvjKKan
+i6L1/mmN8D6C+o+Zd9ewrShHNDRev/kZKGHn0dDtH59bI1eJqwzLbDnXCyfM5Ly
dOZdaW0ePEIolSSTj7t03hUZ/jRr7vIfsjfaNdRMPRGsMcBM+d+PhgI4lSijpGcU
PUuYqpzuxbJ3pMdfedLuk8k5o6weeLIN3No4meyROqmAUJ2HvHSv4aQYnPwp4cjQ
TEUehBz2SPw9rp7CLcllI4U0rl79i1gHTpiz4lLTC+iWe668Qkxgtw3BCx4d96hD
HqiddkfGHc3C5tEkKjroszGlL/g+S6yLPyJFmN1NQDV0SGTvQ8WfS82rfNfyoBE9
RJ7hTtIkzCAAeViwGCGKaqMCACqvmJ5EP2NsLmRb1YLKY17mnI1TTcNhF1UE3N45
hrLio2I1Xh8S//v50MNlp3XgvllThkr1EOHki04WZuZBhgAQe1Bg/BnEfzgEtfX2
T36SwzhdJhk88IzBEgjKR7KuzvCG+fPvmCXgpbxNHBHvkencEpgx9wEuLJ4MOt3M
WswIk/vGshEmxdVZZX2URFD6e9VAAQ8dtU7WjHRiie+CHgIGQGZL7gQ4XXoqOay5
8gI3+q1UQ9PCa3feKmAbUwXFVSuZhE4mZieaLJJBiFCEovr2NwPc9Heg0D6TNHXA
jxFK8P1/x39tKRpct08wPtxOWSIWEU6TlVVwNbTr54viTuOplusYkb5jljVpF+eM
aoLNU+N23cxTXYvDqlLl1Wm7GiWZWUst5z9YX5bjnOiCvRcjYttZVS3g33s1Rgjq
w+GfaDXA1266DoaCX3eIQGuoQ1M5V2hitFNQScPPDUf7M7FyfUIY2HfP92Po6bqS
LJ327jwXHYO2XuBIWlvnnlIJ8DU5wLmmfB2RUly1yFBDO3Lfytz4oAXYftx3Q8GF
I+77doUMJKmxBJGXOMFF23BeNeDUTXyFFzuK9u6CEfzXoGrwiAzQIdI3x9v4VWQu
2TAiKbuKZSHMP2QXAAk9Mfs4e6B7m6WaTl97jnDMDmW0kWZyssqH+4LZDhyvKBJM
ZzCAfi7wDDdrgLUyxUd8/txuvdWJ88UYKNeBifNrateC1E+XZqLqSJ60xatXoYFi
TJquQ6XtWISyiQ8J1aWRFBLz/SnVGas4D6GcpgL3CX2tcU/ykgUW1SH2/bfBRvk8
25XZ2Lq08RQrDY6YH+WLORvHi7EHCFKbZe6doIYtxHkY/bdqmDESp1t0+lIlaMhX
rfA4MnuRYx35oVWesEFiE8+Tq5Li3OBeBoSEnqdwoiy812v+Q5vU9RvNPRsjvbjP
mzpqgWfqEU3DyGLefQuQaXPSfan90Ue85C3cQXqParmKk+5pnosWie+QV5AV5/pB
DMLSnD+y8K8VWUQaDLyeXjWiDsrbL4WJDBBxE3QjfvcSdhouYqnDhQZ+uWqR0MV0
d4zph//hLzD2TtvYXr5H4TRohKcjBW7l1+axylNiDRvrhK3VHBBfghlnPHUBIyOa
bi7qeMKZ95jsSU1jpVcX5Dop9+gfeK8cAmHZXeFvsPCLVzLF4AAGsNNeuAN2Ct5f
GScX8Q/timw3E/aLkK2tITJRDlHRzaDnwGmtEbVjcWlrhCHTdBOyrKTkXZQrPY0e
ic5fUKX8lUExZtVCh4SMllOnPeKbmuthLnXC1u8jhVTZRQE0lbqPYnSe1plo3fP1
6S1XeovspnTFF3AdoUINr1HoG55LrUwDPs13HOiLYvPaJxfLE3QJOCfhq9xExeVv
ePKpQ0RpSBMmenvzjnt/GBqKv9t+Kizu2Oqc2JGiVhYOHCKGUC2ozTs58RPKmRNj
CCcbYbc8AM5Xx8bG1mkwczAk+oIcOydgii95+T+HMwsvmnsUr0qGq5jPO8BnT0hB
aKlBHoRSFOKN17ZKjDNJ9QKr7uBIOaZFliEv8QYGLrr4VzY5I3E5rskcGl3cLtQw
RGO+tPrA9bGMX1E5AN+/fF1CCyshGzi2ssy0D5OJKfCNOfcprdAobP0tz5ddBJCO
3M5liByoDhEx58AM0q9GRPnC5TleWUce5Ggh6l5mtei6cOrk+XSfgF3zll9f3qSu
orTgW8xZ1swo7E/5d7veL3Oh1tCqVRiGLlq3pZ3pk0vtjp635exy9qaUMJ56gC/d
VGsZ0pJu4a7EMEPIyYjX/TsMTkwcE75raohCExnt/K778EEuhexNR6AC2wRzL7IQ
6CzYpf0KOO+FTFWVQ6BrT/7FaNABGB9eCt1sBPByVEXxXU5g7b6838V7PuqP/Lum
PMnfwpbv+t71cT+aUWYvU2S3toe+0EIGpkETwKIWkDahcxTlxiAn+ILmQfUPQRmL
zXbjy9w2xvkuYAqWmoXcKMQEAJuREjPVjA+g/IPRnZi6LNftPyIDpjZdH42G63Sk
2zfVAuqwrNyEMCYslrmV37/b6v7OwLMG086oQZ6DBNd9z8UUAs0KBYERXZw9q2ZY
mCzI0HLxUWuiVCOPMJaZ0weZXxKV53fLPDlqIt82elACMa8wsMIvNNJv7bN/baiN
qaRCtzJ+1p5CzlP1am+fRK5UVVMHk0s4doZHFVNoiJtKqRs18G+aVT4d2ZZ1Arcn
XlYN+gG8nyOJ4juHsN9nf9FnneHlWBxCCJs3x3t5DMne/3fIO9vzobe96MGtU9PW
oLbq5vYBwkuwWHG/i2nlGUdyWoUQFCmBbdMXvn8uvPUYO9wqIh8ggUnQoUJksxq+
yDDxX8oCxp32yz1RxXR9Nbyl+JMReIRvsmtY93uktRo9thur9mmuwaaxrNaCvB55
c2jmqr7kdz+cE+5wzGiC76FkmW20YHAEuzCyiozCn0SlX69F6FEkxhCnoPeZ4Sm1
mzCfqNfpWVG1kyN6WrdMlHwoeu2qjgK+kTcR/rfEmy652qkv9VEbsJb+gR/Nbje4
S8zbDrYwTfjO/vDgL+C4sFYKUPwCUokI3fymnR/kjbS/KUCpJ8UVm+R4NUFbldL3
4agmvYd58L5T4rPlshWjy1owmaVXyz/taFOUpr8HK2It6fZ/zxQS6TvgjqQ7NKvs
+uWqE+XFnfqZIUFkVZYcEuGKBbNw3fpHoFuWP26tXIzy1zBYXXXCtvHizr2bnfMY
cb+Z2e7e9OdmfUBAeL9Vw3oqRVrgVdv/IScNk1wXrw0oAqnB7aqQ7/I6Vg55n5kK
EZWlNQuve8HPoRP9HrbduSYkY0D/iDZ445oHclVmlGMb1o6MiHiJ1m2AYeFtzTan
89oGRfaHjYnDhP+qGe7ERC/nINuS0z7SZrPjYhDvt3YhrGMiOcPNl4kP3OW7suSt
9yfVZg+WwW4NNBrs/UxNfxCkdYtXGWFuPTkLOYber6sQ237H2HBLVuzqLgXC/NMA
T1FWqH96firOgUXwuYFV32ON6DDOGS4PDxbtWwGCK+P4mMCKUr3zq1XdBm/GyeaF
ITqZsg7FusAPvdlUEqYl+K317LMroaiqV9u8vgHQ4ZIXZANZ6LMD3dTVTog2bcEH
Vjow5026wo4WUWC4+XeHaLwBHbGmsrAAFDcPMTphexIhnxUHtofoALOanUMhNQAK
4Db7VfmXzwUu1cEplXBWnT/NsaYJDcfn1v6fo1LV/VofXRma3L0dCYpRK5CUi6Sz
7nq7wynNBv4g/4yhPFkZHCz6GE8kfPwu6LRLqnBUxIajkx7WHNr5IUXbmUns0m/v
TppzNooCxeoFFVPfuiuDmdRB9eKnLwkCqNHOAs0NTpS3OlEyuA3wVSFhJoVbO59S
v65N1DSWbXlBT569XfcLVu3BHnfqIO+STsiofHoO3szPJQ60ShwcXBcW+xYuvB8s
gpl6ZV4MkM3iM+rEoXQ53Lj0Itf9hCtIewBValHN3um560VRg+ckL/xn2Lzp7wyu
p9Sat0PQj+0VtucqW1dgL+jG+phD2t+mZ1wS1p38gQw79Z/LN9WuV6ZYr43GJC4I
OoPtdWSwRt95dGzKL8LwPH/BquHrRRm0WHEUy/P70DSvoMVQ+Q1QLdhImUEpHJQM
bw0b2qDDSM/dpX6pSlLS7zx1nN/1I4x/y97R44fp7OEHlouEGCTYEYFeK/B1SjLM
T8ne9IMZSKIoavP/T8iG0sLv/++h0Gv6Vb2/Ze7k3aZGOtZXBEkFtWEawraWLldI
XviGj42XEEk7F0gJyM58E5Duxo2EUoJADDn9YeMVR5kmnnb8WkBaGtjYf1N2v7ur
IrxjFuQKq5RosSYTw2sRy+/xYMxk9iSyofsAc90Xex0i9Qtp1I0ak4mUnCPdilKI
/e4jM1Z+imIaBCDXtAFd3FYuOmwd1NRQVsNQM1VsiHu1stPuAuvKS/mcFeUJs7/1
IyKN4SEnLhkOikaklxy+8G8EHplq0m/tAwqxQkgD1nRmVLBOBkhqmGEmzX1ACswd
RBTAgemgGMlFJ3dDbKNcb9wM7ngMs8jJXcgDMu+t6lNos5fLnzkOIgI6SitIqiO7
KuGXBXaPoIbg15ic4OaZmdKDxEEzfsxut7AzP591xIDSxZiMyIC3eU472WS9Lbs1
2lcob2tMhiCeUH0/dbRuJ6vLV9hg2K/YeiK21kTKdclYGigKsC8AA4L8Ty+g88m/
SLB3CIX0tTvL8/Nuw1FHwYKiuBMo4HoOOmFeIGPLFTLEHtun/L6EkhelYB/3cYKn
c/W+oTuu55R+G2/Se7lzYSLZao39QL+w2/nLKOx6WHncsYCrcoILJo/PcUqqBse1
3iaVVNjHFgkNA9saUx9OccUZloULcSvTjMeKCtQu7VLxs7AI3NTsblnEjP41oZnk
+NzFEyfxWoDz0rZIkaVhoFfAJu2i6OuLZkZJyG3si50VkZDuDXPvdXzifnjrkiRo
yH9Idr5m3wLoaasVlDw+Ve+WkbvQxg/ne9Hi/xl9CL1NTVK7/KGVq/DMYEyumiTm
2yVaGP3HWXs6HUyXlT0tnpAGfgQqzgiuE01+FPDYjP6JDl/py3pQTCG4QF8guuby
hzjikd4+VOkChVBLj9pdDryeJe8kUWesptUiqL/YMcIw9rdCLASY3kIgF09g6ePh
qKLCl1SSKaJdgT+DVUN4NffyIu4x2Sxi9r80uiEQdzUxaM++BBAKBKpYQnx94bVD
OEMn5Y0iNwavDncmNUFXuZu24bBK0qYJSdelKYMm6rMgu57iHohga+1NhDLcxXK7
ESxpR9QTao7uiHT96F2iHG+Jzn8thFpHx9EXYF8FmH1XwQ7cUndV75dFa0dPiZ/B
VB430vSmcphvXDStdXotvYKSwWJBLZv6XPLeoq/gAstT34erBUMHk2Vfuo2PwZkT
5891PRCUyZM1pWCqAFhrswJp2Pcoz367c7UNBl6esylgq6V6sBgnH+g+jpHdOlSu
Mo119usaaKC+dCtxyz3j9HaJefMazNbm0OHcarW2vazEkfEn6rFTNPGy8AAHck6Q
esVa8t8mkJ+NMq/kQfv6ohZcUtEQWDPUUi0mgy06wz4P4c+dJ1eq6UurqK7KWCwb
Gy41eCH5Z/O4CmeJnylezv10uzStClX1NxhwL0f8MIlmOg2WlufOtW8zVkLRJrFn
I3EDhldLTAwBdHR+DR+k1E5CgScft9RPOebHWB/O46HWldjpFGCyF+uQeCSKPEHn
oWpSFmkz2wxWMfJOi5voBDs05kohVGl7JE/f2kRM2X9i4FZeI7NC7TgrD+KuddJg
hLIOk4nVmjSaTQ84RHOEJyMBP1ln7koO8ODBIU5YZako1mQ93aGzV/OzRax6CvS0
GBSUQTwfQbYZcXGt4pq/MWnvCGwKqrmIi51+p3UN97I33y76sV+dTmlglxW8n3+8
TxQtzqZeemFFNA/TfpOL8G9dP+mohC5jrWytOhUeUddgB08YfL4BVVu73UDd8Tq8
px2GlxG7mcn56dWmMMOlvUHQsxq3uUQRGxS9GUjaQFF2cMje1glEDFJoKrspbOyg
Nb0DfiQiTJEMWfAOM0p3shQ31NgZLgMfrO8G3Z5aGrmWzdMi4gjEj3i1vQ/4G/cr
nyjYbVyvsGjMBxg/Ox4r6p252eGiaqM53a76U07KXjMERPtpLKd9RXiguLws/IGG
eVZgYCv8gxSodl/4AeRznjqtW3y/keQt36yUAc5Cr4x2Gg0DONbgf+3sV6amqEH4
XxGJLkypii63X8PB9EZ8KmjzoibqQYu5uu+AwVQ3ld17WoZzFt/sR+XmqM+lb3So
b+5VPxyi+1yDulib07Z8CVWYnM86SL6EpqNn4RwE8F/epEL4zBmWlGVlrPDT5BhU
widZzgCDwca6V9xR6SQ1zw/N0bV8sNFGC0RRZpQm26H0CLZMzDHJ9ly2XKpqjkvb
iyl7IuDrIulVAY54AWLaHvSOADDoCsJgOxFC5zYiQQR7QUEEkx5FHIfrZtRko2nC
F6AtGiAU822BZZ54fd2vmZs05QnMJsJ98yw54WVJ76vN2jeWzSzRxXUwSnnXD6lh
WoUhMQz5DE5dZf2/QO6dkchLjYbwxXmpW/6NLJAHy7rQIo5h6RCeoNx2SDcj0TOw
NxkLEOLk9BIuIFifnCZEDnlylhfmazw5tTzIFHJGIdsAT13+Wtjj8UQW+FM7JeaM
cuHJQQkmoORLrkF7reYRU2VkmaN3nO//a52Q2/OnHyvBKVugV+jV6Y+deqtnLpMu
KGbZlMP6FKgbkmJNO3pfRqemVRHte3VLZC8PE6Y4210IoR4IKbnWh+arHlzBBbcw
liNyF6oTVbzgW2GDZR2M4VLszyh6dlJC8G8W8qM/q4gnnZ7xTgkdwkjBktmYelFV
+tN+EYwnrsH1SOIkdmLbALj8WoSVIwSkIcYLA4VmwVj6FwPQkBpdQKy3p9B1VBFh
np9WLNelKrPhe84VHxG5wlhYW2Lf9hWzz7jeliB0yUq9QEtshW9aRXHIWTZvZuBs
GlpOEc7LAH/rXRk2hTOQES0YNspnGcys07rq2zMTntw/xIF0gWZu26R1DhegaZxW
YSetBJQl0gTNbSxr0Imjj5PQtF/NvSl1rY4IuEo+noJ3uHUNjhhIgML+kqSI9OpX
y9yNhj/xBB4K2m92zloUaUbr7EirxqfaXlNc7WV+kP8k4ZXhso5MXMC3TuBueS28
q2T4l9YPVPhys4UhkDhgP0ka9UHGqM2oy7fdEW3wX2WfK8RNarThVO5pwN1uvKQ7
ErpHrQmk99/UdKIVvzD3at8H70VgoQI4mzM/FvolvZ7HSX9y8qUx3zkVyQL/Brgg
vxO0cu/MYFlDbeDabrT3BNm20Z5SkfF+28p3xoiEPh3adzr0RaFvQZ1JZ7ledbQb
eEiFpsXi+nayjt43VtwJZ9P7bvQdvwgV0amKg+m27P3noZkSFAw5gdRhlSIO2zcZ
+xxcSf/PP5DlUJiVmg3oaMXtsilcc5JqGW1QhA9KJLrWZiAxo7WW1VzGqop14C+v
72awIksStIy/4HWoTUKm75izWxSE+HsoDDXeSq0T3YSqQRD/Rw+pKrSj3YlKVntD
RtuYvJnodRjHNHJ1IPUr8MRTyuzjdUICpVtzo5vjzeJO+tW6lWSz41gwvk7hQuGQ
60eSEwaMJa5A+l3OrsxVb9elLKonKpoE76yb6M9ga7zOgcRVpSt2wcmNar1K3bAo
ZLZnuHuEqzTbGw7QoOTXWeCRVhVP1Wbud/qKGeUhY+HMvrGlFOvOAyooFgSfkV+8
oIi4Sx5kdVZl8Sc7WT3BVw0zWCLo9LHTy7JVcZxNcxOqC7pi7brQijIbKpg/Vuwd
TecAbdnCwbTAw+oP9x9j8Nt1S45zrfmxOOLYgOZFDld0wFekQg6ujVOPuMQNIl3Q
LC/Ni62v9rP9/qmleAIptm07xg388oZaZH9zcBRhvMKZRQUhGXcsW65qrbQiQdq5
VJX2/7R+zV9LM06FB5O95GaOaWi29yNlXYVQ7jHnFDtaq5jqPgyPAAokKJMTT9cL
9F8FypNWpFu86DABGccBSjoKY4bh6H9RxRMnVEpolisG4Kw2cgQsh05Flxq+qvAf
sb/e1o2v16bWvdPqjXT6CNl0dGJVro0qVBayhpGPnk1vG5YHiIszUZ99K3tiZ5+S
7dIvy6dGchE32NFz5uM9uzE653e0EbDn2vA8hRe9PPt14gs0pS/EQ0uZr3l7vanp
iYD9+lBc6b+kfmDBQBOHiCWBsvY9O5jWVrW/e7lzCX5L/+il0Uh8Gw75xWsTDaSP
1FkrtJshNgi0ZqlvSDbmyPtfJxPg1sbhTD1IPKKEBJ4VAO6pe9gohIYO93PECWMU
9JE6tetHEnq40mbaSJK23XiHO5enEetnjxkmmnw1GQoqlfN/zXTFs0MiY0ONLGL5
X9BCJBAfFmSXktEKpSqJL328QcYNVVQ0fq6K8uOEBwTFrErrUREaUytsOI8RLT0B
0lE3nb5FVWtWvZKlNeoqw+Ww0Qq/BU1eAkqGkjpqYrFgLiLxvGAxBQAF8EurlIGr
DIm9LtSTWPCGpDPlMzhwPgSpK+drEIALghq413mszGhQr1mvZcgbl26lxzAJm39B
Tl+0Itsl7Eb0StWtxBA1vTmdZdRTt5LOX5WIwMAk11uA34mxRAyoeCIF3Fq0LPQA
TN85yWrysCd08Rt44pu63N2KMxFoRYR10N6uSh2Suf/ogWvMTWr7cFL0xyVth/lY
q4DlyNtl9VzJebSprdB0iC1trhJvkCb0/jWRW95oOyDvUVj5ZegQSuEaK+4kmRXL
5y7qf3q+w18MyTFelYmXPlThO52YesOIPo4ZJu/yzdNYC/aubwFgXMqSghFVQfFO
WL3A2R1HAuMLsy3XNS4A51CRZ7FNjELadjS5pvxvmKkmrnMKbUYouhXbTDbwhrPH
7kZFGLliAJZNIgEssw7hcgMVNRDBaaiJrLqOlXfDTMjImpevezzMcYMD5cyp2+cL
9JhQphuuuR50xXLiueCewEwFKo5k5JUYEfltkIyLGTJnWAz9HOcXzwsWlkduQH1H
8/BMVZcZu+ZfA5DKBVadFXUYO9B8eUfDcdyiAtlcqrmO6AKnXCstLcjp2CXxsR4j
YpJhcr/A9J+jlNNLWrnKeSODTEHTADvzD671Buv2nAX0OvOJFYsgKDCyJcOxZuI1
WDnVWwzqaTqNlBdjNvsjkD44sz+uD8Y44Yn0r76k95/bFhOG5kOGuFsxAA+R6A0m
ZE98+jh22/6b38RNBQS+ts//o9NPiZChNWsqoXsB0+qVR3saoWfr3rgpGg9Z04aW
8ajglV5bH8hjkaE3HgOhpuIhIrwYZt/GBAxYzKlxJwQ9y/jWZt+S90WB9MF9njqK
6QnzRfxbgFg1A/wodYcMBDDR2LtTp2veVARJ/uaVGtY8xdxmb3T4tN7Jr2t2YPV6
ppttuAft/qjDbBhhgQ7ZGvGCJ0zeCtETVtgAW/iRfx4IRhadw6LxUpJXXfK2LrH2
CnaDgIGxUn2KcqdbcLr0IYxudoxBbrgKU7B/QC4ZOTHS3EsRekJEREyUUEEgWucj
B9qAontGwOozM2j2E/xgCwoEjXQ3iv2eu82JnCbw6Y4PczoP3MEkpYF6zdHVZ6bs
bAKr/cjbcbOt0sHWM67VesqRhQRJJCDjFhAwqiRUYlICRL4LW++OkOxqGMnsPmLw
zTXdeeZ9rhpKMEfM/qr/GqIHjBK5pZpewpXetlldy67Tfaown2dkNc9U/HSiG7Uk
r7tROTAHJ3n3D0jFn6cH1W1kdFHrz4NnSvck3xMIQERlC73iWQ/FeMynSMeGPV/a
mxb1e1b+9xEdtlbsdjk+Uq3JcMNFQeC866I1pNcP3cjDvEykgZBDB6qp4XU1p7jj
E2CX0QdeuSlsFI5riHeEcnOwMyiEJYDhyv49FhpUYOCbHCF42wfL8/zU5MzEUajG
zcdp0BMvXEoTXcU38o8KrW64MEDRbnudk8/y2wdUEFFPNLLAvVPytj60x2mwKS1N
r9KrSGffEciyIehVxqrionTjtXdkP27dJfM1cGSQ9cP/VFH204XDOS6DN8h5bLGS
+biQlqomWXP33ew1sJESsIL+b5ceHKEMhHzJlyTPtEZPW9mreMWMnvYPVdckRMue
AEcf0YmNHv8aBD2Bfn2GnzF9pYwT+KhsfRq2NChITkz/c3bJr8swDtE7jW51w0YF
S27pQgZlPu65sPz7iXuQCNIprr1CqXF1LzJjrbcBPU738lZuP8AYRIQwZhp3sCtQ
HTX+8ik73sMBEZRVWbm486Jvlj4uJU7/4f97Xz8YHd1kYcqD2elKpkGQ6XkovSWy
HoIdW7Q/gYv1WQd98FTDUHsZw+raUu23urKvE2SSRg4gvhxAo789sze0Ht3g0gYz
pycFzXb/jJF8P9z3UkPaDf/rAcDcE5iUTixS8YcXfOgsrui40YeE1wdTTtIX7Bwf
3Pl4XdvZI0fIFBfPeClYcoOkjpDNTg33V+eGbaOV52i/IRqyBW4823NIVEijW9jG
chkhNlCIll0DCX0brVpeqLfZ4oj2C4r7LiIilPVkEbZ2rXlSyJXEPOn0ASljtKjl
KXWN8OUXG5bXMewhy4YPYDtOIVxUHfX5Ite6/LAXO7yYaiOoooco/+xpmWOPRNbm
/dkKV/u0x+5pKg877Y2qCClZClZ9qkGIv8vHWIVGgYPFC7R9p0b99CVOP6eI4Kqy
oC8cU8xkpJ/nrHFXzzkzbJfLLw75ayBYkId70zhrAC6ubl942gmqQ9l/ZZDxBupj
tT6Zq8qqvRAyH2z7ifDdwgcVNuyRJAO8jcI6RG3zZ7mosvWj02JgBdBvVSfbU8vQ
tLS4VG6Qz/ec2tOSHlfk8k31QescZ4C++xHM9i5Wy3P2HMyIqr0x6gPrUjw1RQ1M
+nnjrteooK2wB0DMGYleFgboOJx+c7oELAn3fMjlk1PWvYdopq8QWe+Yo0ylgcru
ogn8R6I/l8hzLNGClrA3ZPV9b7zPUT9vPZWpfeLp2HTrCcKBpYPBxIX5w3yDJyCd
+K+oyObF1l548IQ2D+WhNz1i/p6hSHVn6fZb6Vs21+buHZr5a8k3knaILd92z+Ej
/tIt+4Mw1EqRlVLwXCBT05xKydUv3xaSvggFmSWyu3fqlT+U2fG4eXtMZmML2kJ/
/0zDlXSIf+3avA7dI6GWYQdQaOu7NdVhBaV2leCDCc9+aXVJn3OhtFx11mW/jW4r
eig47O7dQJtth91eJ7j7ZwlPh/B+WRbXm29KiSVdevKGE05Zs3ZbTJcdvn4ER8Uy
gKZUA1VDza/wuq4foeVxp72cApcZxHLtfslThyGr6kuW0hCF4vdzzJ0PciO2jJHN
IP/dvqnHzEYkjPHTZ4Xmifp8yIxBxh7O4L0XEVRD54tPFiXXde24cr25H3/ZCf5P
9Y4dbiweYZakS/4IHXBe7xjFZ6IlL5Wj9/RJ/3UDf9oJPW/ScDZ/3i7edkzMX4q/
KyA/MgwZg+khI78hH53xeXCOFELXgcFoQkAf7ohm0OGQkU4lHZc3c3NOlcK5o4bH
znRCTf73bifppzGLWH9ObXKLtrXpEfpi8NSeKQtXkrbYZan/1aMnRcSJyBMw9dc6
1o6Os6wiw11I//TRaXSMTJNd+DtPf84lfDepOq9eJK1DSoniBg9/loC5dSf7CkeR
8uQgst9WHJO+DUrKyu2A0aiTf+IYX+H/34jkvHmGbnSNOjuhfk9FUld0qbg7uft+
zrJOV+3g6bPDZHDk4ZlwZjCQN4J3xX8PCFZhwQhea5Bi+IKfJUpX+v+jeqs8f3rP
Ssj0NcF+nZxF4fp9YX7eZBpjOYDvR1LPpKZ+ALw7nporjEGHWHMEyPx2u//5FPR1
4n38rLB8Jr14sTFAC90gZa8I11DeU+ndhNbEFy+Gn2g4KkcauWVqBrhMEP0G1TMX
zjKEm4BgX0xWN1dfcNpMJJutNjvdD8AZvaRak8ZEOPQQeHwkEmgmYZUI5VtWMheS
Xb97mZC9/vFPL5yEZbqPvLbpXsWa28tfvgxyAZCvThLNtrMpDn4PSNiGsfSR5tFp
ZgZQ9t8lIdojH0PHgSNx315+W7yfWeLgA5UY7xlNMWYzQKNwLSi7dTYLH67tveVe
L9qLBCLA31hCX++5mwae85d953rdSMiAXbaq8pFzrzMlG1Y8q2t5n3zdrXkuK6j8
3utKoN0USphme4S1znFtIt+tTsHXHXIcdHvgbgzxElUeqavfSmrxVXcjsJ2br1UO
ylBec6KVhZHi9roZn9283u4YvOogJWptE9PHBSLGx2DU5HxFUwRW0L5wG8H0HJrN
ixh0DjezzmYx7kCVbee2D/V5jkGXvhIMoHPj4GM4VT5jpWkeDIj5jMErWeVmvmL2
n2d/AhUaUqEi3EFnVZySl+Fb27unHkdpwhFK6dSULV+PCF6Us9PpZ2I7V0MmlpG2
ctUAu6k0SYqb0zzWHUpxcxXy+Z+c+RYD4CL0OqBUMrjORYfQiec3Qx/DNmrSZUoy
0Szn4Srhq9xO9HKUL0C69wONfuYH/+vUNvUwGQF07b8eFeEtgcr5dc2tROR6BKjK
ll++lzWcEdSJosmpOPppNc7BKmyWIIR0ChCleg+VwUTMeM8z5zcB/gz5GhIVm6Dk
+TgjXNnGJPG30KlfMHn37BTSXvsMUd4uasPxoO/s/VYcxregiO21+VcoPElpH+cG
O/ig4qbAXhhdIwJCUdx6HY9NA06UicTdscU4XKzvJ/+AEZgdFCa6kpXokiEpWHYB
VOSjQb7jA7U4J89F2VYmX4vdl5JFQ7uEZnkko21ftycHKR5qBKI76H76iYe9UJeC
xhRhirorytLE6DSgne8tqY4rJLBVSGgxXAK5wcSc0PL8/O/MqsUuxl4uN+kgVr+O
9NaEySFcL0UsiwuFalTbP1D1Hwc4bBUMhbjgdzDSGSlXsBXyLo1EcrXcRw6HHmkv
tGIuoN050ClxfRjeyBZXR7/psQUs4lgw16RuFg9edsRnDqMo5rhrbkIzwVsSkWu0
CrCCNAQOGHGmqdKa7PbnF9PNtMhiuB9pIzUpbpuzpEAKNvGEvWkhetpCZ67gaojd
wO7r+5eymv8bYC/tmvxXRAt6ihEHBp5og1AS7b2TxZLPpmba4Htg47fuwLHFyPI0
EQupkiAAAAUP8zDRf4ojwU0HEHGOVJq6THhNGNkxEEhHPTOO563ZUHaVo/bShCof
Ga4WsxxC9Zj+A3scPGELn/iwhRrc7D0MwkV5B1E666HpV8mrWqeQiYedjiyfDi+Z
CTbIcXbpxz5CWNu5xijUv2gjTwmKeHgIOleJZZSj88mozTOwRw9VQsma97C3mI39
bnBbCkZSDFEoZy+4ZYOtLncNVP4rVBF4LSsb8OdwnnWaQ7xJOg9KSP2uZ7E7tEkZ
B5Ux9LipxkHJ6ZI8RDRtyw3ShKkmsHj1nAS3QyxnTlIVGdH6lX+NIrhufWc9owEY
hE6HIA7rAn2zmAGGP+v86hD/oYMsfmqAd7CUbVnftmQhmjW2sHwGg0yhsdbg+rZ1
rcflat5tagRB51pQlPkh11PdUMSWPKGn5+0q5M7Tm3TxBtwqNKnnh5Y4JF7HCYNS
sRzjViiRhfAnL8Hez2aA7QOXn011NI0ThSiIDV2gqMM3HfFMyX4P7t5ydleYbTgQ
1SCYOwq+0Sz8CLvIBKHU68ce67Qvv3KKO4swsEfEWiuYmrtxI2V+6Jq9JAcA3/CI
ogup7vvXdaAJfPC9+H/f2BcaVyJO5udW5bVEGcF1pmgQVCrjDjh+7iZtULkGQZR2
zRq07WbleGWtQbVlsld8P6TeqNo8sSwroga3VoQW3M3sHWzD3cTOkvfbGM+lHux5
ubnG73xJLtWnxy8NLqyeM61HqdqkkN3k2VVZimQus6ykB8fef9Mc3aY6YdSNYmpI
T+vEJeWdS6v6Z++zXAa30HGhMnDnm628marBsworW+l8LOF/IysawG0e07ELmIjG
Wdx/Xg5UXwHFWJ3AGtrAt2/XJNt20FlgvbOv75byRckgpFvnuAt3akyWaH9LL/A1
ZLjvjcAfoHLGddKJe+fFr1bDu9LAy1S2ay/9vaThfin2HtPvbOd3+yWyqKClrRjX
9I95lWsEs/B3Vlj7neSlRQVhKCGM3+a86sgdxk8b4+q0ZzXzgd7TE6pw1oCxIwrR
L5350FLDLWTkEnI64sp1ZO72Bkd5rm3YA3VORNY+fJebHTfI55CJkHB1lXZB8OBb
XzESC4/gO9cUONAF/0r5Wfmow5qMohV6QXOisZtngtPNCTp1fJV0piJ6hkjhZnnN
gVh2gm3A9iR/1ki6KedUwW3dBxpybycWal85htlEkHVGREoK1CzkbfXT7w6+9/lT
C3Z+n4G/Ne26/CcVlVx7ZNMHDjZZaxSiUK8qImjLW6HFM9yxmhb4wFJwPomMqoHy
xvmgSgPWhLDxU0gCAKT4tj1+80kZN01rVf/fbs3k70HcbRtHwuVUpV6FT0jSd4GR
MiNKd4rx7Qj4cLz4eaYS0o0D77GQb57b9W1rMfbf6JO3E2bg/c6bHvF9ePzozyxf
4BiZClxDiTq1DVJNFEpx1GC83kVN6l77KVP87EcW0GbkBypIN8O9wdNORhiWKqhF
rSuiKCa3qoHH2aOA3LvM90bf9OaxqzWXaYb4hz1PaTNWyahB6ChShsFiEGtsXDyz
jADMat2jISmGbFS6AqC+7rwiHgL7vOGogVEY5UWiHSCN0fUkwcwjxHRPzUb9+s/h
Rull3HZQhtVcEuvOYu8EgzXjZgU2QPTCdmlDzGsiZLl4kYEkIeAg/sYdhGXYiMHS
1W27Ba6M/UgSq7Hh4GdN1mrjwn6+ezI/7KugSHvq2Qbfl1MK6GBcFo0Ve0vhL4bN
Lt5YKbcOcqOxya0Ke8kBpBwFJYUfGuVsOhEQSG+iG0VURfYkAHqSRMx+Md80JbYL
3Vhzfgp4eYoh1IWeirogmtjYnt4E11xEMJT7DwKvWWQCdDWNJbOH84wGRBa0BM74
p8LtKZ/IlOgmgkeESSVrf4e4DQEbiDF5/zmlcdoL+WFhPkuSET7iKtcP5rnbXr6A
nro+BKKQj8LecyJp6r5tGSAIQoKVMc1MUE0hAqtnXGtasZ0fRQ/6OD/3065BJLFx
nEwmjvnpNGlKB0arsTougVUeFnFJMDTmU5yt090seWg3zgAWkNbpg8HmAcubRTmS
OuacUV0fM8Ikfk9dTqi5LB4Is1csCIcTPbXU4SHoEC1IqZgSqiooldEvYKMEqUK9
l3PscjO3lRuJd4hdzr0OTtac2GTfyKSVamkateUITtpVtU0FnksSystBH61SIUw1
bofp4TiZ9DljznsDGgr25pUp4nqoLvdzK8/bYLJ0oILNvBWyirIGdpjTDSCR0cW6
7fupgzp8Aifcp8WMdLwYxHsGa1NS2zQoTmQcUcgovPeIw4qr3f/pT437n1OHrX2+
T8xSDGZzfW7LUTFdJjYesHqvb84Qln0gsQVbVWw1XzRPxrdPb7kZl8+GbQG5IenT
bwP9pjf8lIKsio5W4rcJtWMwXQZ+qFoqTPgs0erv42+xxO4S4hNK7j2qZnB90r7e
AOr9lY4/XL8XRE0VSCNtpU69IKeXhPm10fkpYyhbKhRFGHXuxTmW4Ce3iMcUPa9t
Ym05dkCYsL/sUfBuCdUb1qj1UTVSmI9ZGhWCmFjsM/D23BuAZYmvY9D2aARx6Uv5
6cysLNnHjDkn+xdNe18JVpqfN8n7zgEH4pSleOeaO6qaIZWSSaNwrBfK3zeTE0pX
DT69wxxVK9CHL414p2NvKvZkyOSepzELNAbPTUWOd+tpaDKNgCNQwWXz7LtsEZMi
63fY1UMYCUUQHjD9sw8tR4p76mZaeMqXRcF6KI6U0zdwfpNBbEzuBy0SOKR7npvJ
A7OTI6BIga09mQ2ezriTxFBK0KGk8O5i8knak+bh7/f8niJdm1qvVh8GM1A9XkFT
/yKPmNz/R9B1W93gHEjwUP2Q+G0h9+qUeimA1rTyzBq+0Q0ltfUdvx4BFt7nIYqC
jnG7pirUJxQlgUzLIIm5EjpdD4QjLCkuCNd0+3gdj38ITuYLrt1Bkm30GR+Qjokj
VsWSIHunMe55KB1DCBsvsYr6+i1OMQyVwENAeZY0pdUd9Em6OZlVtwMadKixEcGB
AtZKlP793tvYNcYdHdaDXT2jEMiaK0zVjT7Hh0jx+vlqRdGOM49xby1pSIPbdv84
SkvdA5iAmc41hRlH71F34IlJspqUauY1gmopnxu9fyMFERq4GsB7Zjfn2UI7lxWg
PdJHBJJXuIFx6t12zcFvxWBRJBYCgybkc6Depoowjh5+DV8tV1aLfq7wQG21I2Mz
zL2oFR0kn5MAXlMebSE0O0t1s89KdpK1snRny4DhP+qzSpIQQ1lWlObNfdRbfxLs
7ns7tfFSPsSsVmdn4lQiqSivkgL03eSxGNZotEczj3sDqcJ3MYkvJMfb1lbaNisB
UGzk0EuhneeGjReB69AeupYH+dmbSDIHaISX5D+BoCb0dJcFIctZpTeWxlx0TwEJ
xhHWRzsLWwa6MIvws9DaqVgzJfYhHYyamfWtNEzvA0g0Y8q50Gp9c/Vzhb9ssMl+
Nw3LlRKDThWVR6EwETh4D7IZ0db20ba6P62nk/5qRmBHkIQ1apS3j/oax/CWUo6B
pSfx/xh/SvLMuBOIXrOpyS3z25fSUJAhrtUCe5Z3PI7ydarfK9Lg+pEZx1J5EgNq
JlXcQd4K2hPXMudr9Angzxqggqc4HTWj72uh2/LY0NVfhvNKc6h93SQ1Y12g0/Ro
AmJ70lZg95Qy0/aXXaXAFkYXkMvtBxWGje7bUbAikbbIugDWAHr9uVpR6za5jRdo
zrykqBzHGriSEQRJLUE3V48r3UR2ljfGE4x7A2xp/WhO87dePA8oMoaKYFCm6N+i
ed8L/5+AWN6TCzk0nmlBMXixDhzQT0/yXqXqQItPjqP6MEUWxRmX91srbfyXViVE
TDKF7Qmh1GYElpH/YObl7uBl+VvfqTTgdoWlGCvPerSFgKtZISFfuayGrVp6Bdod
nq0fLl9hStkdWyjKpbzsSdwIMZJfP8V67rBeSpzct1HW4EQhrK/AaoflKUqZx7Uy
0z+0KfaEPKYnVPhdX2YiFB1V7oEszNKE2yXGsg8ch3XpWhiIBfw6QZ11OlR6J2vl
+9ttogkgRcjK2cCDv15fNRHPTvUdOKyuHUpGP8DOz8HIdIDlSFadtUOcit1uT4Mw
62zmEGfCbQgcQL0mGTa2cylrw4ITxdQIj5Gw0I0LQUTLrB4n6/HGZk8+1U6QUkzM
d+0Sn/1Jo+ySxm2i24OYGlQM7203K8CpdpB1Sb/JoMLjz7ao0jZ5pUB1v7h0N0Kp
SiOr5BTff1gEA3o7Gj9ShbtcaGCPRuE4DbHs/EgMYj12dVT9jPqey+eEYuxwkGvR
Q1j+vihEfCI8Ys/2A0Xium+gGe6GpxXqhmXLGd+08a9R9J8ey1uFwLTdaI652b+E
NuvnQtgeE5IMc9lFZOoFhsgrQ3VXzj1lSaGzdJb4t63czC8inj0SGs0mckE4TjA3
Ix9i1R7+4a2nG2MWYZSeQ5N/lsYojROehQiqi3EBSbrS59oPPy+WMP3TyCrrTq4P
KEdBImTf7jR0XCRoYoAPTfjj9LNaRtQgCM6OCWifQM4iRZXKrAaeXJE55JQ44qRe
hlIEnv0i2eWbR/VgQ5PsXv6ph/WUwNQpDAEpMVtaIa2AP8KYl1OxqMLiWtBRQTVc
a2yQ0WZ1gotLAFZ+rCoGbUT/I0g6cPljOia5rnwCpiXZr5m4Q6MH1EaxU0Vwd5Gt
mV0DjfQX1W2MmJzixQOXBM+LzwFcVnUSnaoV51t5BTuw/4+tGaviK4xnKGoW30gk
WfO4ot4LQc2qQb40vNDGBPss55Jt+Lz4e/qvCKq+paXoxBV3QWQEMT0To1RhFRK/
lLq8Qp3gSta6FIImCzdCMvVvMAIYmpXpwc7uA4tuQpY9P/wIia+Sv2Fb71xknLyp
N6Ng485cWEjAjPcXeuCobGANdOXpbOyPWrdAJ+gmAzoyhcc2p/bfiT5CRMwsJm9n
mZIKHDeM/gK7K40bx83NIb41q99jWcvJfwyVgpYg+f15d1RTdWDuuoMOon60F7xn
L/x8GPhiv3eutZYeCtR7i7MBab4L7mxS/mzwE6qtvuUo6m1KRE17zAp/mJUgZ2OC
SfhUo5mU1uJEl+RCOJ+nlJUWEP2p1w34zW92EB8VVJvpxWrIZ7d5SoPv+1A1/4bn
NqxTYBwi5CI8SWItwRPlYlyXolEXDo0pae3OJKwVeZNecSE2uegwu1u+kDuYRxFf
RHeEqvL7VdiO3by5zaWG8gw6MylR7BM75Y+i+XcTI2Iw2JIi/ChqI7UzJ/lyUM1m
IvxMMjemZS6Lm+xfRO+6KWm0SZ71vaYU4LyLzag8lOxDHrcT0t8lRPHGarTdD28o
EsOI00AWyPT1PXmYCEM9dQni0wUN7AK7jjbzIT6E1AbHbipp/jiwbPBThs3NoqDD
eV1o36yrqJHsI4sUi/KLvtvPfR1gC+krAXgm4eQNxfm3LSJ7U0j5Z2Qi7NODvr3A
r6rHGZCWZt6R15MjzEWr6F194KthssICO/Igkzp79bA9sfoWGK3zoKN9a/RAhhMM
rqQ/IMlfo2xBB8CsVH+I7UdShJNBufz81vAj8XA1vpRDzNH0osDz+rp3IRwLAMaU
oOjx0Vk6rAMYJZtSI0l7k0HN0MCxmuX3y0pjNp+xJm5CXMnOfx4tvKsFDZy5pB+D
RdJitFicZz8gkrjr1sjCQ/PL5lDk+rSh/SewCxoDxZZjlPlbeNE4VXn988nLgmpO
KKnaJ0y0QR551o14IR49sWwyFQ5nWfio9FEXzIPXVYN+COGKOwzGRBKnY4d1YVCK
Z7PaZyWh7DauhNCSZBUD88ZY0yS+6rz8vUYZWQcE+57c+MUJs1fU3pNhgIkmgDFx
AUTVLxu0Ius6xETZsEcvY2rVekJnaqE4Rw296pIc7cD/r7Pl6y/TRQ3DCxNJCkmg
LaTGQCDLpSPSTDFZDZWqdcrp4bN1+4NVhIKIi8VdhRDoGDuWyG/xxYAIsXsVP+jG
dnQxN2ItK66376YmX0GbUe49bRjYoguc1q0vFzzrzaOKJxlpGflkGd20UGMviw4x
Bav+62WyLCpNZYyZvYuu56LnRYuqRWdMWsQsNMxTkr3dQQXQzTKJNeKA+QdjBgTj
IF+8kayh+OcI2ZkTr5OXNPSJxp1CMhT9j2jnOCXZfIVw1M5w7KXocVcpxvy0ECuM
NXTSWp1mvq++EaybTCJFSEe/K8mhvLnULz+dy80erWjmhUJllTxtsIoizOp5Sdol
icbJ3Ja5EtY0FB8vUGzg2stUsIYkzPjyz+Su2a5O2cJaz6QmxBbLO4Yg2Lb071uE
JIc14jK6NzIxCrjX+Cue5yUCNrj4fr+9/hdjnei4GlZuQGMugUUeUbERlBxFdHVK
s3RQp9yO/c5m2qFo9a80wCkCEprStBAZiNj48k9Q98X5rDrIwQw+Isrgk8znkpF+
uoCa+5K/gqVaECzeMz8uj0SeNV5Rub8FsgDIeHx8xnwor9cYpXaO4wIl/cFb8PZe
NZENLUq/pZqPHnKIvuFiNxgZY99MJyRhr85qoCciFGwETW2iu45NQpyDrUwcBRGt
qzHNcz7A62m1osvzswIR2hxwx7a1Laf8UYLI5MxW8hOFZrShkUeLbGn3t1OHl945
cMsR7tAiynS8V6YLeUrwTkvco0XUmvfkhVyirysyyM8FiYC6aDRf/R+xpO6u46+t
kG+q9Gic6U20bYNztxv3HnwW8pY4gIfOWRd+gXKThg8tdXp78ZrRIzQEXyUlKF9p
gL/oaaHiK04cCxJnfBHgkcwDZ9+Hm9yLo5YXel9tsmrQTxxiXLGOx+XOJGiDrag+
YOpel4lJ6RstFNZh/LVhSZRklJpIXbzEWvz513IvHbJKyuIlOgmh7AkuzuodxonS
azJy2df61DflLHuYd0aOKjjb/SyxMY6AzOU7M4vODjkCfYvTxZlphCSbyi2QeXgj
FKiY+DNKYRFAemZ2GGwbQSRaTx6kSuBgHrHlx3XXv/Pl0FgTC89XEKaUzx/ccbSo
J/FiyMo/pYDQVRIidFTBxl+2jX079Nr3LDv5J/rzu06Gi8UHnXfc4kpG1yicH85f
uLQBaH9IuX+tYyUJjgDSuAvB1tkfj6cupS+RWU5gVEYtylemgLTKftcsxbjas2Q9
1M7M1ERTc12o0sFJhMJkipOdX6n2DdBoBUFianAs8X0LL8tEuotCAoNXFAsmxFrA
xa3neXmGdiDTN5KxGPWsDho3giEvy+Ot12C58uDlA6ZUnfKJB4WhEOtEXp9mp4Zf
QvUuktDlfVLULapAm1CAfAw3rS+2WjiQWTDyQYnAqSV+GVo7TuKp9eZ20T+C7Anb
Si6xAclEB+MVVfCS++fb4BCcXESzZzAFEM3+Ohzubb4ZEq9qzx1Ier+CTDZT4DNe
70kFbquwRBGw27kH2u9YZP/Wsa26UOlKbW9w9fSEENkbDog+Yy++jAGRfWP8e/7n
+E+BX8C+GWaXeQpApyBEuk9LpNRcfcsAPPu8YXwfoIVsSbY1raU8ZSnAYudvsLZj
sEic7MJCyCM6Vq+s+RFHED/TkxBsp9d6qwVLYGUDt/km5X1/LPIY1p0p1Dx7A5U5
q/sksfwlSSlcPRWCsu70RzspjNpqsvOJdeO2V7hdyH4yqypJi5YoNZPIMttbVI9V
kP9W4sxQrstRomjNEftyAKwIMlDnb2HrZkkLb9RI3Z1GaS/SwDJN5fCJJ8wroThD
Ob2W8pD3CQbGQlNBP3QynGp6Z+wd/2z86xRinMr+3xHXevve22Xkuam+7LaIsZgC
UoSiA+XY/EnFkXIXViz5Fm3PZLjabpObOjZ8q3rT29kNVtxDpmfiCvp7LhoMVz8o
gJXBZg/lE15FAMEqh8bt2d3m5sxAaKXPMDNmuOCFG6naaLZAwl5dE68pgKby1t1F
9ATi7+wN0HfpTwEBO10xt4dFlh3OiAiI8tTXLK50+MTuLzhXX/l4EtFaD+VE2fEk
UEecZ68Fc9++n/L+V+Ggqz8M6OOsLlO0vcH1RGFkH3oK6oHOJI3+m48w+NhCgH4A
FeYiBpFAW+Vhmud+VQtiYMEfoHByOyXrgT9opyUZVZN8awkIt/u6dK40mRY5A5pC
pfF9Aur97AkfKhXYlj9KfRF0LHsA+ey9eS+b1XBBQV/fLuEgVU9RH+yjitP6Wa7Y
5wANlFj0moGjIDjrHdd2zoLhIcxljdQU3a1My3QOguSq6VOcx2r2ECa1Q65wTle4
yM9ODjKV/OeVs61WJW1xkfRyP5afqoM1EZuEYm24s02Ig2o9Luz+p6ohxAikdszE
EyBo+IZ6a1J7giZjtdE5nutMaG1DK/8WmP6dMn6FzdlGm/sB8JDI4LdTHIntge4d
hpoWkFeoOFlxEoMi0nv98rQ7ty2diSyz+ZCZitsgyxgecop/2wjGM6mp00pDe14S
h6DHP+VQawDP5UU+YwRx02O0mTv0APOuaIPTQeFNmbfgcErvrUT6mGiF7gAy2VlG
CyT9looR0lJoYM7sogdDEACxFAnCjdvZsRPggnwR/JwL0A1QI8OWNSQOfzNsv0D9
jv+rXNZci434hoCJYa+VWpjM/WLyAlXiig4VFJVeU4Gwp0wK7iXLb8YT50H30IfX
9HM9TuIKZW4y5BwwKX1io/fDRv5FkyEn1Uh3tj6WqBcV1zxGEPegzoYY9SHTOgkl
hVBkyXkhzmulYVdPewF38njs7el8rvuZU4mcOBSocP5OfT1/2G3grfjDsIbCNSkz
o7ZTuwI1bKeEAt2vrSj7pxjL5/UGCYvoNO2EZxfeOi63FCsDfBgb8lW+5RlAc9qf
3bJG8j4lQ0un3wZ5fBFvBIQPhzKvbJ1lVTy8lcQJd2IhwD2QsjwUuThNMNtcBV08
/02SEtp9ybA04FEDWr5mTSrC1B/9E2rsMsyj452TSUiyKVSz57r1LYuTKB/idRNV
Q/5CNrz8Gew/7iMRUUzZEzq3/EInLOiL9C64H+D89Lm6rsRzABIZiqXpoDJXKVLa
48KR+QpPZqwrB2W1pKHkcXK2SGhG+60HSSyOqyHeTvsyi55MPtvTOdumNrgbhnN3
NNEd7d0dR+vHLe22DWyIwnh/PDfz/FsZaLJnJsk6odK3eRSxIa9z6mqal3dp+NUR
OXvEOO8N8EXb/wsABKvAuXDCQ8csPh9Ph+geufWeTTfiN9nLFiSMYtkEgt+2JGI2
toWrHP7qphXpL5s8rp560hbhp1Rb8jljPU5FCHZeezLTf9RjkBSXsG09wdxgyZrj
vp47fJI2VeaIwzauiJ7chxYLik9SLg/eoImnaZFpCYXg06CfxpppOUgW3mHuQyRq
5NDAkoZsq1A4t95fjz5PvXJSaOmi36yzXfs0ga+x0Tq0/6xTBhdJOUdJpr+GxjUx
FZiQO3WGyhbbc17hj5jpwjxjYwzYd0plD8zWhHkWOCzsZsTOpU1hTjHfgFvWAwJb
rarujTvq0iVv/TcpPFOblmO5dCHXXLgCVBbYwjg0ug6G3X9al1qvuHqh2b1UYiDf
eJHiP9faRtO18lk5I8qaOsGFByqEUvW1GcaaotSfcTiaXqSlZIIImUZP2Egf6X2g
0wGIOA+UKj7Q7BGFGNsEfoU+GGwHwdodJf/QP9yhxLe+yFKqwYG/A+iDvhNAEpyK
8C4BAcL7/XVTaiFkSn5/rWf869YbVERRVS3GdiGfWmgO/j7ftlAUQYIa0hI/DXun
5PNob7tI7Pyyi+iuq1Z89MTPjx1/24UYILi0Yo8nRDNVU8GYgn1KgFGnRja6Segk
VehTV4dPaLvTENoy80AWtYoidvkjCt8NUy2Pyz38Ltp1soHvPIwvzTrp2bnkwBn+
KVa5NjI8irxB/+zhfWzfbL0ag23hnRmupPgVdiFIdzhOBKXZ9JBpbOYBARK3gMzS
EBCw4VELkbFrOo3H4upxzhiMSZTwbjX17juIc8RoqVj8qwgP6NmXACHM9XEfqEuH
heH1twsj8PG9QR+Y0wpuIj+4nT99ipKrA8GaqvNJ+2nXa/b8ZOuXcqvtQG3xWFdz
jAsBf5vCozsig2NfpNCu97eaRHbDfpLmHFq6mrPvhYJFg+Z+XEDF9d4JK3iDbXnS
S7wQFPMATLBliq8mwGaJtJSTfhxyNJUntWAyD+toiowHOcses2NHMeVCnmhVwUku
pDPIUbj+ScxfPF9cVGwy/sVOsUm9XQUO6lWGgkkD+uYEOVEexqNt51WAz+hNgrGg
iRP+GoGXMF7STBxI5hIY9qhOHbt3ekU411r7UK46BqZGL7M6kpzVMGOtIKLGY2IJ
fqBmglEqWyt9muFUKvZk3J1Zq35Lrm6lUo/TOCIxrLYeE6LIR8W+2Nw+covJYxeM
S+5h6WOZDG6XLluHwKHeDvYi2aEPQHxXQzoBnwLF/CIcrCBUNDBVVPqigMDfwi+L
2csstBjurpTvkwdxQcoCMsT7RVJueXd7e2IbcHGPPBTMRPN+01VWd/z6tNnIWZU0
N043rbH9L2kmCugYagZSJ5gnV0OsPIZWXDvz5KcMiJtt0lwh3ESWGcMkqKq9f4RY
cj5QjeBAiTjs3+X70LGNSpmSshSq30mEuYWf27bLbwFT8DB3XB2Hf8XI1IAEUYUY
hDxhT8I1lMl8kJoIEnebp6wZ8ffY785ZPllKe/rcjvNMziGu3I02awzNU2cv4noR
upGpStniEwXwNj8/bF13JXvSo/r566sMSnf31RJ5SNvt0HI29gVG+BOQjnnYhO1d
qU5R89fao57iI0FvxrhNPetG3jHZ9VeAsBqVgPFGdGWQ4PYxKxCdsUsusleohhFU
NDmeLQJoCg6xS4nEMQbV26B/jAaMozcbUhM2REUXkFmR/HnsDEnGs3TXmzEBacLa
PyC3VTDrX5++lyCae2QH3/XsCHte9VbxclbqbucRERNUo0Qafjuxy3N05a8TSEhJ
nrMu653kdx8MtLZ4V5xqFR76I0z6Q9NR/jeOgB8I2pmblDNVoyfx5s5qgRPsd5nf
JF6WhDbaRAAV7NFuaB9aPvUDWjssXhI0UDzrU4FRjKUkG/MohZfYio6cHw3yQngg
kgCZyRqOAwvdFVRcyR3+bxzTmczN9moQQSJeB3oHsI2QC4oDVo165rzfPn4EbN7r
fu+D6ibNV7tX1+sryZqYZ0KT1ogJZYGe7mrtx++0CGhzjFMpydl1+XrvMmuh3MIP
v8Yw4Iyn/0cjoresY5aGXS86hUcTomcyWcZvv1dW+KfHQQW/Fxp/2RVZxCLxcQgF
j7TD0EBhbteFA7LUvYysRaBJCxBB/eu5/XPiWgfRwxr2MbgUZsSn0xgMoEBL20RJ
1VURk2AUQUWvmxFqLby38z7JKqWjmUxIYrJRZXDtsTCXQc3QcmXE8HGFkYvtCUDJ
xA4LDArj6q69AcyAilpE3XoEjC3BY6Iy+CmZnnIQUxgZ7WdRSUc07QIHIj+g3Tzk
vouk324F9MjYScST1dUVfECktpKJNMXO3zcdxF7SXr+Hx4Ni5Cibh4KmyQ64IFph
qQ99V8ynbRB8niSyhsvetexy4Vb8vBlntFN3ziXBP8I8GrQgX3Usm5eEEDixc06y
AjNoqjFCtAPuJXEDZ3eSp1MiDZOG/RnbGr5A8LmUJjiH2WJoJJulC/8qVTYvXMpa
6+x/vpfDs+TZJxssZSUG5SINzeniMCGhgFaEwe9gLVFjUfuz9krUCL6JTQV7fF8B
BeCSw3tg3m+9z+IUZgWerkZzDeRvb42KzGCtSDYPopQ7vNDgXEqoXH5ZX48yTsb9
wyQq+oGdPd4wPhkprvaoEBg5ZcS8gtCKcRa+C23fo6jdfCKXXhw41RYrQa5CU6Qn
hj4QFTW2CqFIe21slrd42Yos/X0nqIxOc1VBy9th0TBXMpiyKsjbh3fx3tooCk0f
O/UyrjLg15TMFfxGD2L12NnZvCLjL/LapYGnkX+HLGj5N8cIB8xu3f0plhSRbkL9
D/bRTnoc39y01QYFTv3JEyHg8owhIG83B5JwTJzMiiW365glVRpFWXu8Y2aoT/Qi
ClIUrbH6PLfQOAE6ZbkD1NuE6NUq3N+egICC93GUC67uo4Td1NbKzFmjP+OzRqnn
cew6CEuSzl/z5XDnuTcdBPgzS6MoiGchSjj3SeniQcvcjBKC0VfRs1kclTgJyE5f
9JiYCIEY1gJ7aKKnrSFeuZw97aR86cU63TyrMiWczNaHMB6WHMZaDWtYCoMvaIka
rkdSnbD64MPuXXvcS/9ZkukSKBtAHc/nFCQdWp91/XgsMUzPJoEausC6l3K/eUKK
2+ZnZzrYnNPQ2jK196G+hiu5do9cjTc6e7teOQacIP7N5vpX+clWQY7Yu4H4SWAL
2ngLIfewzPAd+vQZhgfQSF7H1Da8yfVBNuMqfAvzrEUEUTegC2hAt6WMqQrc1Q0+
1dADX2tzii3KMuhJ4cXBLYtq0gytTPT5lJD8CRYXoX00X9uNuOqUzv/NqV09Ni+B
Fc9OxUTFy5Cf7+m6yn8RgmgeORSHZ4EPrpDv5KUHTY8reMUBOKRW+LVgMLcXrpDd
VBUEmdZ/GfrBCNE0l16lvkDLFPefNUVSoftYJDeNafdAHG6bJ29NTm/HhMLa9UOF
jHRMaIRL0TqdyEDURL+y3B7PTuuDIlUYgQgM/kQ76cO2FD5dKiGk0dpgV0uT8Jvy
P7SkWDpx07+tWWp6XdWjLA+qIAU8jrA74KVrmt0/xqlCHt89SJ+RvttKJRByehii
vjd/IznON+WloF6pM9JlbibBJkrNWC1Kt+NI0kBdiQxuzQO3NuGiM3pFQh3rYiON
TnhCRwQFbn8iAOtG+j49fgO9H5qeCKgPyrZPNeOwQFy8ElMpKAoX93D9w6FUo7lG
bPDY9u2l+B5yWMmQOZn8Ea2dtms7lmVucYxf2loJqywDjeq7tIYuw4U4b/ZGaDcj
dAzSFLHHZD9nD0VhtWY7A/8p5GDpVIhzEdCfAHJc7t/gQERDN5yLXmQm/PWMRNN2
eHZ6C/pFRvWE7je24tyQdQM/R2WDKZ6V6dC2bHZ+57m80SNDSMHb7t317jmKtWJi
xsaaiNTmGdFhv+L6dgp876eSUZY9xKpywyTYfEnEy/8EKHJNqTjmiKcH0B74Zvo7
c15Ijh8/QMkqjByaS96aYz3/4D8MkfTSo2iLOXPGwzoDTNiVOccQZD84rRpmbEIH
yg6Q9UanYtfU6Vrj/x8NAlLL9BgV9NIB5weq/YZADccN3PVrdpi/Hib+D4pLJj/c
QO+v1CxCr2hIQ87n+VTencPzQPFSNdqtB7DrYy/df8L1Te+NzuPvjyxnL46w5YmE
w0Hc4znow87yy8Q0Y0bXeu0oNqMtAePaYXCUvfdvyh8fFDk2gc5hCeZbFrURmrdv
7R122b0nnXNkxSz/Par7dyhjTBtXDN8T1X7ezri5QI7SclxMaYhF/1ysjsmuZeXY
bmxzOXxO2nZp8C9fRu/Gfd7UZu41N/Tl0ZKAveTqlb3sCS7KexdGCNXKvIpsBt1H
H8grS8BxpCweVPxDB41gfG1h+a84Z2DpnolU2g7Loeic21grR7nkJ7sKU6emgJlR
iKRuLOkqNt3ARgwkdYAiA/negoTqp0fIWG4d3YdzNwr4rRXnnn38g6QEN8kc//vb
aDSanxvxbw5EtwhDZKuaz9hIphj3pLLZ5AJ69InznqT4j+L852uEe3DepsRSM4y7
0wQ9lQF4msXqcnrLBYA8o0Gl7U86ILmFlkkZNGeGlbXcf7e/EOD2d7Hhdx9BQk4x
AjFVGxRFVOlybxpYxod0C7PGF4NXTdsgdSDkJVm4XwUlK0Iaci+fRb8sTIv3Y45i
//LVvZpeXWZRvZ3CF+AvWwu/TnbW7UNrsMEo0y6/T6ueP88IrsVeUlM71zXareiN
/MnNNVsGjiej84cPqT+tl7L5sPCi07zzhBCj3FC0BeZWbWdGO7ANe/Q7b9v/pXNT
Hub630AJLXWEAPdtAhZnBNWnNiRYN7NS5nht5d0lAa2f+RDWU8TwWgisDVIqFm4G
3s/84HGhMiiR4a/j9NKtWH+JEwbqplYLoH6lAzan0/V4tvBZ57wrI1OGyh3IFCzT
HInY+lnBZxgRYf7seiNA3MwhgClNm67La0P89Asde/et7PKFMcLZ2q5yp12Hpp/k
FAMq3NgSEkEeroUxUKkS2XXzso9wCCqpgY2F/pgIa9gzVaKZ2Ku6IiMp+lI3KHKW
68u/lB8E446Avy+dfYbxl2Nud8yWdgUl8Qeosu7turpJmsuDtMQJ9mvSGqlPpftj
onvCho5fo/T6/Xx2k5D5CyQk1+SqLGCQQK1Zht4KzuWaklryyC5QLvIkzml8z8vV
oSjP9YnPJRB4iLt1+dQSQrbIrzFHc/oefTzmrKCLnnzfD+WTyjlYUCizjjEO/+bg
BP/AZmQieOZJbYCUPUNXIiNI2E7pR6k6SLO4ek/4mDe4TXU4f2nDKoB5PtuzKHUb
OIR0UiXZtp/4we/Rioc3wPAZDkfaNIxZ/VGIAp+NdKqNRZwu5XpRc/DdU1ZUa5xi
ECD91LZO/8Hlu6K9lrMlOlsJ+YXUDtdbo0iH41C4uETQGIAh0wlTWI3osxocqK9T
zICM1v2CDzWC75oNNIN4As4Yy2AOjAJQnnsPwhIqvLpbLr5CAP3iogBMWSU5jYwh
+tky8nN/dpHuMsSzNac70Kdr5etZFfVMnn/ZpEzWhyPiBmlJfU0800dGHvb7qs+F
x8XIBAphOJRScXt25G/7eHHrDQgc53a/gh7jzRbLQSolqGJqlAehvS9obLgkxJsi
VNKIYZ5zWPYY3w27EBv8EtIB8QJqr4bo8ErAp5xhJGCsxLFpoN61JxVhhpn76Ow1
a78vaodw1QMWI3VgNnrxIoxbauL1Qp4clL1iwF3f9M/Zo/HCt4BZz0yBBd1g4WB+
eq7Zjc/eoCQyqYr16c8xwvxRPCO8+JymMTHVTq6rVp7UhGkrgbfCmMk3BkgQurM3
5F3QZh+ihcjkBYMTvVo4JkAOI5DrDMCll6mha6B8w3b2mlSwJjEDoabNLkDBlzWY
WaQCgES5D+QwaVs4kOsumKklaTIWNnnpy2+HHL9inCi2D/JGSsux2MoaM+YWjBXC
q6h/F1AgaJ5Bj28H4QkSIsYGs/9JMq7K+AMIPpFnhKHUSTjVEw79glV0PgrIxXkh
9vmMgmRvcf3VVKoWjAD/rbRWPL6df3OuDbkU2R5CH7wiDyW6xVQMnczqIV5T07Ai
819BvZArUrN7jXOLm35XW6hhBSZ9XYu8IvmDKWyH8ORrEg5Xgnjac2J1+OryWOwm
wBxAtKvORfccnfJhWJ++MpHKnBfI+CDVBPm2LeR8gYr5zw8NkDG39923Sbp7BkGg
2Z7ovgqJzpxEIH2Qs6Bl/7s5Ji6vtX3fBZJz12Zt7EMzHlPNGtrCLHOFD5+AhxKu
a5kF8qhF3AHzLRAqid6SGdyDoWwzbmnst1sDjdC3hiM2W/cW8205CSZYJCABBCIc
R/0LJrziFc4VIV6SQlZH4xxHdbN4rHt5ICACp67hTazlz+FXgk4YGibuK1PtIzgY
UUSuIWli7VOxZbx0ZFGr3U1MxhmsmK6svlug5HF78xRoj2cJiNZds7kgWPzrrvMT
LMflBcJpqdxAYTuDU6+1mm05/GakrUX7QBNTsZWQfzaGYKF5R8BoWtUkCO1tpoQH
6lDiYOpr/GMh4lmT6YT58QXt+kqMHCZwd9M3a7Pvr+Z9r8i9Gvs8SyJ2RXrHPJeI
6ke+Y1zDv8S8SK3YQ1oiU5srV4cK6ixytVp8B2oll6Hx79KQy+RXQOUxWXVgLcir
mwypZKLY9Dwks7Md0yv1GG9QjDY7IEowa0wZht8XbIyZc7oXIfyDTR4qWkBO42eW
QmrL7ua0YLt0SfGKZvOezok1SF7vsxTnw1TTPVUCuwXH4HxcG2ejjqDa1Qa62RYp
JOLJcbHpe+ij55BMadCJpj8WhZ7PPhyxVVNLkH900cU8tKuM32wAIF4h/ERejVUW
otU+U3QZMNLX3IdBe1R6z8of//CcKIgK85kYNlC4pqOuWbw7k51Fp5tfonoL3yFW
WNB+GewGlnucJTowk1Q63X3Z33/TxgwrntZIQCi2KD4J8yCmFeXvGj2YMYqJO2xv
Ow9xYAo3joEwTEUvuPzFOybn6dtaboLkMe5cvV5BgsOqwf5BxFClDbgapTb75inP
vvI2bJW8N5lpoxq+7TaisUJjrYjEdXxdMFR/gnqxlMrMPA5lvHJ2YTyOqpFcfbHf
qg9voNMb+3XxDn8CspX19CDNv3oS/sJn2h6W6fRPTngIlaGPvdEO2ECPCSDCtPxw
PfLmUquowDGxC6cQwmnsz9Dl2Ao9awI2ZKtucMUj0x/7kE/CgQagX0dFqGPq3hro
MQwVnRa0VMVolcHlmstFv/5E4GCvAhZ4srkq2hTMvuhRHPreQCs2jJjFOFBhZOxm
btZ351bp+VJoM6wQ5T/KPlFgatz5fqlCxlEPf5wejM8tuh09A1Je7S+Z+IYqIRr3
0Bok/ShzW19+yhEHiL3Z6ClYIlfWcdJoh1HIA+lx7quVWU9I3U9z8niie5QXnMVZ
LqUcDQ7QU1zknsnB+Udjd/ts+tNDA5jtMwbH+oyFowbyVY3Hfh8ljn2/NPKsc5K1
Ju2CbqF2YelANmPlnq3ZBlPH/U8f+cMqVw3UxTnOCZqS4IVLjmzh/LXFLmyNfeXX
fXgXiufABzZMWlzrt1Shm3nwJuF/snhC0CM950oN7QKRdqW26KKtIT2Hc8+9ksMT
Ta2b/JYjNyGDEHM1NieEhIR4nH24a6gliK77+K+DhYqM2PX41VsRf82GJfJgwON/
Ld7DYDbf3ETPxurFRgwShIGTalWmAS3sw7INZmuw68hjuw9njwv3tBjI0OgBSBD/
nWUngacVSVk0ur2Mm9JFb2jMnmW15EoI9zuuGJfZ+f8GEa6IkE/aXslleliL0YNK
ZxDgChjhEKw83m0y18sGb7CAmG6IY0vCmTs8Jcrq8sRStLwcKDrBXwZPTyrs7vn9
VH4mj+sz6Cg+HIQJSvPMIxqdBWDR/8aB+/9xnItBP9o78vewIw8CdsvN9hhaJ5TR
FUiFP5LFL5rLOlmYCxa+kbPjV61RwrXc5kj07NU9+ArD6VXDdp4BZvgk5AOFIwZi
tCGUDko8gkpIhwABe9EXypMyL4Jr7ddLNGdp9KY8icAFi+naXw4V2IZduqbsKcIr
Cc5pfJvIrgcA1cfvhTfSoFfKCKy2JX51o1BplUsohFWvpj+hy6QVC8GvmXZaLkWZ
74Q3/ZASMZFtStOj7HGEYf+Gm8/JkMGX74ojF19kZR7RSkgTFKnnEeeaeywqFO9T
N5M3NPUPsKyXCvH6a7j4nOtRVsP7VFmWWoWs+6FL4y7OGG3KJk180d7bVRyX5GSR
Ca9zgi3YL76Pcsjhlie7JwwwkHSS08fNfse7f42u6EC08LpTjX1+YHJ6X2GmGx7Q
Yux2uDH2E1AX47OxJo/m/V49vPe8o0lOmB1WhKrgZszQ/Z2hGmprVtLmlrtSM3ME
XOWghsTAPLauqM0AEh5PO8YaNcJDEIot4zMYPw0vnq6dFyggZN8CU1/dotTG08MO
MabsUzxmtMwdi9qChTB5dx9l6StZyGiE1k9k+4w7aYcBIXv6C+2A00aFfc4xSu9S
xzH7u4UuO/SHqg0wHIqwMoUMJ9ks2nwnsrpwh7cUXlfjxypUr3m456fmeE94J1Ze
r3qDJJ1IO7KghMabA4b+8NxtfscMGKQm8ZRsSxJz/WLynfCH+AyS78LGw6LO/Mkr
VWf2phQQMjJXwR8uRgYO6ESsgdbqUydb4cJPV8PTzLZYvOWeQmFC2i7dKq/ANlXw
3JOTmfinAqYBEayCsCePfQTLClQMTiXkLYQWsVhJq636dslaC7PnaiBfvQVVLVxm
Ro6UYwTIgCncxlYLVLla7rWYngzXYjNL85XGZASCtjfrsYO+EQMZdzh1Ho9FFCIc
kp3cceXhcZ7h6LKqRARytyvZX11lnwabdYDOEP6jGsnHidC6egBYImQuuzViANYy
VaWeomz6xPruJOoBwfygep0p/s/2gla4h7X9y98PzDL9nDjSaNm4u65MxPaaVZ26
AduwgtUgwAAYRGWaB5O0NEsLLyXaVoQx+M8PXB8QgH+x6TXAeRrvzQpoFmlvZb78
y/kuT/tviKHtYQ9suxnhZKhipfntIXPVuCUB+zGx4BBEsn1jTdMhE71ik4dQWM8n
tmIbZvekjlBtDaJbTS02+AEkXJBuUQU0o7Mktg5h3JN0i/pmnPC2YnF228kLcvsZ
3Z2393V2YQ7/RQK6Jx/bipxLGWmpkNl9/+aT6cLZ9BShJvM+K1ABbnAdN7VhBRu6
xBs8owuvKH/okgbRFlHYKNEfJHWz4bH12Io4YT83Rn2QfenaNe8YzzsgNhD3hkTd
8jQSAwMEItKex//ixCVtxn2yDWBu+votOBQLDW4uzbQ1P3dFNtFN4qDduSQWgkb9
Mj1lpDeQ0zV90Sof87KOciHiZ3/MXnAvijAHBsptx7Z9uoVhVSRmOsDqiIEvxdG9
MZFt4UI54GrdOaVVXwz+nDq0dKt9wBwh4DB4rE7OtlRt1jwtXqLx8UwKAPRW8VFP
2Rc2VXdR97iKFobIqw13kDVyGWIeCwyFh+1GVEf1PZGJgFaPk/mgOVg8aedtY/by
4HRePjtg5gFNZcOSzZBUUntfkGDY9PafGfGrkcrQYO2uyAXgs6hO1Sog6IfyOKBE
d7qnL8dy6mFvYuCuSjE6M4tYR50s75wu9MmR/7ASRfSP19Xv1ylBbhuOA66IRGex
bumQJ3CVp11ygk+VWKeCMYb/tJL/ViPZvqsOulwwcheCSzSR6LKQeX6RXm3Wk9ZI
yls4/ten6/d2tOtnNSM1MV27ZQs/RoP625wEQq4LQAAPaxpaP2sx9sh8HlQiG7AR
5Fa6b+p37GMUNPydrML63CFxDeZTlWqOkCfPHcA3Xj0HMk0ZfPI2p+B2oFMGx2t9
NKqNvxDPopJdpe8NSD53q8HArtIq+1jgCyIcsK+X8fJVWVyJPnd8mnh/b1lA9KBR
X+s1ev02841p3eJzram4RQoarevjDAuaFXCK9pd/B5cqWYBv3Tf6wwO20oFX2EV+
3PFkwcua6jioLUVhT9orECQmZrVZRhMO4NVZRS917dmcP5Xxi3X9IsroIcSTQikJ
MRRI6siS25wj9xkLLLd/vQLvHFTrYpOLqXFkfLqxzmknLU9KeWW7YGNSVEn7bZTH
f9tmsxw4JcHNa+3O1+YHupzh7Bb0nUfvyluu2DpH/uUJ7WAWAAl4A/CK2S2msCtK
GlP+TScB5xkCYcrNf4RYo2HEHFPWQ9pM9kU9qtz3G3dAuPT3gNaSFaoTHmXKkvUP
xUFZGNS+28NP0XY2e3VSt94q8YqZZli+rcWYjsG6yAO1lJ2CTQQvvnxJ3FMZ6Os1
eubrRNdKle7yze8agbMpmJVGiLjQ+5F0q3fEzShYx3L+bw5FkiuMoPET14po5O8I
00nQEmsrsPhnnNQAdV9Lku1n4vrSugqRuUErDsITd/xJdbt9iiENkDmaCf1H3xHf
sx4Islm2RZJGUsouSwesh5QQ2JelvhsCNfk0Nx8wCMPZdH/SdAu1+NpAgYUiKo8l
ZcFzTeZGoC1h0YrQ9Tc4OI1aB7Mudn0wHRZeHXs6G4mpstQ2rWAdadtqZWsX0kIL
7F6WBbq8S+EqFYvpvI/d5sNK9lZGc27bp/UptVqi5+C2DJ3fKXMZx2F59J25tlgd
l4mGHiMgE71s0u/QVx44qvEznudMxWfP5U/zSde8kE2UaIfNwweoJ7tlnaBRC9Tw
HgChmutr4gB3WwTVQHKI73RC2ple1jQEMdOSfN5BZcH3yx86FDNyoQMIhjub/zut
o3nPJ+cXKUfGfsop1BiEYXTLVd2JH0J8Otmt34ImHxxRwNO2lyxoo9DI9OtVD6lc
I57pg9iis0iLbYwrGLcSitgh8tTFx4w9il+KiQdy9MuokUnvDA9/8ixqvcWwcQE+
b4EwW3JJP9MlqV2YP+/Ih2YK3GBt7OuaZrHtxGVb1IhsTFSzB6TX1rUNupnBfcy7
upFp1aHqhH6WMBFooSotBHeMYcHmfwolcC/b0PJNWGlXAxFEA8DYc5vOig5EKKb8
Gy54yW376bGlHrWAMggtbF5B9pmVlGj9VD6Cj3F0vsfBMCypB3fMIYYLTavOknsx
+wv9h/B981PoSq/V1CinlG6ZPa2wKc8HeuuDKDy7HTmi2Ie5vrEE7w3Q+WqVVVGI
fd2QbyJy3/mPrzQ7KIGZPSHMh9svHJCet1brgux+JE5WD8wrCYENb2zNqDUrksVi
4BiwCXIoQaBIyZ0I7P7Fy4qXde7scOldfLGZzxyc5PPuB4is0zUDxBY/xhUd7C/m
rpchGnFDjDIBqakegkFS81PH5kVxXqrbdfWb1MzRZOApd3OeOfAKTi/v/R4ATFkP
KXwX7T05eJ+fLXTdjaFPj34XxllqQ/vBT8Pn8G+UskX86jgKytkTLQadXH7/VlWL
/pWSp2K/zTdiUAPFSWLRa0vIxZaYeRzC+ykNLIgA38d2dkl4z4GJUIE+sZHOCl8e
ulmEoshOXzA1O/KUr6ZdaJZc8hOSet/bCw/7bgtJPwUjT7c47STdmW80wyrcXPx+
MWw4hLXNUNI/3Id6XMhrsQUAxtgAnLwk85O6XSvAoEq/WsBjRoDkB/atYDxeiNMJ
Q5jaX/0HPeTjX8ZpdKG47lblhpPSyNvrME1ZQCFj7NEENDPS3ZNjqGDF1mUi1uFI
UevY2iU9fMGr6zJgCTRogvDroOpeW2NpJKXTnahpj9PcEkWpBMDXE9S9dhA98sx4
/rEL7RPzA+m/PrCISjXi0EGSma48+30OQ0vKpnki7wjsiRtOV4wEtYQXAYB767nx
xv74LWxMZZlsuP5A5wX44VfgC8bQ9XDDAP8/c2r6RrAyNpO59IPRJmW0daMeMUHM
RtW2Ve1FRYCIr8ksq6+J8zXK7YnWOV4AanTdk3J5LisUycEQCmGY1LQysB06ynVg
UK1ENprGZ3gAvDn+DTUZpI/enmex2f/4O1gEKuvwt1aS0OjgFMhZyvoJtwZMswqL
El6v0EamYnKcTuDbgIBZ+i57jbEXjYMAxvnU+g3h4tBaSN4KVP20qp9FGi3h0Sj5
wDCH58dbOcsi0qEkxK5awbRhJycxeUKvLQn4iHHwNtyZOEepKdWJcvHdO64tSvXa
DkRCpj6xmNvxrrmKQXvISvM6MMi4pbPliIyOfxhPBI/PImhcJITPpCy13ESecF9c
wRzahWUPo8cWewonrDaYu/3JLef1o57I6a1vJsfaYpAxudY4aWIn9lgoME6RMy2s
NwtfBQYBTuA8WpYC2X0Gl5QSqGIAAZ8Fgcwo0mfMt+sFg+HislNZdPDABdX8zgg5
lI6Z+hsZDHWM2vxk0yIyiBR6DMqgRbykXGeW32oscaqUavkrsJZSlqoS7ykqWe+9
Nobr/wNcNk0MIOrh8ufFvYr8AXh8oZaJLUlMN4xccFIyv3EZ6QSQxaDdj/VUQtHZ
ZHLoV1sL1poOnWJT9OCtNyWSrUeUaDZq3V+f0CGXdKMTIVQE2xrk9agtOfblGXGU
/F+bcirk+nX5Eoq+rbadB9rgcBLu9K1xMpcsoXr5F5QOEXoxg6blSi7VD02BtPfo
RifhSWr+X4fp+/Sz6UabDCBCljrxsJawWukkrqsRU779n96n63Nj35y7CxKco2Mi
qavzvK+WGSTj1uDYTBKRL9V0wX5DIHu3p0Y+rqvg995LRz8TgzjXE/bzmjy2meDH
E6CWQO+x3HbhCWpvgZyHcgMyAgiE28lTyMNpxkkY2AgP+BOsOqCpUBV81jpNnVyd
44qx8Tfi/FGZVLhyKINqGbX35OLQ4vd/h5g7rRCHZ4/lKd0lkaLQIADcyUaG4EZs
BTzeGTOPCCWlKoqc87F/WIgwn5aYkU8AwQS2r58TyIJHurBKN12fjhd5N10q/gyX
MHAaZAyN/9e7Q08axfbJ1zIeIGsAicHs+FklH32pxIApjdy0/w6SHM+Gb+cyN0Lh
po9eSMghXmL0JLiD/p/hg8lQpBsJNugDWV96oZzsfY68CSal97l9pnCPaFfyQOpA
octBb2e1WL/qy1lgTrsVEIHeFXk8nZT9upfzlqywKgD+rwqaxKsP1L36G2oD0ngA
8DZHfMAvHZEIXtnp2C7In/XHN3ZZqJmRK8yLkEGSkVfFwPZSQo007IUz/lhzs4Gc
4v1R6XnNWNwAGC5ETtbA3nZgGXiiyxfRz+33Zr7JJbWE4xUcNB1aT8SDisrAzZBg
/SvdAuecVH8Gs46RdaiTEUqgBO0XK0cVTkM1jH6RlVCBDe6n0+iPBLE3qs9mccBb
iePcRKoznKVKHAlSYYfQYcJkAI6vLgeG9mWRoJRGhqC2+zb5ersg74KjePWWNNMb
ug6Xv4YCzME7B8dcn3lcZUES/JgmVMfhC2viv2wX/epOAmSbjz3TXLKp0f2ggJkP
Vi018s2OHAZm+daZg/gr1QqCq0xnxzohlTP04X37QpqjwlNRutn1zzn6CpYRUIsv
+zxld3OOzeeS1wIaqhTJjGeBjlBoxEkYjQt+I9CL8Gs+Lf9M6cDVGVNDzM/qMRMi
getkBNpMHvV3tV+2pGvU6JB05F7lDqMrOhoouKBbe5SOKP9MwOw1dvuZdnKob5eo
hip8KnQMlr9++sS/mswVgx5oa+mkKMbcClPM326zF9Afm/XwMDH2e7LwWNIMvLxI
lCw6BR6BjSz7hdN1Hj6ZUG+O5uslF9g1PYkpSdVjYIXDIh89XtwncM8Oo58LmGkH
Uip3KAf33GsWsxguD4JwNXIv0WO2ntYbFz1Dc/ofDzrvJ7UbvhNlSCSK/3m6f0p1
VMZLwtmrW/TAJaKhlDgaZ53ijVC1KbDKzVMzElcH1pqR4AflS9hOVQWcTUXdiaof
YB+1xxhPFOwThRop5zk5rHxYSwC5lqXQOpyvMqEYmfEzPmy/suegT8jO+lqBlN3z
qpUKkIqkalxRrE+WWk+wuq86PjOrGVuFTwHd1WqnkMvIjtH6cReNbzgdmyqxpv2S
2WmGX0b5HINzfw6xfn7Sgym0yFtTaVaUa/xrqn41Wi4yeIOZ1ctDZySbLeW03edd
uslK5f64Kljl/xGzSGFoePG+0EqHE1P/es1/s3vXclvWRK9j87q+GvI783N00Yqo
nGWnvctGPbhrHZPlZp0LnlFOUGhTurwLKXbTcwkdiC+MfZguHx1gmVQqjU3jXlAw
2n9OkhCJ5ncPs2fO4R9lHAaOgC3BrCCyp39qPq3ceks7D3/njB+tUXDauGoo/y8R
KsBeBDzRnppmu51lORDeTUUGxD2SoDv3vGGJbM77CJLyFpSldZ6/IKE5MkimxAbD
PhjMbU/3ljax6pN/9KWgNJVT1hAwQGuegdl7gpDiaSR044vNJ/eEZic5IGAmaMRf
wjimHcGgPUJ5pL6Zu2Eev1ITCM8qehNpF0o3vFKlrK8XODJCTI3zZ3qeplck7hIB
cvmLtx5TUBYCX7XGXJhnkp2eiRVwQ39FbHB1qhRyAkMWd1KGk5RDk7JkrI7bwc8t
+IEaREhtPg16HfnVopoaghq4qoWoM70QW+4jt925i7vNysFnlD8nUzrJNSGnirCS
0GOegCZnkgA7Fq5auSpj1+vjh8lFmTWkeAac8zO9mLU6rA9IxSaVwOe1uD9F8pbq
um7E3LPmawQw0qcE5RvZ9h/iW2/gVtPGMXdkIX92T7XBoGqfoiwqtVGQfYeed9yD
CEcOkYRktBTQ9a+J6MFDdE9BM+SOqprBsY/IyRmm+ilrARpqbQ7FqfzWthBL7guy
fcdxNKJwSTyt8F+OcJPUZtcsEvTpr//eTH7Zmmzr8vBIi84yqkdXQVH9ELvVKB5x
uVlimdLi/mGDApo9vOVXBb17zQg5pB9fJ9OSPm0XBxLwIyIGZTu48DKgqPwN2CUI
bthCRMchOKLgozooN+oPux9vFkKb4WagV/w7u9UC5mKAHZueVCXsLylpcF8CiKbY
oGA6JDc8kqurLQTlaj3FNtXe+7RxCiLCnMulGeAU2FAAw5ZUu61IcayeT5p3CY+p
dwL7fWG8ULpxJ0UBa/FOS/vBD00qNbAApc+w8aYSuJ9QOykkzzsKAIZbs8WDfIzm
Z/C8FiASZAiWxqiFZv1uWcqIOxj6FEJytYD0sA10kQIHnavefhZEBJw7h9FrPkLc
v/AP3oam9s4g2zdRsJUZMaUk/ErEvl5SBsenAa7s6kfEw/R94TPpLOmJwtQzNcwE
BYg9mX0qUh+lVJU5T5oWnz1Dtl4y3MqMTpwXeEow8Rb/uYt8qVemRyRubAv469VZ
ezsMPpIZltnjCL8Qsf8ImXOKVHY/LVDI2P3hPvJTwQw4GxGN54EReeCWpXy17u5Z
Yp5a3P+AAdBqRr2BSZhnPnllJE/m31lIge8sZNvurthfs2ul56V0VWZji6ehixMr
hFp9Z86vNkICm429KhckPOJumwNL3FSUc1rzeB4rF6f7Cvrrk2mLOTwAADisxS/2
7k2lzdBbzVhc1bWI0nHm4a8XxvoPj0ghS8YuEOvjYe/8z6mkdx8WsiYGsf3ugdX3
i9iENsMxJ2FeDIrE7wfuljFPfnHuaXSsCH/wH5aUY41mbp4Fkab3MnBcpTXj0+YF
Dw8NtUuZs7hw98RL8nwYvRo+3m3ojPQMW166Ht2bDzb7hkuG230QA7MMWT4BOd17
6hlIQ0CpXwf4+dPUZn1JbT4w+LuCs6NZahr+Ns1vZljF7mc38+2vNRt8ywRyZUNr
ixU5IX08ODgAWE4/vRkt/+nCMrKAWobP4OT4ZJdLftfYP3pOxj60ZMuoatihF1es
g86q5mdM2uwcf/p+VsHUzEl+Eq1QloVEkDnn6pawH2d3kv6bE6FhzgIurJVfMbK1
9caZSxxaiz/0W7Wp8BuSkRthCI6fy2OQnEECR1EnaNgVOLt1yl2KyuSj+EFDscXd
pELtEPIodPqb7M2WwoQQGMWXlq/5N4SdsM76mPEYq7gZMHiHOcFpgVYMhqu8LTAe
2tZZchuVPJv04brG5WbEVwZc+uXktbTq2jbj/fHcyn+5MUxvA85wTv1GZiOfRz5g
4erStEtzfoR/rz11LizOqEW6E4t1f6I45vpkLUhR7jWnfWUtWCRuIIq0ghxdVBux
Lr5LHrCtpvgUeNWMuq9o11cxwaDS1MGjsx2LlnFNKIKFPIn7IfYvJPgBUyLHD/l0
soGmLTDWTauCoXQPJgCb4Lv33yF3fWgaersmPfQknozhxuVZXPg8sgM+bHqNLSsF
ZqsQyDf8HKutvkJ1AjEcKB8sVxqQBIoB9k50OY1QOO+NhYVT+TxCJs3+InEWZYYp
w+h0u7Yhy4Cs/Qa8nO9Tb0oPUrErQaM1xsdsCXq/gBxQalAn3PiYxeGdIeks0g33
d31u5ymGcr9u/RWqhNl4WVI4ot2oum26Ffum5IDRwZo6UXs2rJh3K328nbOnHU4I
Fps6ys016zi9Zn4w0HANgzGeQQXW3ccLdGrs0IW1Nsg08EFyKtmv2FClgHyHyzSg
EQXLyisr1B/9siB6N7wuUZtuuryxNXpzWGl/9l2BcUeDxkdXoILjRyFQxvbSj3ON
kZ1LZ7wiYoaiDhjBDunURV5nQfAq+epaSxMLn6RDOe6CHKzN690O5aeXTLwK914g
qZT5TXkDva14Ol7gpoIrCC0jS7pivMaMumGk5Gc+LVNF6RviV1EE0Zx2Hgh+mdB8
kKASUVwHTdpn6FokcQ3+/bYcIMtkYrQHU+Pf5v2tZyhMsrgSk6kVBuCd8BaCsPuz
yUVvslQQW8co6RYXGfvJT5cJuWpSvdqCxpGdTGwNiqJvA3vX9lG/Ee88BhxROX7g
IwvUC8PPmPtBnMnjb2lba7KIvBAZ5N8ae0HVX66hNLs504oEhrQ247eKlC53SGJZ
F42msFYJ99sedU7MmwRWPJBjcx9KLnMudMYGSLNJIFX/PSFeBRGxc726KwNFQsDp
tHb/iPfZFST+mhkQVgrkT2nQWRWoEjWEO0A484+clDRgSwuyT4t0bIyQ/x1Ncraj
AdZwtN4+G8jXNaCQLf7/aJ3l2rG8wrI+iesWCkhE3ezBOaBt5w3jtnGU0Sfpv+jx
yyya54pxl1rctAxrIURsgceaArOZNpBvccx2c1g9z10GnyCuX3/2iZ3fp167qEPz
ra0B2azGv7byosMqDf1b7sceW9Iv9idTMQ/IhIhhRtk6g4JcN3tJeKMZGzQpgi2t
XLRGDPYdkw509O122fUOYeO1FJ7Y9Nk836hyzrsmx9QWuqIsptXKLCg1pPrcKDnp
IHZ5hsKvwDV+H0sa/e5JaV/BnOz/TM1pie4hiCRAi6FOZBkKhrxd/ARXdZMPvYO8
+bgcqiqb/vjd2E5CvheDxLCiEommwc3PNArYtuy6yfcpYyHX43YzUchGrRWEMsHs
LvM6R4TdP2L57IQOdCswxW64LRuo6bU4bvw1/0dA2GVopk3FwRuoX7EdHRWy7etf
TWAYjcU1anauaq9CVO3T2H9laAtx0cINS5tS3GAgIeeeELx3G+dIsV0J5LH5l+2m
vsYdUxMmiEXrXyn0plzWwsgDTfyGXolLIDwowaBDGm6y5saSeZGczTKuHReDACD/
t7EvHX0/zVHoL6UC63YfnekdtG7PHvuWMcKwGLE5mo6FTgQUqV4oAOX7kbNqu/nQ
rvj6WVqsovajr8tWyKUD6inIAGUKk2m41mbGjQ/orJbwkSAoSBJQhcexhQdxbK/I
IfFPLmsZKqNUC5qmbnxTfem8byWhl4lt8rbIoqKLxr7r63RyBUHz7Aa30hhIH5Tl
rjiTDz1kQS+1m3Tm3qrj+PQ52xvC6OwmVHMf21HDtHPVDAeSaon/Zti+aBp3xUf5
weyDBwI2qZI2QjaC1Jm5IYcgSPvntY9B9j7QE8vaBVLjVIWjxwXV7ngWEn0u/6wn
cBhkEV/vD5GDt1KR9DkE2wGDqYE+KCg9AwLAh4inx4OeyPPnbzvRrHU26f73rkCT
R9iPQDB/E6Dl5BSLHW/if89Lu2Av6pibJnySFhnHuK9eeMS/OTqhQ3hc3HBGeXcB
vasrizSBUKNjtZKkSGOqRrLF/iG9nNWb3rN81oPLJbXuB7PGAAjvpqrHGona2hjh
CcEUxCNM9dfkB23tvgjjNoHnTwxlBeijQW+i6Hl4XL/XP/1HKMbJrkdRbS8UAhtI
dL/IbdG9cJEUUlFYz2DPi6EfVRNuILjpgoRPDey2rk9EBGumTmXD61+hRQLz9fye
lLyxa/4vM3/YQKandTchgQu0qvSqsN6UU3X+65lnPSq1Z04Q/cgGAnWkjIjRPVNp
h75Ge/QH7lhnVPbyFg7wX6H7zF1u4Aeel7wwVQ2t1BD6DwOthSi87Iw+/8XtNCJ/
CZiEs++lJ1vBpdXrBlaDmxIsRjejly+mSqFl2k9l55BgCmRkIsNB7Wx3fCOv9QW+
Ms8A16C3MWOxViKqRln1UK2ZklsDCIUHw/QuS3vI6bl3Rzi4u2g6kz0Mnd6SRrQG
EOuvsbS6Auwp4bpYieAn1FQa5gbXZhuE/df7lvYdo+UrP4rdphbqMnu07mC7K2fI
MmDxmKxERmo8x/I+rUg9KSp/hp+eVP72BF7AVMEtakFWmTqN5J1AT5a9K7E5Lf0Y
6ducuom2QDgg/nQr8hf52dZSN9Aige5I0J9ZWblm4EHJlkJ8e06V/TPBK3xxRXO/
MiGfut4AUE4d1ihHxu8x0scSj7gcD/U0RjyKvrHlRZXaSRT9vAykw2qRoM0u/kcM
/nvqpbFwMLDMMYplNksMZmJe2G+eP+guF6L109t/0LXxVvLtP5mVEkw1R72CTCXz
uETPgLchYsCWKngXqi4fqnOiCS/adKLDuWzR1QzjmgW8buVaKm1nVtNCIYFdPke+
j/IzOQBU28SLhBU6fHzoIVJlUy0B9+zqTc6AQgG9uWEfvqkTY0moLWN9l8CQF0mL
T9dYIoFN+8jwq8bokJsLddkeNBUD2xmwinWSlky7NZo8CjirnzGpa6VXeJaNPtpg
esCvFTecxk+7hmnd/BX40wRtCADKCM+X5BGimNiDyVXScsmGNCVocCK7o8YAA/71
3eYCwC9m8HJ7cv21en+4AMGqRYJoHh76dIgrX/y+zjRqsXf/1TVSFFGerMdZqtQm
+ARhcPoeO6+lsZqR9RfsEpyLYDJPd0o4biM0u7EAw/m/+k3qu5l8BN9+Agn+TIph
Tlrkj7EYJR2hc9JAHelno0MfVHKw7HadS+IYX7mrFkUiw6fXoKzMlHuGHa3Z8OWz
3YNlLEhQZ5+HZ37kG/7GzEePbxpO/SGgGxw6C0FwXNQD2qE9CcmdT67DRSFn4Cze
ZQOnvi4R9J0docLfzkvJcK/nnL7SVA2nPMtv6uHcgtz2dYY9MokTDMCbTcjB0ccU
ez7iNk86tnbe2EeGIjIiFqKO+H/Ch/FRlFwm32otHmWeI/DFMaNy/s/eOLHFhcom
vT4uYHtAfIxm/irvZSE7xyjFwXjnoeyaLZHFtnKc8vRZZgAaW0zl/r80u4JX/y6y
gGRcc1drN2tzWfVZWuuSkDbf2Bpd9nUEh2lHgtM1K11z0gF4G2YPYYokDhunLCsT
+qtHB0kvnwdGmqhmUNHP+SIoSku/5owi98tEBSBaIhJM9H+GmgDSw/0VgE3B04l/
ilp51A3rlM3lWtkDy6H5Zho40KJpEvNCidR7BaRgekjcFfFF4ZNfMuRd9vpYkWyp
l73ceQlwEK96OXhKChkhycKgUwxY2+4MEBJ4hPZk12sbI4EkaSk5ciOwicU1o1PG
ZOJ+OVO33ltVsrWJRarbDWCAKvRcYmnLM7S+17qxhKgEu3IHkKitM5I5XA4CD40G
V5vfy56uap4J5rSFKD1WK4Uar4b7VeGdWCwcgoRYqKeKylxUxxJX2nyc28Jqg5xj
GUv/njdusFJJnc8dhNpOg8o5KRrDd6VZc/qoT8g9fgG/rwYf8W3tTIZ6LBr2S7VO
dbhZUpXOKStourPen/8+y0cICIcRiEyVOqnoKJx771iL5Sb6N4809JWxFbJl0n/a
NQ2TeheBQMJ16StgO9js4lj5MOqV3s68kzW2fAoo/rrfJD9Hlxm55AlYCpyINk5i
lrANtSE/fIhvWyAO3ipa0VbKXDXlXa7ypmm17mvjy4yLo5jPDa37mrV8z84I2Z+z
EAeo58NHuDrBreBZbX/UqM9+ydu00GXWiJdW5IlmKYZzGBtdcvolCF8v6tA/2aD2
h1dlJtOfN71yCE2IMZxXCYqjtkil7bY8hEq1b9PjRIVBeUCvBS3DabHjmJoN++wD
rNp/gZyHYxwO+ap2cB1z3cKGTNRayPmVJqdrZn+vPaE3oFnHn5zNBzphmXfG3IV9
z98tOdn3rdXKLvt58B+4j7DvOOroC0NZf6dsLWwczkjFiU74e2HMm/vFcx25c8FK
Mb40C8HkhJy16QYSTdi6sCdy2pH2CAhfgIkbdh36pwmYTiNUvPGxnRdraa0CqasB
Z/IEyPS4wIaWLd3KleKn+otg5fLNp/lURuHUAXxfoeULXMzmlCSdhqOTw4NECLhf
dhz+uMgvi2Z4qWarirCDjQS/JtNORtgOO/+sDRmO4aQYhjSojJiUt5lGXSQLg2El
1cJoMO8CDpbAVt8fT49orvsiwxbGACAFndtXTtJFgt36hEGzrSv5hlMETIVBIgSw
mNwuqDxuDmXrMORyNKGZISpKNELX+NJjFJ0A8SEaB1TW2MTk+1NAku8X3tEAaG6T
p7+NwDXGidhpCBNSj0O+WH0hhu+xV4V81xK/rHYz0Ljz0uRVe9S8Se72YugASoea
Dp+IfJK17A/nMeoYbrKiG/m5Kagid0EhdnwIbBNSq9fzQDfiwvnBTpwYj4hapYkw
m/COpzP7Q7du77NBHWTEp7X+LNfPqoBeiMSXV7CHctxJDZoYpNy3XdZuLTFgWQch
4bnY7SWFAS3hbMaN7jnvcy3KSlbV87jLAqpIVwaqTkKHnLAfcB3ZRt7wM27VD7yZ
KcLtTOhQa4h8gw91VEbV2GpTfMUFIB1giyIIu2T7Sl8NxuVcnptE2oJGAUgxl4E+
5BDu2PId4rXSeGZBWejqJB8uuvikgRNV766k7W+yVHGg7xRehFZnOstXMJcLTPK+
5wkG9xoW6BzoP5COwevcu3dRRWUMdua6/dfdCKQ8D38R38DkR2qEDZZpGRUh6392
su8rQmKBdMh1qFq1hfZQGRy6B9WCvT4Vrm9pHuCzrAND7eCRoNMeIiPEhpb3GU3Y
OG7Hy/rITNr7P96sPuK8q8xuGGqUe+l20OdpFVuPnsa9R3N8mNRt0N/zlCoDm0jT
B6TIxHa6H49NQLQeTg0kFi4rCyFUu2FvC2nYLiGMkSFXtWeFBWUgyiEr6jCP+vmo
KDKVDPSH7vxmQ0GYsFIfcgOthUmRxLtgNWKTwxYbsSlsrPD59wjSFzzI+pb5x+2j
EPn8nFfNf1umEX7ScagN3RtduDltkiiVFmqqhpbmZQMnXOz2G4kYz+iEFMl/bUPz
MO108+x3uHenNgFS+gNq8pq2Am55RrpPqJ9QtZK+UX8eiCvkzO8Cc/GrRxiin3cS
So71SKk2ecFmRmOMXl/wR8EqFLl+PLLcwKkoKVVD3jSBQ2ovRD2h3qeY4U6labCc
X4zyVq3Bg5VpSsOUmPudXWQl9mJQCz59V6uEXvjYSn0pBO5vUUEeZ78aCW6FRHWc
eCa8A9dWTHxr8S1I92koV7PPVVKfRHQN+lK2q2QulEmHur2eQrsTx5yuThPvS+jb
+pXH2JY3zPMSkwB5/AJ72uF6YL+Mz7E7CpnuReEji5sxtB7GchUeACujIPls9sOw
EjU6UgrcnxXPwtrilbLZh4tipWOBlB5rCwpSwyeMmPWXNoVvheAn38EFl5mX7LyF
1Xce+TxCj22Vdk3WpHoEpGkbVWJRsb9uAkRNhfE/jJMzka1iZad8VrcUgBOm6Lt/
9sohhONQC1O86b38LCRvs23yZS2LmkP9EZ4ytGWHbQsqo5J4clImvr3B722DG8rZ
7RF5IixvDfBVuEbKw46nOKJ+1AsZb0ONUBIoDOSM3NcEvBlSnWcpoPwiuJoYkOaw
NV5/2vV2J5a9C0Q/lyA3We/gF7ar9IwEcZ1TlKOQIKmrDiVx/+z0u/2rKbCFinYk
uZVnB/M4YTJCRKCPra9gPlqmEsLMcIo/Etwm3i18uuu5VlP5kZTfDMqTJ8i7ntj6
4B3MRl7ufAgFBVUJhdAMjt6g2no5wfMPE6ZLfm+8QuHpc/4z8y/jxWHmpXBh7QDP
8JZ6ck9yvLo4l+qDceBKE47TiLXRG9Kat7mJHRB78nhrAoXyH4xZ7WEND3oNW3BS
wsYhYxI2upg2j7WLJdKwVhwiFpDlfXDiw3LOMOl4uEMiVEh/SGEynoKCb8PmpKoH
H8AxYwypqyPeR1ahfOwRsc70lG0E62ozoGqGLd9UxK9QroTOlTYl2jXSTUT5u8AJ
hKg54RmFb7HvfjqFp2rNLld80TbmpXeLguhCWp0tH+mH8zQC4A1xviffzXVF3jDn
bm22uuzfLPdHF3NtO1RnKQzwnjt5aXjf3Xi9MbNOXojEVgZu5ZU3WNxFvYRcdnjn
raSwW9XGWl4sDsCoF89S5JS/MMx70rFgzK6klUE239GkteBlYPurzSM3YGkHdNgN
f4l0Bl2zn05hfFFjNNllhAdEMNcScKV5x2x+R/eEzSC7Gpp4pzaRLAKFfAA5L/NG
OWcNZIR79ZMWZEgs6mNmAk6wtbQEK1zVN7DDiu+6WX50tucPE6dupNdHfY0wGi/A
6zLFax6YesdvmVPuJa+WGQbs75qm5IZIarryHumZ2h4n06y55G744L/ll4Jh0CDs
aqYP8qv9jrFQGeLE9BSj4h034fmDIANNzqB2Z8VpFhqYryEQMlkvd3B2sDvittYE
iwYTdXNtzjPso7PvcO2hjRpSxM4uKCBjK8HnuUHWuhyi/Rpn0bpztiEEFc702MTW
AvdwtYb8YQ9sEQy2Y8D5cIY9rFOUnLg9PEDA0AOeXy1q2g+RNc6N4Pm5Y/ZM3jSa
vmX+uPvz6dRraIyOKcx/Q9MQbtsukBZKYM+8K2bzVBp4IuNr0NSIzn8dAlKgoIWD
rbuSwx3hQTDTZ811ySjORVKuaQ8o3cZKuZLYxLkt7tPbyTit498moCKbyWvqbtYH
89knmGMxL6AdKJOGtxja+Hh+/XRcsvMu2Znth7J9cXZR79/5tLS8PXWUGsPfOzl5
IQMexNdpA4iBCCPFi1UfHx3l2A56gm5PswzD9EV06Nm0xSqjlW3adJTkxkW3RZ2a
KUzc45tujW/NXdKY46WY6VnGjvondAdVfqFONO3T2Q5B3azqmjHdcu5EaC/eiUVA
KFWUq7UiwxniUAq3RThAMMphKhsvGIl1pxS7zcEkUr2wUK0OqiNNLt9QY2obPOSw
visG5Q53xWA3IBhI05Cdu1EQFPqjAgZtzcK5TK07thdVCSrhxZ4ScWUBjc55xjiI
2494e7lzKTTkJ35x0FFdqat2sJaOKcJljAO9LsdY02QU2aV0nXs9nbRZKgoBon6C
OITs5Jwd60J7KuIDZ2OlxbjZHUYhqWgZGQqifsu7C80aT3AvxQz5yISxsYpbI5SA
Z8bazSX6XwFMMR9sR2f0RslidoPomMzbPfrFe0yDpQFyqKlzl8W54ddumK0ssWwm
YdbSS4T7O9Xz0uEtRXbLuoQcq6anodcStseDvaKc5tsUnstZXVWEkzhVviCPLmJ+
NtVnGS5NIa5tHT7qMqb9T03El+jCjC7k8FH1qtwBOm5+DZoPuAazhWgLQoyXCztu
wCagy9R5G5mkln4rO9K9D7VWFbWnTQ1idwVjYz6fX2aEGKu7JpKQUG0EOUWzohsr
kpuIdsTudD7PAFQPvdJox4XMaFhus0DGCAoa6wDXxn7WYnyDuypoxsSOJ/uKl1qq
iCEfBgh0wge/3Y9hT49Fjpdkhd41nCCLD2boLrXnS/y1ZNyw4cEsj1VCyhBAtn6L
rRQSvsvXSBhGbZQ+szlYhCan3d2WIlt476G3uKqo5stfhrKBWDTsUUWbAlUw2NlR
263Aqssofig8i82OzaqFEBXpPNVsQj69Q3j7puDM9KxuwxcOx5aB5Boi41OBPTiT
87dlKI9c2wX7I08FPYEHPyFiWDNnUFephi3PSeRQLewI01PbXawcjTc7UhwDEDY2
ezLFvQAubcQdoGYhm0DMvpQ1jNiYmTlWf/xi6YhOkxG0YKh50VkgS6Ewj5txX9/R
BKmfSms5Pa1WxzJC2yCYONwJKP0hmxVcIuaOTK+C/ZDt/U/ZR1XZWHKUTbW+u1jy
D0kLD9fm4oEsydHnIlpn/Idq7aEbeu1JKYzE8OwLo10Ed1lPgsu89VzRWVscbfNE
gyo6/Is5jcQX+mjdfo2JTUaQDi/CVXC+nxzhrSxD5pg6HPZrWjHZFVhE3AZe4YA/
iBqQ/6fYjCeB+MH/lECKNvcm6H6mHX+7SfOgIn4Pw3HlMq/FQSApC7ET2YG9dVgu
lVSHG3mSDovwfzZJ96c7OW0Do7KZKWf6g/vcrlxefFZcDBjs3BBP4JjyPP5vS5rR
K9wXELoALVe+cRiE9LI8DjCz/3W94dBA9Qc5m4WTPGOLYeuqKOhmJlCjBTa4C88U
xETQL5Wri2mNpQClLZZ03XE8JW/02mP0SoThu2wGUuDz9v3uQ8lghsNZTRGpOCUx
2NLfnb7S/Zbgo68UNY8DAuxzSfLDzYuvi6c8abujjoA5LH7OvDrA86N3BcAYlz5o
dbtFXqRRoC9451+z6t9ErooOctEKB1J0gYClNVyvSNFJgAmfEYV7BWukmS/MqMPy
wjOxbFUqDMIYqWHvtL/Tw663LRTIi2tlZN+0SBZvLi3kbUmtJgpW4+xry/sAksMo
RDMOnO2eKCzUXe7+3+pKcudcisoO3Fd9hkvJ49LK1QIIjV39aHS0iNiFyJB02hMI
HFm/fT5RKh/1CA+D1f8mwj585ldTCc6jbgNWBLlj7AS8SI1KYl6ioBNRLDFFQZOx
rOqZBbr8nT0hxCf1VvMvhAN4CxihBLLABXU/ULz4X2FF9yPc6UesRY4kWFiEd3Hp
yWv5ttNV14m0LMd1FSFRLQdPsYgSok1rdXxKEZyeiduMCagn+5CvjEWLMy6SX2fT
03OT9BKUex44zPzlPKNTvMK6p/0VLAoiozkN1CYt9tgZGCK39ntM8rdpxLV02IXx
7rQ7MbymwATtxJjoirCtJhQhl1OUX5O7WCdb4FiKQEqWaeSNREu+3qzbexd+AAUK
2TKFyOEPOHOxirRVjr5M6ztvXm2GGsmTc509xnACQEsY4C0j+u5VPnG2gZGbrXDG
V0mx9riIqc3qtGQWcQ92bXKPyXw7i3lLOLkPcQX0V36CpJwACubntOwvfAy6IXJ8
f/CHCDXYFrS9ruaqqMGfG2fmXlqAtkbx7sw2jkESh2x5tnHWOQ8JLjfwg4nLpYPO
L7EsYdXnhSzQYx/xIGZHCRxztiEvKqoOJsvTXCbUSiHmaI55r6X0x8Ehe4gZiQND
X9G2FDj1kzjHpTF08j7iE95BWsMrTvFCaWWrzsKyUDXZywGqRfu0dhuA+7DTOoBx
/Dx3sRBBV/bNNDygjBTUD3GLxsH6uw1EN+QiXprpq/HfonNEYHB/T/zYfG9rguNY
doboPwg9Jjtafa3k+PZin15nagWAbX2+hCOT4RyB0JIry1P3Lne4nnrFkMASIjWL
dr2Y7YHybcKtI4Ai9mkGD9LbukH3j9yMJuxKVOD4W9iEPrCs0cHB9FPN5FfbaXfJ
9mVdw/VAeKbT2qzIDoE4fPOBGBUS7qDdKQ3mN/y0LjapWtMl3M2WHKrDCjlMecDd
C3e+lV0++Y398jkVkC3EpR6LAyRXTOu0kml5qc7X90zci0fLJEKCNHAPlS8QseSO
n97dclHbVJjjp7eGCkP0IbhdrqFfbrwnjXwueuWMa3Op7iMMqAOZ5e8qUVpRWnDQ
C6mSxpZUio0XFiahNTrnq1U+eor94ivbhq5sIL1VTrIVEs5jeyUqryCrsL4GSuiK
XCRR8j4Uo6w/+DZo/JnigK/vamciNTeiT1qKO7bACK6VqxZxlMVpyGDuum/uko1L
VTF0P/blUetlxmFuRrbxcfhi6mkberkaK2ST/5a8B7bu0NL1VsVqtCXSJcdvEAhz
qHvosltzvaCm/KmoQ2j2+OUs/eISALbUJFJ/1DVC/zvkSAZD0E5SH5UtfvoPdjrY
NRVuG01Qe2/3gBx0KW1KBecVZPsv1RhzVE7roQRUJ9Q1E4Xq4BqPQuZRFMOwK3Tr
am1rO3P2hXQ7ZvuygeDjLdSAvjEMrJ9+DG9jMc8nZXPttlBm4TsMxXmoqb2tBLAD
luVR+MY+WpXLBL4IoTHH90gSOoDITGJabj39VWD4V31vaEMrgUO738Tl54GHIjNe
VHRsQqnW9jd5WX/UjT42Ygk4EMcvGyzjcv26nsShbAzMFajlfby5GD3MAbPZEA5C
XypZcy2KLCCgE8WMVuYI+PAek0CeWC/ecwCQXEBd2hTOjoA6sfmjPcUuuT+qN/PD
vUZYRgkagKBIRy+oh9HDpDyuii+ur+8pSVmmkdZnjBAqtBNsEYQBxrzxJqjlngGX
hYvnWOsUEq9+0Nlz5EPotMJPBOZYV77twHa6ssqqWoUPyCoAgay6Ae3RwAXHIrj1
4xeM/iEyeSSgazZK4aJPVeG38xmE1Q+gQK6MCxrFybzJDnNiulddmSLG+zvMJqYP
2eSUwGvMlFmCCDHtNJcb4aGfh4B1r4co1cVjLjw85u3kUUiUIerPI02K4EnoCUEV
t7vuRGeJTXL3vrGWZnHOBzpqBlzWch+uWzrS0EJQTZsfkooAau35oo9+85qOUkXL
OmnlgMChJyt29IPsF+FDWbOHV6NqKy+qEPk+tEo/Gn+pmTBuVFfkRQkhhrhvM0ri
wd19RhMoIGwDLw/MXqbXhaHA9P4Bjj4KGorBko/CwddJmSXSSBAcPTTI76bmBfy0
DDzVskYnmGcvxBHbSuNyF5IjxcgFmpM6Y9KgnwNrHI1fyYzqYZr+/0khkK2apSJE
hxvaxXfvgH9qajSgE27O2AeT9ngQWx0/67ct6AIY7XpbhLent+r5JGJf106R9fQ6
4lXUxHdc/HRpBlrwE8v1hlKxSF4f0jlvRxcodkye2zMLhvz5z3ev/Rd5UOUPmvnR
mKOGkcRAjIFkYNe4t7Y4rycyb1yajvOaD2r7q8+nl+c4BO9t3Dgf37wELQUkCbmJ
l04kyHgymTaypZzR31bS3pU7/GIIKBYGVmpY9I65LiUU8ekLh8bB6g1jpIZp9dsM
qFcF9QQCzaHpRybbQZpHpDUEuQ9Y+fI4sGiK/u6Q15W3rKIfwoH9NB/bHUA+Almw
gmHw2UVmVEjNcBBN76djYI9nHLD3/FuqFXdz6IKyG4eh88gQjLIW44mukFQePBFM
6yivJFQqqZpK+dit7zKwqqQcd+CAPoNlaK/2YRf5v4QDwvQXB6AH/PEV6/8ZwuVH
GhDcIX4EObwPMrSnNOVsUFKLhigMNYpgnWwlCqjKTRcpD68jzvgX25TjYW41ykvS
jDwOATctM6M8uneDWk8bzqVJARR1pRUK94LVdlHmYtheoR2HXF6KM3thid0KqEtI
WIQjhw9MD6Bhecpk/xjCgq5Xs1qHlaD8ChsMlWB2NHOipvP14qD10WZw4+DX5zxP
d9K1LbBQ06xyfA+9qkhrvfvWX21BX64XvnWjHpbAy+KjUsS/oTdjsCwhLo5DXAck
uGApr0LqQyQ+zyBxzc25EBc73Rfd5HKkl3rpAvEa3ZHMRFhacUj4jI3NV0vj7tTg
/90fNMilPHtTmi7DrtwW6S4eLAHV5U/UH3PNP94LGuENsPMNnNIcvz+7dPfS8ORh
a7FfG+9Tzq19lnCPWvlnnhI6JW6lcNi+83LyLowitBiTes6fU3WlTaiS4d5nwlFI
Gzk/bpMl8v1DFJjvb9XSJwf2/8haIO/DWvl9Zj8KdaVH4QnLcKbsbswodcg8GBfJ
Vb1vfy6ldTAKcqWW859kpBHzFxQ3GGOFdDEtdN1CjSs4yDA1lwD2FqQEVRoRaftu
ws7Hv/L8wwx1pGq+W3yV4hM+ExEBu7WEnWEWWO9W/xf9GBD73xHpo5SIvF61qdY5
O2enAD3IBSSYV6ARYnDse9tGv35zurc27o0Lsd/0dKFw6lWnte7HMkZE/lL/iqjO
c4Nx4MI0GDOSZefW5LTmBUPNh6yx6M/bNYb/Z/Qn9kLg6jqZg1+jiCa9wyUzZaYC
vcq8WNlV9NQoBvBiunX1dXdvLvpYqeAFXOCcte3ncPLZSuNuL02j3RwBWwCyO1lT
uxmmssjfGgrYuME8GchbEe34QSGGS1YKv/BxwijW6iK5Xldgkgmqj91jgMBfZDjj
q+V0Oay+2xR0amYPaT/zNv8gcWrRcuZGVxmxH2oLpu+KY676JAxaI79KuL7h2PwV
rpVIq/tRzr4kvLzfz9GkqGCBJygDOA63AiSB1XPJYyoLcMH7P+uD+pEqK7QCEr8p
fAO8vSguxbZzJfdMeILA1LQ3XKq3v+PDIZvL1u4n66y8q9mb4JhwPWizM4Nmogtk
TAfygDFodg+gAbfC/8OvlcU6BUWLA2epbZ6vOktY0ehC4pnxCgPgq8IFP5HgGRT0
N70wgacWoEmbt9nVk0lQBonPC7AnqwFxNnsDhrw9U9+g+dhmbROsg7BPsMvbIA7p
iPh6PnqBM6xijBKs8EVN5/9OJZiRYq/5eJigmwRpUlj4EpycZiaOOpN+bNfIGxuL
97ej8J2kClsA1QYjw5Ifq0XE/Q7RnCQ6iA3MuPLWxwI6BBC5PlT/ZJ0U8HVCAL4N
SoOFSeSDvIIR9W4Yv09hCOuBj87334tChVj700bmoCUurcqdGvJlIuzJYveHC57i
vfmjp0Ub7yM2IsnJ9gMsZhC1Xihm3dVhzI0IsfxHsMKrgmet3l1xmifgp0LMAPv1
CcXC30LGnW1SP9H/K+mYmeyC626hVk+CK5sW7xnfKGMrOeT2VpGloUQ4lBsMZIsg
P7ouJ2a+44co+cnpod9D3sjB7VdKD1OTqsMON090eU1SHVVMiL7w+zLODOJUZ5vM
cAiFOLCt0cQ4232PxzEYFqY5BoubK8hc0gBXsChG1QGymSYHHoadbdNaP5iAGNDA
cRcCOCxmWvn8imtrXdcVP67P9ZDF2gB2oW7zE2338IDms1i+/oTABroJ30HYbj2o
3ozX/r23FP/njnIt0MkzLEb19U/L1kwphGGUQ+bGRKVFaX7Q9g3SR3Fnvej9MVV0
0+/Ji9ejupZmPvP+I3KWERThm9uk1MpYd84CFmbFVfgQs1gB9GF5neIJOcB0/og8
iiqkM/J71FmFAZZpeSj/pvojBjo18xEgkYmITUjXRTRUfU5AfZOnQFL8LsYAZonb
b01SSXhtGN4M9dZEZiGhLN4d/TaS5Y7zk5yeklg4F9zbZ0StHkD19UkZTj36NDxJ
TJdbzKy44uaWC8igw8O9bOa228fSmTXuqiGf+zRl+NgT+Rzlrx3R73VTwCdlwhYI
SFeG8HbMf2c0sv/qgMwuG5jjVGd76U7enkqAHkBDn+R8sXZy0+IrcUdJ6u/wySBL
1ko4AvOjeu5onXxTGMkLt6CPYkGeDVbvHj4SChJder/9X65KZzLKk2Np+lDbTmLl
2ex368enP83j5b3yD3J8tgjI/V9fBKunBCfsOW/aYcwFSD9omjfpKzmkf8c5YeaP
pL43akb9HtFLpzdXfsnYFnx5Y4a5J0AGt/xBD6oUdHzeuokj1vQgb+rwfvWfcT8L
bhjr1s6OsRbs+nla6IYfqt3YBqJ3fARn5b91WSg2uun2F3+JiSpZK4qGT8H/PtSd
keb9+BK25oLfmqYf7bMLRvEJnPUE8LAUbIUrCmyMF/7GYZM+/xKha2sIMC63Tclm
JtumjK/lELZQxelRZinYEYBnn+hjw5iD7mrd8g6h8maqn0Qq/rVISgzx/2fpaQOw
jzyY570hbkTds8YXUhR7O41N1NpNCF3UCT/EDD4BAcKEFdHbTsOMvOzy4a6J0Hwv
ZpX/3L7NLgWccyQbE9jxxFjOWX7MSQ0/cR+06SYDRjZORSfViGyo2lvGvu6qL6nS
8uS0aEw9WwyKNgR0wJByWOfknhnp2QGq0aU8Lzx6J+AnXlNjWZb20Rjd/E2nlpI9
txGexhuYwQl/BFR6vlPRPQaFe+tXtyhJBN7u6elUDRlhmCmSov4A70b0II0HiBCY
4wujewFoFarG7cr2Ak8yTn+gS5T+o4sZB7rqdWtfKXu+H54Ql2dEZkWptkDTxUS0
s8b0ebyG4NVzdeeTVeHiVhVd1+cxVgBBGob/GHCYxESE11VM36ZOCf8RlMmHD/Sn
u1ShdP90inQ6GNHnIpoCFDIZFQG9161Yh9v5jJhAeyTs9wiY3lkPMFWSJg7RekWs
NSXZL1mQXCvUxWZ79e+hOegGyB1gl2qKrkp6pIppQm/a/BVhBOxKOEyuftH1P4IY
75y7ep2iUb3USNri/AP3ZkX9vqxRXXNWxnGyS1EiTnNHge1TxS8SSWKHLhjE6ozJ
DokHOD7JinsxZ1nan/ErPBxdOmbdEiX71/narGgKU5UDKTMI45abOvXTIt/jtRMa
/I/4e962flS9E2XxTHJb7lWNii+n4RfvkdpA89cDb97XIA0/Zt1EWyxRKGCyAKA3
d16XrG+AXhC5YIsqMQqQaAjq40GZUHz5xNtogCAgScVqi4P9ZILMbkHpm/5ikjlC
x0h1a+cgfYdhNOmJ5/fzSO7aGpNzzgZ0r1v3CJIYu5tl1nDrVUq2MxJmah5nt0sL
lH8ELQKrglwrvzMz+REa4+nly+CbK91gKbGiKyP2V0fqTKJVZ+VYSIqStvTUHPm8
R+hhmuxXGQgpo6RmCK20UTxXDeVGl9DZ+Ac6ecPWqDZZl7lg+c4+mxVmO/FoerwQ
+k9KUFiBCtr5TmKCfeZ3o7Tct4KzEB5DI638uoT2qSA=
`pragma protect end_protected
