��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_)!{�J���Bh#��\/-�N�}�5f%25:Q��Ȳ����T%I;�x�f���zZjC�њ贠����<g@�6�[hxpJ�g�EҤ����G��(�����l��ݼl���Oմ
o��Ty�����1�򸳉I�$�/�G�QQh��X7�y���x�]�C���}5=��g�)��k���:n�f�ɹ`��y���C^ڧ\������'JQ~!8���nh��F�E6Ħyc�B�~�x��Iɳ���O/�V�RP��B���ӆ��z������-3��^ڝ��Hv�������XT�d�w|P1�Y�H4�I9��zf�F�N�_���Лˍ֚kV�s�x/W��}�d6k����צ��up().�F��ŹB�iR�^�@�D|�k��_J�5�HCť��Iֲf�n�DwD\Y�c�1�<��@#Ŵo�L:ģ�N�^�80d���8�
�����c��tNL3D}e-�vt5��$�Tho����I��zy�bHt���n��6�"�6�w�)�L���Ğb�#w�LA��r��x���l�MF��^]�j�t1��C=U�a����D�� q��#I�>0���a �5O�8��8����э�^Mť���e�� h��3e\����g�I�㬱�w+�7�Eu���>�=���G��B��+��/�*N�,=
)i����P��n-�n�a��G���G�Mp�-ᾼSb3�;�}��C��S����~��������VO�E&w��j�'-�=g³J7�&��Ң��愑���X������А˭E����C�Y���y�vdPG�ƥ;�SA'�i�|�� 5+B��f�����{�d������Ɵ�2;CT�C�C}l�WbC�}��0F�3�����+3�y�A3<�eΗ�4V�D�^Y�m G����(4ŋ�hy��W}�x;e%lS�N��*�p~`Pz1�pu;V��gj莐2_���v�L��m.ݑ�aX#t��%�F��w@�l0��D�(4:�ʸ���a��"Jl��V^��	���l?^*b5�Zh��n��u��gݟ�y
:��ڎ�k��}L�xc���We�>�:%�3t�a�5|�!u+e����-�3�* �,��P=x9�QA������B�N�^�^�������K<ok�n�P5�J|�5������n���'H��JY�<N��2#�v����a����E� Vc��zX_U�E�{���_���$*ʰ��)�$�4èS�d��%ȥ�k�v�ɇ1���+]0^�Y��́��%�ܼ��u�QSƄ�rw�����j�t��"����o�Lz���tc 也@��$=$���2��M���>@1���8?)�_���`����(08�μ�]�i���|�U�(�7��P�˲}1!����LSb�v������k���"m!�]P�x�%��dٕ�	��a���{ԼEލ���C�.1�_H���(@kb�̻�����C*����W�������"j!OC-]���^�£�˰(�lqC�+��me}w�jNչ$c�����nL���O9�|�m!�|L�}������(��R�?f�"�o�Qe�rf��T"]��S��~�>A�?�wK�P#L�K�[�W��������k֞1b�46��-S/���_bs>/օ�|Bn�̏�ǰ`�MD�Դ�(�L^p����Q��/%�ط:�|P�O$�\�(�&R��2��(|T�LlIrqTcSᥒ�=����켩���O�a�3���r,r���E������1�A6;wwTbDꨣC�b���ĩޥ}0ʂ�QZ��\�i�9S{��D�$MZpg�g�	!$�����C�M�ĸй�%�����:����,�]�'�S>���-��lb�C�x+\�z��Np�(����͸Q 
����i�����B0bL��h�1(�~{�/%�@�r��Zj���'���Ho��"4�y������l�e��50�$������6-�v���6�J��=簾�
E��YJ�>�yr3�g>s�,J� ��z�<9<g������!g����{�5�?N��12����&�f��!s��䅶�>���P�h˔ȃ�]�U���T�<�j�P\�U��:ݍ�֚��^XY��%4t�����]�-,��.]b��g>Kkl�]��A8�w�y5��I��� ��З��/ҙ��A��a�����:���l��фlC���.�zY����tr�i�aR ��P�w��f�nwp��������Y%��x�?;�9$]��I&J�c�Wv)��`���U��4�t������.��8a�7�lg3�PW7K�ą�'&�Ei{��#	`����j��'�db���f �{���o���zd8���e�[�I��pR���1|�2���l��MVs�WM��N�����,��uM ����`���M�v�?H�V��NKŚ���������)������8��|��=(c�jb��N#-F� ��(�3%փ�{.֑�g����-�Ր�n//X�O�l1a'o�)7��0r?�����0���Ȩ_�/q;s[��WhR�|rߑ.�V��������&x?(;��q�q�qU�p�+H��U۞㬊M۩��~Ynd�:�}�Uœ��Q�U���KD���O��������h>�7��B}
��撽��ú�R���xz���,s ಀ��&���q,Vdܠvm'�DR�t
LǹC||�*�0q�G�vޱ�|h �P�Bn-7P  �@�7��h`�'):l���yک�����NW�N��5P�d��8춟R�M�OG	�`��#��_�����N�R�I�BղZ�y������I3����՜l��2�H:5p��4U�W۝�s���ot�,{�MCe�Ѭڹ�Ʉ���%�L�V��S��6bJމjCML����USe[ɒ���#r�LPgo��ߑ��m�4�IV����j/��x8H_�M#��a�>h�uEU���[�z�0�}@[[=�T�L���;��'�6�~M���f�CQ�"���i:���'��"|�Ϛ���s���(S�p�hnX�vՏ4V!N����s6V�8+����R����Df�^D��-���W�j�%�^�QC��X3��|/@��3Z$j5>x�h�������w���\{5#����69������}�q�0��N��ڢ7��kH�
vgB�g�oKT��kdC�'l[]���(5�rH��0#V٧�ћ�W8��.�O��y����k�[&B�
���'�0w��RΥ/�U@�
�rN� ������0���ϯK��C��zg��-Py�.X����Wʊ�������Q��l.8(HM���=���2��}�9�w�gbx&�|��߈	�Nt�p�����s�Lw�bEWi��}ֱʴT>��:	���3<o"ǭ���ŻI?�Q$�~8�3먿a6��O�.�ʉ\�13Q\���6T~�>i���ਂ��@I�Ɣ�yR/�Q �jVy-����K���v�'yn�8nE�w
eI
����@G�]�����:-zLީ(��Z�@$W'��yt�x�?�O�.�!q��e��c���y���B*��#6U�\�ؽ+��\�r���BN6��EBI$�~�(�s�-͇C;�K�}!�$�+[I
h�&���q���r�u/�0^@�^���Ik���Q�}+ԇ�9�2����.���fhY��a%��P@g|�
5�bhA."��G���xD�%��m�M�����{b��n)��V�Ε})�o�M,Oƭ�b8QzAӔ���t��o���/69p�g�.�7�R\�[�M�$ٷ"-ع�; f�+n%�_���Tk��~�R��_Q��*֦��L?�:h7`�OC��Nxu�{m�P$� !E����
ݕ��������S�E������.���?���آ�}��4�au�M���+Vi]2������5��o�s�Kr�t���6� |iwi̝�i��V���)�x[R�q�8��y���;b�@�sD\����NU�rd��?�*���F�����V�U�������W�Q؝Z�W�_��z�>�Ȟ�}>�4s~íBē�������Y����������!k�v~��i�&�-�����Y��&D��׼4_IP-i�C����� � �&��������e6Ub+��qc�g�����e����N��{�M�s8J�ߎ����F�T��)>F��Jx��F0�KBrɈ�C�����!ҙh�|����&h�$׽M�Ol3N�c�?.�f�vG�J�-�b��� Ω؁�����_ߢ�*b]Yޡ�;�����6�ߔ)�(�#���}q w`B|�H��߇h("R^�h}�Cӻ�e�p��Q7mTo�h���JOk>�5����B�2��Mʣ{�6T��t�l��J���`3���^	#�v�}I����/wʳ1ɇ��j��_ 4Jb0�9�atw�嚾��&IMf�Jg�Q�l	c�M�X�7Dn��4���㰄�H�q+����{[6��;{�f��U�N��$�]tw?��9��E`�r�B���x��3ְk���yD�N��7�J�Չ#�^�V{�����~)mT�?�x�����'np�p )Gp���_ ��A��CN֙���O�{�_=����ov��n��8�	�N7��E{��r��"���=V��B8}�e��_���a��Eװ�������:����JD�O��r?�� 7R������A<_�s!�{	��W2.�=z�Q��ĳj1�5��S��g��m����̻+
/M� c�龇,Ԗ��ȝ����Zl���YI����C#I�N�X:�����5
n")���1�����9Y�Y6$~�D�5�X�|@���>���A�̕��/�����Zlݯ��`�{�-����I��m�}��(!����r�TG��#7%H ��MN�0���!vNy�'θ>��rw��]�����;�M`E+�^f����U�F2n?�2G%��"���e���<��n�~ �A����Q0�x�sJ�ڀ��Ĩ8a�]�m^���.�XYѡ����\a�%�*�e���q����v^fE�RK�XQ�<r�����.� �9��:<������ ܚK()��S��vE}+j������I�ݚD������\��Z���Qc�Vn�M^�Ӻ����L�!(M��I�M��P�re��ÎS�Iۓ=.;ڃ]VA�q��~}����s�79-��l�+�3?l�x�&�?W�\M����|i^� ��J AB�s��Q��LHW5(�n���� �	U��,��xQ�viPޮ�eX.w^m��¨���8_v1)���Mo�o�$;���H���:ή���_�M�@JX(!m^�ݤ��A�}��7"Ŷ'_�fS�K@�:ܦPc�����q�u�0��|���|JtVe5���P�υߓ�� YZ�%�R�D���7���n���ʊ�A6����&I��@�]���x��˝��H�F��v�b��Ȓs6w_�hc�j2+�7���, �w9o8�X@$����G��К�H�R1�Te�q9�J��f�F8l1�_�R�j83U? k���E���ph$�=��f�X�ܤLlv��[V��P��cȎ��I�%�r�����n�i�7>�p%7+�����Y �?��1 t�:3f��q��o4q���M:8=,~� &fˡ�� ����>��R4��S2io������r��J�0|�_�0C�i���0��)@b3X4���[��h����pM���*���+@P�Q=YƁ�1���$�8�����%}���?���~oo��F5Rq��z�����f*'�����y���FԼZ���"�H��J�\�h�d;���S�l��H7�@��Na����L�n?2�����p;�>\%B#��e�һ�>�$/���{�܍�ȍ��/H���Ɏ|Ρ� ��#� �0��a���\/U��ϣᣜ �:j�HR�X�Uv����p�>�s��~�d��a���8J��)U�&��hL�6!���pe�V[ +1kt�[�����t��A�E*}9���1�0�KC���A��Ţ�%N"8���x�bW�bTD���Ήw�I��#�H��*�?�^˗�q��Z�����mNǘ�䉮�˻U#��5�R4������|)@��{�q-cU��Ҁ^�5`&�:��(v��<��1Co��Vw����0�D��?[���6���~�����p%�).H�o_L ���ܠ����Y�y�%[�Fx�~����˥��(e51&^��F��eεd[I�THIb&?�
չz�Yr�pKe��ƮoA��j�&Yv$D�4���C���ᰣg���\�{��dÊ��B�q	*��A$����ڭ���k4����U�����&@ϔ��*�΂�q}�\�����&�����"�`�Pk^���6���7J�v�k3~�,�xv�9��}u��G<B��MaM�ʉ]�1
�A��m*%����(�u�Y���!�bש��,�������x�G�gX�q�$L�FTc2���n������X��U�Sr"z���#��͹��o�T���Or#jI���|�s�:7���梨�F���b&���Z��2J	��󄳲L�O�sQ��Q�lhW��8��?b^����9.��r����r2�Yy�פ���Ig��oG��&jo��T[���Q�m�I�l�	܃�%.����!Q��Ф���N�`��%�x8}<T��|�xt5溈�h�8�����nE����������;�hï,V{
x�W�A.�?��Ϡ�[6-hK��,Bk��ܠ,Ŏ�S.��,|��X+Θ��-�YA���K�.�mpY�;�x���B�����ט��.�#�{�p��5,$��cҧ�4=,��]�+ |#�EB�~̔<J���4	�a00qa#Q�I�t�F��d��0�+�P��9`@oK�6B����7��amJFF�B#���,���B]�k�t./d����M�Wǉ�c���_��=����H��rq���_�7&��J9K��#�!C15Z�2d���˟��M '�E'Q�r@��|�(��qD?�B��d�\>���tf�&��
���n�A�Y$��]c��4�ap8]⨅�.�X�FĲ��pVw.�a��b<����k_uR5�_ۀ2�u��1���i�i ���,�u֯�F`�~��F�OZ��di=�QZ��4Eō�%z!�z��.���
w�&�뮬[B�É��V`&�(�JHh���@���4�����E��{�f��W����L,$��@K�ǀ��4�kӜ��C�o�.����V��zK>oGh�r4x���v������S�����9�q��uS��#���}D��zX� S��9�d��-���ƍ�;k,�x�H�_ug
_|�E��>+�":�O��0�>��?C��ݼQ��FG`��d�̷<�n��A�Nk������'��M�6ŎڙSGW�
�'�t;uj!s9T����	^N��x�$Tx����^-W������g�>��M�ůɅ���B 	�xEg(�J�;>WV�ڐ:��Q�9�8k*W
lo�L�����@�r_|�����F�fB����V0)��B�K⾑γ��}���(���ɭ]md�n�`,�����U�{y>��֯����Z���:��_�@��'�D�;�6�jK��Y���o�w[�#�gm^���F�<�|����� `�2�;�C�i�B�o�ꀬ�OɆ�}��Vc
��Kӫ�l?�t��~w��e�.��Ay�:c��9rn�nt�(�.&t�E�O����]	���ئ�1�H�1~ �p) ��Z.s��K�Y�F)�U�3˅���9�UJ0>>:���*� �=@�X�QƢ�{+�%�BAn]�4���|�{�.�^�?�	����7s6�8�'Z$\��2F��w6XH��������t#6Ea���.���8Nh��D� ^^-~s����S,�`�r�"/�o�/��C��N�j��s�4k��`�������#�e*�Pk�����~SW�X��wrHT�=|����z@O
�#�\3��c�Wɬ�u�����p�kx�����8�Y�UF|�|L�ʳ�ie��`�xE��;h�04�@*[�s��>ndE����Y�{?)�A�9��޳} �?D�1�MKS�d[��������l���P� نl�ѹ��8�u�s�9
<}���s�3��L��)���w��t�0��@9�	��3ڵ'fb����$;�
V[��i[7���ю���.�"eZ����|��j@2�h^�p��D��� �+�x��X���"��P�	^�ɧ��0��e��
���t���i��-ҽt�^��C������-��e6�Q^U蛮�dǙ��}>R`��n0X 6�����ˠ˺6���5��k,�R�f���M��3�1�V[/�F9TB-ޒG��
 �)v2kP,�-����55�uy�Π5�1����cn�%@��ϫPo:vw��Ust:�3vb6������4jX؞��7�\ݞ�9�@7�}ֺ��
�	���%�9��ʪ��rY�������d^���.e�]���(�W��X^P�h�H���uݎf;.{v_�b�l�/���b�4���N?�á�7�?1�znA�P�G�����<%�Ml��3i��k�j��+�n���~�$���B�e[��/^�~z����v�3o���~�g6��W�-R�0�3�xK���Ԝƙ�i�
���x�ǒTi�
x�؎%_O�&���d�������xґ/rg���k2�X�~X��n�À�&р#]�ҳ�Pڸ�u2���J�c˭��:�X����U�l{�OF�%ً�`���5�@A��C!
�+N��SͪȣW!j�����
������4X�|�q�R�߾�PS�C��"f��[���i 5�B�nc���~*�db��l{/��-ކ�Bk�$U����6�$>ِ5���EM�!�]��	x��t��6�,UgZ���6���%���l�=5,w������U�@��Lv�[s��g_���ӭ��Ӵ��"�&m�o�D��`?m=F�E�v�����a0֔��Q\9
� ���
U��UV��ኜ6����{�eC���?�.a���=����&��0d��y�h��G�H��-z5g��/?� `1M�V;����~��-~jhΫ8��V%�(����+��!���Q��00�>�{��C��.�晱�&����͠o����mMk'3P�W�l��T��~�	�M'��2G� ����3N�T��@EK�����<t�H�^:l0Z6�Y��7x�>/	�N��ܒ�S��xp�K�9���:�B
�TY�鼌����JeT���̌����)�M�E�iۺ��y��� �1����d���@��Y�Gd��Hi#��'_BG�t����U�T��7՘5��hޡ�6q�+�\�i����Bn��� ���W4��Re!�Yw�8��x�(P�:Z��0=-<��!��5�J˖�DjAӧ@��z�<�h�,PTpeW�8�5����Fhwh�֠�JXP.`E&��y�G4#)�ӌ'1��n�ɺ�S�Ѭ��."]df�]oK!�0��Ҟ�@�7VT��!�;���y֘(�W�����)�r�W~�/{�Ȕ�)��Bݢ�������;1B�`6W_�~#�+O��6}A�(PS<�E�$m!��A��z��2 ��ش�c����  ��B�G	?�����o�d)�nR9���ep�u�k�A�ET3C�9i5
�� 2������ɸJ�fT�@u�4����G3Q���������0��4�չ��l�΍5vtb	�¡�X�Qt�b��ZT�fa6���(���"=���� ԕ�S5��S��6�*9@�(��x��`Ʌ%V{0&���[��Y��X�ph� ���e�UE���f]�M2@a�`�z���%��(\.2������O�@&�j�,��/����߮d��4�$����О�D"�r��3��~��D�������z\5� �Ȇ�����N�V*6���y�L)ɑ�v�o�fF�H���srꐯ9�tZMc�W-\�P��!��?��LƔ��@��]u~�df n�!H_p㔬.�Lx�W,����5�P�[{��YlT^�C#�;G�XC��PJ���Iܼw­�
�0d�y�=��h1�
�wz��aZ�Sx��JkՂ~���ޑG���
�qqc>usd�Y>��P�r�\���ɗz�>6A�y�Ȱ���R�ss Ð7aOV`��d��UC;�~���pΩ��fQ��uF[�<������(<\fP��A�㖄4���h�[E�=Cq�8��b�Y��.A��<���I�?�1��+{�Rt��q�$�5�N�Կfb�ZNή���z���ۡ!0�C5����`
D' Vs��)�`�U��,J[�L����Y����҈j��{����T:B��*A;�����`s���G���7��ɸ����,�-������� s�>8�X$������Ǫ@�B��(�����)c0#~��"�@(>_<y:oAO:���H��1�oC�F*�6�� �(�͹��:����?2B�dӴEt�G�
��@[ZN�9�޲�ם��p���a��*�Ŝ��Χ���P)׳@�/BC��Х�ח��{T��+��k%��_L2UR�rG�>ʣ�$F� C@-^ě��af��a�y �	G���C�!m�μ�3 �sh8���r/��|O�#�NAv�i�n���:��]W�q�N�[�8Qv�L�
� �G"�e�rpT�M��)���i@�]�� �t�&\�@e`'xzy�.+�?1_T��g2Nt �5�����@Od5m�z�`d�ޚzv��#��֐?{�)`a���;`��u8Qv�Z�ć?��'�!�C옺=%{��#�~�c����I��*��&�˫u0ӎR�L�,��k��~m��&�DU0WN���7�,��FH\��<jQ�^tӥ��/dװ���������s<�;vq}C�{3��o����u���{�u1z��s�e�9��K8[ų��B�6���ú�v���"h�I�v,s�p�>���&1	�]�)��Y���~ٲc���P�ķnT�M��#�gs��b*{G*�b~�%y���qW�pam	�W⇄�Wez��ޗ�vO1~C.�I���&�yl�\/�OYꜤ�p�+�#h�@p��H;�y�����ұ�7��$���ZWj�����#Ea�ʊ��턷%����B!Ǻ����1X� �3=v;�w"J�FwD��i���U3갷:lѴ���{?$	���ɷY��Bi1�}t~�2gJz;|���z	�@O5z4y�����@���=six��t�G��ً���<�7�"G;<�簒�������}�"��tm�MKD�g�(�\����D�g��p�<����U�a��<Ֆ�`/
�2��x�sBu'��?���sF�wރ�p"��v�C�aUq5B�W����{�����f���[2�'�
��tFa��?�l�M��2�`|�?B79E[�,�Go4Y�Q��}�����̗hk�pP�#s;�<\����@~�C��2Xl���ba�g�<Z1�9P�?��_����h�KW~��DS�[c���4���NmN]�)��д����~��*�j�? ���ze���i�=)��+B���?���?��x]d���VV:
y�z Z���kO��:QD��?����Y�A��$�
��lM��tWɪ21��+�����B�޼m����O�7)�{ �ef.��zCU��i�h��Z���\T-VZ�������$�e�� ��.[�ά� ���c��Փ�1�v�L�j>���Ab?�m��rz�,GV�w"���dX��.�8+P�	�艈$���\f�I�j���C,5�B�O-�s�m��ڃB��E�>{4��ז$e�:����M+@��)�``����z��:��WA�.Yz�M��^�f��1[�R��Z�Џ6PؘV�<�f86Fa��6�ˈ�<�#��}�tv�z��^��_������%E�߅'*o�$^�Je6�+q�-s�sp�֎�I/eJZ���ZUb�!�d�M���C[�$���
Mt:Q�㌪��)F-ڝ����o�b 6�&@�1��D�~_3	ڛ ��R�1[�N i�����.�\ɇ�NQUJ��m2��k�,��fX�i ���\�_u�T�Ɓ���X���ʛ�sVYY|3��M����v9���\
�f�{�uJE}�ۊ]V���>�k�q��?���# �c�?%\�j���;���נD҈�顀�g��kx	�m���9Q�ġZ3q��ʷ�7I_��e� �p�t�̗��q�|�e$���5�>2c�ҏ���'��X�#*��U�
�RUb�m��d���J!u�om�����"1j�7� zd�OUK��܅Տx��#Q���oQ�������)�͂�2��$t7��[�W~05Nj��R7m��`.�%���gs��Ϯ��s��[q4i�B��_rY�X�G۵����{t�ɹ�<�U�ne�䨪�4H���ewB�@~���z����ã�LaIL���ԷgN&���~��iH%��x��q�xe����K�}d�Of�T3,��X۰�/�ν���j�0��2]�T�,���'�.o�c���PQ��ܣt�I��Eg�D*��9 ���!Y4b[�X�z��O|s-Km���ˁ(f^�N�pDi�{��V�sȑ����2���4��"g��<�g��q�V��'�����\&����)���\X��T�-�8X8�96 ]`a/<�#-�%�b�܉WC=;	��fi�U�Ȋ����A`�ǧ��p"fص�kp"��`����j�}�[��1Aq�W^��z{����[ �/ԣGh ��GA���yC����d�;��[@��E��^�0+�rՠ��oDܲ}��{XC�22�n��ͪ����0(9�5�&��+w�����+����>V!6@h�I����۟��}m\De\6�7n9�P��7��a%�XԴ�Ƿr������w���m����MA�F;=�@b��4f����W����t�GBn>�k9���S�K�RTO��^����.Ħ����1��swj˒��m>�m��%�pu�ur�ӳ��<��P���>tY"R���&f�ym��l`^ȢJF����"�.�#!��0e�պX܄���Hϛ	��ŗ39��ρ7���UƖ�+�����l&��"�<
�f�eF_��)+�Tn��W����2m�l8��<"}k;�,x����]+�491�3X.���q%�<Ɛ2������*�v1S$��=����\���������1�X��x���D�^ ��҆�}h����9�;��ל�q+Z��,��^���"�ݎSЎeڶn�(����襘��]��k�V�u��T�:�QN���J�《�D������|A`�)���ӓ���D�5�r�vO���7��.粣.}xG�MUe�jBr�%n�	*�^�V�o���O�7W'+'���{y�G�=�O ��;ɒ�
Ӝ;wZ%å�/�^(�thnmᠪE,�Z�ڣ2��U1I�y���������s�
�JMk�xT?��(��&�s��a�<S������S���aA8r��ROV�͵#���`��E��R0���n���o�(c�{����z�C@��� JQav�����S���trEi�4���d�Y�Gnm8
�~�t�az� /k�QG0����x�t��0�b���YOxd�]�sdf�G�UsJi�ő�ֶ�N��@�M6p~�S�NQ�5P=D������F:<��Z�LN���)aJ��9g��eֈz�@`��=��N �#3�	ڥ�9�p�oM�� �d��e��6�����p'��G��% �Xb�����ԢH�ؾ�<窦u�0�,ޖ��Cv��v�_�c_ӐXǩ*�;~)��C�t_�� ��6���S	.Rf�O�^T����LB_%�o���W�>�s� fc���p�Ii�0�!u2`�@Ek=m�5�	�y�M+R~Y���/4mk��i�k��xeQ%^��oz�^+D������ϩ�%���(�tsK����|�_N����n�zig�=�I����#>�Uҭ����Uw��^k
����aU�L�	>�K�X��}�b�e�M(��}�m�N���ܜ]>�/�3������ㄓ��9������?C�l�:������@�Ǟ�^�[��$ᮍ���˸:��TW9Rf��n.@���k	a?w����k�(�軨8T�wO�i��։�i�r�uΎ��/�c�����9eGƆj�`��nr:]ޯ�؜��V��-�p�s�=L��p�m�:[���$�����y��s�?�H05n�<�?U`p��`b�JgH|0U�Hk6�L�D�*SI�a.1��8�r�a�C��<|fǇ��_�Â'Q���!��Jaj����L�����1�rˬB>~���D��ߦ���Lܚ$�G�E}9�}Ì�x;��"����f�����y�-��2}��
}��;�A�%�$=������%�͟�g����ѽ�f�v��U<�?PO����#;��ϴ�c$�BD���t�N�݃!H��A�ٷ�A�e*������l��򭲺xC�����6hߜE �/��y�h=�ߍj���"���J�"݊4�#qa\��Dk�(,~�g��K9��>]y�j�$P"�Q�?��Ġ+w�S�c��a@�t�E����B�l>�e;�A�\
���u���8j��0d��>�����J������$��0��ι�/&A"��s�u�Kdݏ�{����/߹a�'��A��p9̠g�^K�( z���� mAyV>��j"�ɺ%x�)���e]�l���v�4�g۸��Vb?�Jŵ+CQ�xf�l4V.r��t�Q�-4?��%�_��Y���Fp�?fے�ru^��y�,*b�~ݝ�d��1�W�l��Ѵ 8�.�1�Iw�����w�����&�(lP�����;�'���kWTN
 \^���S��)j�6�IvP㯶��F�~�1�h,�N�Q�X!��Lh��}g��iW�kɀ�I��*���=W!%Li����ڸ%��$���Wj]��F�=f	 ��ŜPV%E�n;�_�F�*{�>��u ^7�5�b#Jv�
"uhUV\QÌ1�v�hK�ȕ���jtܡ�1����Q@��%�妝��'y�n���r"����m�G��g7�5��Zs-�J_�H�j��Ws�z��nT�:�^�	[��J���#�<3hFo�x��|%ȸ�Uѡh̛.Ź��2h1��,!5�C�Ǭ�1�̏�Y�f�Q�2��&k����E�@���J����|"R�n��l#�57���5�zg�& �"�i	Kl�=W���b=p��*�<���G�b��?PI� ����)�ӄL:�Zw����q��Y������;Ĝ]�͸ڇ?���h�I1�ܮ1y�G��8�m��҇R���н���j�1��ރ	����KO��Qs&�AC<}���]v���kY���8�1Spr�u�;ӓ���UN�bu��#[ ��o��ިRꓬ�on[��9��%�[�+J�ʎ4�:Շ�V�?��/�X A-&�B�6Q[��G��o�{b(S?�T�݃�NJ�F������s2��'y��sԤZ��^�^����{�c;��d[N�AvGv?/���_�(����Ur�v$�G?�L"�Tz�^z�g��N(㟫T۱{��������BرL��+?�8�˻#ޘdm�u������Q;�%���������MB���Hc0>?���)B�F���>_c�,T��*Kfm�X%��+�MCq�����z�x�H��PcQə�%�����c@ŷ�u���3c�%o6�`�fD�JU���_�4�c*F�]��-��9[�D�����)�0���K��ۖF�q��IJQw`3��SR�������l_��M��Io����V�-G���/�	ߓU��F��č�̞�������Yp��K%J�mh̵��OG	~���25���{V��w�R;�8�֧�Z?(��� s_)Z�0tW�%�
d���!�� ��%�����nn�Ǹ��p�uzGg�ʌVO�H�>ο���K�������<w�e�,%i�Kk#!�z&�7>��z�|��5y��^�n���
}Aw]5qz�#�O��ϪX6'L`�I�H��+��9��
�,1p�,�{V/F��J��XR�����!Z�Ln������˘���M>��|A+��n��.�p[ب<���#��$y�����Uh,Q�AeW������r�#lJ����D y������gS�~��͐�`9*eM�.ȤԷ�V���E!�6De!/FW'�i=sO�*B���q*&ע�~���KT���L_�d�Up���ğ��q���׷�f�4��dV���q_1u�8�|އ�L���;�~�9�Rrt35��}Hz`^��ӄ�&�/P0�:!�T��%y$	��8ċ���.,�a۫ 1�7u�� ��]����u�V5H&GE���Mᾳ�J�f�)��/�C�M&������@(���!b��Ԗ�5�K �f/��fy��0��~y�0t#�_�L�A$���B�]M�ʪ�O������ٻ9W��2�M���v���S�����O�ۯ�>@O�j�&�qA)9�`P��e������D@%��I8�J�;0�����
�ΥT�V��o�Q~�/�}����R~�0���	���w�V��6ӤR�v'W����2J^���E���e�BbN��9Qcr�t�|�����J1�:�M�M"����bJ]R.� ��O�1���!rA8<�l����ɼ�����9����'�vN[��Tf�9�}Z� �g��o� #��B�ݕTB��*0�?ϟ�m H񲼙�r��ޣ�����o��h�`d�WZ������S��}�6���ڛD��������H�'�ut��9����=�?=tci�L�ې��u�Z�z��"*0������,݀���>Z�#E��\�3���.^#Uieʽ��ա-R״�B��m?�Z��hb�dє�t�/�=��7 t�ݒl����X`6ľ��T/OkI��7�+`��C��b��s5���"�\`�I��,�ȹ�k��'��`���������x�:�T� [}�IzEhPw�Y��r�6L����&+����>�6�O���}��I���~���:j��'W�-ܫd�D�ɣ��1u�G�)��֊��;"��|.�0eqd�%�(*;�E�$?k��Zi����Mtokc�%"hI.rg�AK�Q�Z��
.�0�:��9�hݒuޠ��o��kN48��-��v���*|��m��.�=C#J����.��S3�l�~��P�c��	S-�����n�^�;�il����ߍ�O��-1��6:V��<������H�#��\�-�3{�wh�����M��Gdҭ���-F�м�*��w�Uxe���ZGq�T�͌�d��P�+|�"��Zbš������m�Ĵ����N9�[��E�����_(�y��=DW����:�jy�]8;����8�1��*�tv���Da�G�)���)�-̸����0��y_���J ����~Uz'�XԳ��H�L�x�g�Q;h�j$���͏�h����O7>oAV`(��ok��O�}nEH�\E�K�-1�s<�rv-�	<�՘�n��'5���:o@Y/I.��`��4)���eӮ�� c�U���R��MT����hp�Y�x��b��};�ry0��0_�B���I���7*�_rO�"���8ғ 2�����?��)���Wȣ]��R�ц^`���K3v� ��8�I�өQ;����$��
{F�sV��z�ղ ��sl�TL
���w��!�m�S<�c��^��Fݾ7����3�7�9����{@�D��(�,��&S8j���E6�`�x�l�܁P�1r���1~W�"����ɑf�G�/ѵ_.M��𭡛����H�z�L���	{eR�f��i�\���d/X�y P����>��YA�Y��r����$,[̃�2+�0�D��aP���Vr셾Xc��㦐�T y�᧳aօY<�=�$������b�-j���\�}f�{�mx���e5��^���r�)�S�s��Ǎ .��i�ʡV��U?�\،["�x�^ZG��RR��`���9�N��u@��@�G�G�wI����nҿ�Y<�u�f��@M��t�.���Gb�C,r� 3�o�9��5�-^D�l��T���OҒ�p����>�>����o�t����ZE'
oG���I�����(Q�Kٳ�����i��+G��{%���K�:M��pJy!+q�^e�%&�o@!N�Ԛ~b�*���1N�W�{(��Lz�~ �{�jAť:��Aq�Z��[N	��s&�P��K����>���2`��fr&~4�t#�Z�-+h�3������y���>�}>�O�7�ij���c[�����~4�<�-�!;\t:>ӵ �8D�,�߮�^J�``�Ͼ�w{�ğ���Kd#�G˷|��7��3-���KC줟4�Gj�w#�.���c$����(k�>�$H���T`_tw//}�]o?5�f3il�Ww��w�ecyu�c$������a{"�q�2R��� ���잀W�)XFH�,��~\��Q��&ƔX�g��N�1D`���Eg-N��<�l@U��T&�&m ��Cp�3�MK�Q�7M�g�`��yO2��A7�Ƨ�An
;�y2�ԑ��ƒoFJ��e�!�ٗw�^(��G�K�~BCy�}M��3�DD��z�2t��"�l�������k.x�m���8�j3H�*�����Tz1X�_��)�zܝa��_��)�2��&��~㵯��1
��2%�����~����tGRyFt����ح���e�Hÿo����V�ʮ��í�O��d\˹��ӘA[j��o�=4���0�RZ��,���Z��W�O�U�T2�F�G1���Sb	�����tS�C��3���qʄ�6u�m��7�cN�E�x�im� ^�,���_�W��	��f�%k��$J�1ڎ�����d��V��I�9�A�� Yqwd��4 �F��J8>vVR��gi�f�n���g7��l��/Ά�*��p	����K 3䢦���%{�"���5����0~T����1��'o�Q.F�<��x�[!`ӫO$>��2�ar����S��5�t3f����SZ�v܇ud%>v��.?+�^sA�r�z��8i���#��%������He���Q-�5׸^�flA>D��'a��9%d�1݉d1�KBy!>qBNlJ�C��� �1O=8?[M�CM,HW͘`���,�v�D��Ẻe�e'ُ���S��D]�gx/�3�t�S��!�7�����p�%+6:��@TWKNe�\A;y\�C�gpXaa��= n��_q��Q]��%�7�>�z>�ZO]�3��!sȖ�����1T�I}D�U����[:���]�9�_E�b���������E(�'�������M��O�.��쒩�g�s�\9"�͡M����H�L��|��U��]�=�������;�����`�?��P�m�����½ף�_�݇�0��M�iLA���E�C�Q����V'ݷ4k�(�/��v ִ�ˬrm�;ˠ�&J(d��`v�H'�S�"���JB�΍�%���8X��x���v��ѡ\����%��h��;�}�И�t~"W�l��cg-���\��l�-O�X�@�f���Y�wy߯_�2���z�'g?��X�̛T}�W�2�+�k�!m*�n�fv�R����`�V(Vm�_��>�����z��y f�1}cF�>D��>���@���X�-�7%��.�A���R�(#�ءY	\�C�F�tX2 9��e|�zn56��R#������4QM::���ɺbR�r��INz��E6z.^�q&�v�tdo��U�'hV�d��-��9RWRZ��;ɞRÆl5�Ox�����}�xS�� �^eE��^�˼�jy�||URz>m���9[%C4/�V}ӼI���u��9l#�%�I�f#p�G7���͜�;�ߵ(vX��vl�!�~Ӄ1	�����WB�91�-ݷ�!M"�,n�9F��R��7�>�^GG��Q���1�b=I*v�p�H�к�n��x �M�~8���so�|S:ȸda���_�tq|�5u�=q���s��l��qC�:���%N:�@���j���kLK&�p�@%A�@OK��y3S��ޛ�^�n��ƫ�}a9���[��3�U�h*�Q�PP|��j'���AE"D)���es?+�Ρݪd�{6��(�v����ޠ\�J�	hK��e�V��z���t���/k��TC$=�o�Ұ��i�3��*d-k���]�-�R�,n����:7�U��0ҍ�^>mdU�u�߀z�e��yt ��¦����!
SZ,��n4HgU��]ߨ��(��:��u���X�3L5VQܰ�F�aq�.��3�ꢝE��|�޶P@ր�tܾ+	|��*�#=�_�j�'A��p@�����Ֆ6Z�SM�)��)B î%�^8 nz��W�L������Q�)�W��C!�N)^+BM��������Ru퇕��26��^5䊀|5�I͋ �I�P���"��k#���'�f\~J�I:��-]��3l��yO����N�0�Hf��r	���y�{;4w�#�G�t(z��s�Hy-�iK�I���9���ϩ���%�rsT��l�H�*��'e�T�1���^"�¥�� ��m�Yqꡀ�����׭�YMR�}����2��M�o�YiP�T�$��N@�����&� 2�� �3˚I»ԙ�O^^c�����>;�Ia����6Y_��;Բ�ݴl�6�1y׫G���F>Ȼ�g���B��CŁ=_��O��^�~<V|,���O��WySЀ&��p�q%Xj��JP$������8�*�z�,�ָX����n����7ؘp7r'����� ��j��k���?�]�[��o�e��&hP�*�ыH�� ɍ�:Ta��Q��������:��qe���Z��Z*{���da���߈�	I�߀_f�� ����~��T"�Y��vmE�ii�Y5H��7�I4��k^�HNU��HŃ���؁��35�{��v�>�ET`{yh+��ayI(�����>��ko���>4�GL1�4OIT�?-�ɗ�;SЕ��{0t|﷢	�A��!�e��gz����X���Q�B�^Lq�Y�0|eO�ԣ�	�̑�^�*���T	V�Kȴ�(�h|���;�(J,&���F����>Wg˙�|$���a���>�9�{~�J����9zP�Y䮬:|bky>�wRsד�4��,7���_���A*t�vL�V�NU�����3�9u�(2�R�kg�5�ӻ����:��}���3s(�b��$�
�v�o���Y$��`m>��t��=^�P�2�$*R��߶�dR�]&�w�������&��?ϛ��}ׇ��x�Q�@�!��5�wO R0�l��b6I�tis��ixQ{A�ݺd��UbT8�Z��j�(|�a/m�:)�h��m ѱ}��������W�0-XpC��	��^˵!9�j�l�U�?�j��B����LV7W�D��ý	���.	������a��U��ϨY��G��&h҈Ʒ2������\��iϏ�d<a;��g��]�
GB|r�v�e ֗ޔЛ��T�:)Tʝú�'7�hf�(�ʔ�KY23h�~��5?�Q��<��S��k���3�۝�f�G]`���U2�b�6s}�_�$�W2"��4�HLfJ2G�b�.����^��|�H��0g�B�?	.��*�������o���hw��
3㾁P�<xyӪV��%�>�h�7���\PpGؿ��u�:զ\�!�`�[yE����ᙾ :�w�m<�rg�ɀ�=ǆ�Q̀>��y����N&$䓮`�[nx�ày��;6�v�S]2��i��[��{�o�����GDS���*:7S�0���9Uv�4��uB�*|�:1G
sH��>�:��X�ꩿ�(��������I!��������N�ۖY�n3���^�����
�ɍ}�A4��Wm|�_P�8rۛF�%��⌽�hd��L͞��Q���]�4��l�Uۈ�<;�{e�=P���-����!/X�ث�#���w^X��h���{�7�Fo�V�e�v�7O�W^rL�%Rڪ� )�u�N�
;��Q�O���5D^�wʾhj���=��� �Ǝ�H���%�Zel�*
qck^��8�Դ�33�m�h�������X���]J�䃧��f$��1�4Eft�d_��(�� �.  �ŵ�ƀo>O�YF%�h�+܄����2Só��]�E��\�'��L��d�+��mˀ�
���D��KfqL
 ��.�7J��(o��X?B4qJ��a���q�Ѽדͺ�g`��q���[��Ձ��gM��mCXHIK-t��ccy)�н"��\��\S=���P;��6EB��o��	`f�quM��h1_U�pآ@����A��#��V|�Q� �_M�pO�G|�yjƍ&�<����I��o�6����L��'��`��X	C-4��E4��FU���.��9�xa�Q�c�K���(c�T��7_n)�*ص�o!��b2^��m�s�o�vG���k?�n̪���Bq!�g�_X�5��V0-���.ȯ7J��x(�2�6l	�u��?7\�,�|��[��~;�_qU&�F���MrZ�:�amw�J�ƈu�4w��y7~���/8Au";NG�a�eO� `�ȱ7�������Usl�ƥ��<�V�?{"�ؾbd��I.[�]��1o+��GrkeCD�	8�q��f�@� ���BUY'c��~`�s���V q@��0)����$��,�_�����4
pP39,����}�d�T~'42)#wC��4�S=-c� �����j����ث��?��F�j4o����ʨz1��9V����P)h5˽(�8�qʐ���[�
���E��7{�T�яW�j�(N�O�q����˦=��P����rI_�����`�:�O>2K�#�������^� ^�$Q�F�c��/�NQ��M6�\,�"����7B��?��|y�g4B� ��$�i?��>��V��c��ʇ�|��%�K��]��7�����(Ҳa��v��_5u�H�Y������馫V��^�f���޴�+����/^���XN�Y϶��1/=���2�p����s>�ʛ�B�<�H�p�:���<>�̠l��c� O�F�>��+��P��k������P��3���/L�(r�<�{TҠ=�zf�9�����?)J8*������	|{���z�*�� �Zˎ[L��գ��_n����r��o	�oZ�^+�e�D�Ϊ&7���|��_��©��]Ɍ��ԩ!�*{���{�:�QH^��9��'ťe��_�I�?����k���K�.��,����w�&�_�^�j�Q��E���.���9�j<�Ny�� G��Q[-��ퟦRD����9��vp�Owg���nRj���H����Ŕ�F
��pgV�0ţ%�߄�	p�v��f�7!sƐ�(.��2m�������ጬ��Z$=���5�KH��h�}��:_��dm�
r���1�EY�Smvd��J7t)���X������}�}4c��'d����{��p���~����ܧI��=�?��u�.uO��3�:ٗ��O0��'ͬB��_W6Ԑ�r���W�i�吐��&ğ�cY�	�}G/gk������Ӡ|{����A��˵�,iG1f���k��v�:q�Җ��^���Ư)2BP�H3����{14�rP�=�%���\b��Z*!�u�N5OM���-���7i�^Cә�{z��\l4���6��";e�>a�����kie.��>���c<-�8�6�
�"Ъ�d��X,�"��g�C_��փ:��h�aZm2���~�;���uL|ʎtFo����x�.�xoKZ����,[^��g
nm��AJ��H��.�o5�%�=)t�I�eHUIn0�U���
ʏ5,L�2��x�^jJ^]=���1����'���?&,1"��l`�C}�om���A@�:S	�/P�X��-;����|�,6V��5�.h������J!@܂u��K气�J�`��ƾ3�3y�_ؤLp�1TKE����?)��j�i��⸘�x{�SՍMJ$��G�2mY���,W�a\j�^��(:���FJwC��V(gd�p�l���� �6��`��-�ō��&�V��&�Qy_�GH�J�4���Wi��fD"�(f�����,m6�����3u*C�,�F1��l���3dp)Z�zzBI
0��]_�/������l
��5__ni7n�g�\����)G��MWHOW\����a�
�	�Va#U�!��(J�K7M��^4�6	8�I3�����.�0�w��Ufɢ�ML�{�n�z��-��F!Z=�%�z������;�[0})�Rn�-M�ڏ��!��Q��zc�z�:�X�V�y�ܱ��[��a`W
����z�_ƹ���J�6�mŘ��&& 8,S�e�aC�I� ^��^�6P�>��W7���)�-3�q�	wc�k��N���T�qR�eJ��e���+C�m�e�<�/�C3��D�!���^��Dm����K�F��tw��EL�XٮCY�
+�5��o�1��u��4|�S�H��BՄ�(��.�1��[��0�`�߁���"�M�1�ef����ژ�mz"��H�42Qh�WϜF�6���m_K���>*����
���1�t�R,�z�X���YW	[�HP�)��M!ă��9�{�y<_}Z��.
q�Ԛ�Bһ�5x!ד:9;qXx���3�Qx'4�b����z���CI�rΨN�#K�Ɂ�ϟL�aH쐟`� W�����"�4_� �Y��O;���υ�Z:���ܢ�^otoU�9r�=��[�z]��@������|_� ���2H�r�쮷�՜:q{t���64#�XB�O'���Qsl���KI�t�X>=���z��@���3zqC��Gj������!O��ܔdے�Tzi�D��iRȰ�{=��2���w� C���r_~��`����Yb��]� f��tn�i��_�XVg_� �]zGܺ����@�G^ő	6�*d؉��EJ�=�f*���' �#��<И�Y���ҟ����OndŻ�C�z��||\��.,�v�������x!VS����:��Y��&FT(%�7 �R88j��?�����������Ld9�mI2��=�}������[N
en��>{ɈNE�}/[�>���#��=N����n�����i�L4\X":R2{P~�&g\/j��Ӣ���eQ	d�	G�?�R�jNP��2������AHN6�RM2���:��&�8��l��m8+}|mw*��N�c��1'��UON�u�]�Y�ea�H�{��qe�M�������'��q�b*NY���M�Xy�o!�ݕD��芹o�T���L�a���O�}OksB��[���dvc�e�]�8��*o�.�y���$q�nS�+���a���Gx�g�|��D){E�Dh��l�].ֻ���^zj�*�F{ο~9�E�6�=�C�lr�:�	r홶H"�q�gYp1,4��Ѻ��Mc�%s�Q)����[����t�T��]���xz�	WЅª��:l�2�����Ww��,�NV�r4g�!�����s�^ٵ�[5���jzJge?U� �ӿ�	IӏAw�Q�7���'�}�[;��ŀ'F|�IK���]F`��{�à� *���A�sz���?R�9Y����K�V� �Cū��O�dAP�؛����(�r������!����T7Vb ��)\���X�
��#x���⎡Ax�s�j��z��*j䟾��4<�G$�x��8�A0e:� ����U^���T'2�"_ �ԣ�2��i��z�,��C�3� =�Y0�ԌM���)1W�[����}e�0�O�Is���U�[)�&�/���*��
�DY_���F ��b!�����})��i���T��&K y���~|.��/�R��؂�Vs�&~2_�_�&ӡ�v���$c�KXg�� �p��t�t��������*�t!���5�ש����(54�Ʋq(��I��f�rn���p4"� \\k"~C����{L�|�U�w�P�zB��3d��p)S/(:�X�Ґq-?����nn��J��qƩ��|�0c���0����r8�#t
�
{0�y�B!v�&�S��ʇ*sC���N~�3.�sA1�;6�3�^� �!Ǔd�� +f"N F8cTI&�Ŋ�?{bo6�V۫��@?hD�6��nƶ�oz��T��N��	�W��n�k 1Z�?)Ɔ.�I1&���,
xn��
��(ȿ�a��_�����^C�Gvb:D���ֺ��_��rg�ز���>�� J��������lI-�� �9����vLg�;������i�6���3���T��2ژ�"��E�M1�uL�|��ʀ��t�e�;񈇂���5�t�_T���͙rld/���
�e��@w8':S�ޞ��l|�V:4#�z9�!yhz*��E	̠Ř��!�iT��,�t3~�Jl0�S�ٜJ�Xo�i؆��ޓ%.œ�i��_�s��&��2+ςc� _���,�19�8	kVO̩v�~o+�:�[p^��=G�B�N; ���F�l_���,��q��d������_����W �(��$U#�9#�Jf��}�M��:��R�k� �z��0t����.���8����±M�h�Qxs�_�qg�6��Q�d|�Pw�̖h:]Ͳ���� }�A�o�Y{��j"�&|@��&�'�����:(m��q;-,��/�cOv�����B����K���P��RN�\����=���ݱ��"2�R�^*H@�祅���z�7�pS��5��(gB��C��m}2	w��2�j���nX���] #\��@�ËҊ�g�2Í��� "ٌ�RTj�N`D�بK0�ނZ�g���'(��#�����^l��r�U�{g�J>C���+kE`��v6�$��]e���o��(l1RN�.0s�'���E�Q�2T��]J���M��p��Χ�W�F��� �� ��3=���n��X
p{+-� XҲ?*~�flv��&ȝ�}���=�ʫ>r�O��4@t�|s���8s5�s�Y��5&������4h�u`���Q�����]g�r������\l��S���5������)`����`��N�A� g_$c�K2���"\�R�-��}��d~�"��2���' YY��O5��_L�#�{4��=�RO羕�� bm�#�P��|ɩ���WR�?���]��F��L��r��ʞ�4��n����f�X_e#�>���>�l�d+���rH�g�rњ{`��X�W�n}��rx��)��c���|��y��yr;D�Ԣ��@��8dH{��^�OS3˕M��BЏ��)+���G�"K	"Q�&��Mݝ���R�ު�� ��,A�9��03DN�[�_T�D��Y�V�����*Y��^�)v&��j%q�r��:�Bb�jݫKN���y�;J*��]��lC��5w'�!�NX���hGq�^e��Ŏ��d�������>���8wcI�� �axF
k~:�(y�o�>�Tӊ���f���w���Rv��t��S���F3�i�����K֔��]0���j�����0�#n�[)����bH���W���2�Q��"0�$\�_7���E���}�v�<��o!�i���,���'x\�݃Uǿ�6���M&���1���&���N���(A���V45H���b�3��M ���@aM�{ �fXb����V�Qn�=υzt�Q���M�89�3w��D�V���TJ������%�>H4�eE�+1�wޝ ۊLLhǸÓx��X�4侦������ۦy(o3����=�F��F�A��΀:^ͽ��r�[xa�w k��z� �	��"�~�4��@�jF/�ޣ ��<��i~�<ida3�Eq��t�`��6e��2vt��+
3�8�8��P��`U�ɁN
l��)M|A1h5.�3�!<���7��ωC�!�1�C�@�n�84���#�W���`M!d���,�(	l�aK]q��G�ݐ�
�A����țb�68�l�j�f4Z�g�sVU!Nn�I1k
M��N�:4 Qg�d�$�X�2b�<�(xhZ⋲��-.�a����G���_��y����`�%[�0t��qnv�������&���ʕ��'ƅ%	�f���)R!jH�a���:���%�ln�j�/Rb�>b�erq4����%,�M�C�'�f��$�j���P�,��o����)y{�#]����Eh��zl�/��]�+���[qќXaqeO��/��uO7O�� E/�Y���!�5�&��T�g��������ƊF��<�f���A����!�k=���xR�ݒ0y�t�ZX���=�]��+P0���)<u���٬�q��;���%�*ER�RWy�]:�4�?n"���]�=�g6%�mr�
�f�S,u�T�@2k�
��	�IF\<�!u�	��cF�c�]Jh�*��{�G��Q?�Z�T^�YxR�hV�F�B�ʨ�~3�s%��s�}J�dB���' 
Ð��E��+Iz7�)c[{!%���;��i��~��K�;�LQ���������|���n�#�<��X꽈���N�'�-A�C�ȯ}9Iq(QO�t�ja�4�e��I�y�f�;�A޹�G�� � ��]]Ż�~~S&�oW�J��Z��0�z^hk�%�4��j5���	k�o[F,T�-��;�쭤��_�[�'Ů�og�y��+�ʬ�(����W��k�BV�w=��]
R�<�w�%�u�(�����zE��>:��K��\�%F[�3���:�3x��m^?��"MHxfao��H�U�ז˷��dBi�H�e�?"�@Qb �TJ;2&m�����T.�e�¥q+JZx������}2�̈́����{L�����ǘ����c$��������A�$��Z	�����m��9h<�)�k�J:/˥�7��|Y�5�&�&������t[����RPI��r2����J���"�G��v	���/ި���G6��O��:�8~j�ú�y�t�c���cGC��]x��z)uַ��e�}��L�:�WnФk�TS&oŮsf���Ә)�.d�)r�?(M�*p��ݟ��>���<;h�{�ɾ=�0
���n3���q��hH�N�3d���&����V}�Z��4�Q���*7yi�O�i5^�_����V��),=�"�C���u���jB��{����nZx����7�,���o�U���!�t&�Mg�F���"�n�}�p�t��Ie�� B:�x����0�J��ym�~���4�\��I�����L�x�S��!�3�{�r%������n�0HG���=�a��i�.�Z0���'9�C��Y* 6��P8U�2�n��Y�l�N��ً�D����̄4� �x��������r�G��)�����PE�����@ڞ����*_X�G�)o0�^<�ms0&��|MF���ƑӺ���:�}�M�=����Z7��Mo���?�S�F-���Iٯ�U���|�(yd��\�?U��MUh�K��`��`���C��|2e������P�4b*\?#���TF���+-.�m���af`�x`^�s��������(�t�Q�*39	��{�BM�N'j�����������Wv5�VL�8��*O��9C@�?S��C��s��R)�V��g<i�Av0Q�Z�}�R�\6�껺_F|l�Nm��_	q빾��@���_�:�@ ��%�bt�]��`΍�ZdG��?�kT�]�;��5E�ͧ饑��h�bz#�!��u�6�'~�����48��4����;w-du�gx�
2[���ƥn6F}��e��GӀ��5�t�T��M���x�Q��B���>:��<�Z�G������|o����v���q�xJ�ٚF"�"�"S����b�SD�n��QiC��
*�9s�6Ky�����V;�+q��W��q6w�D=%�U�D/�&�mX��X&M�`�t)�Nv����U�q���Z��;g�.q,����K�i���yj�ź�D���&AWnI/��R�"�F RJC[�o�$��s�F�( I���4�E�ݶ�����x�c��눖�U�T��E"s��85楸k����G����s��X��|n]�_-)�>���T�ܓ�e��*��Z�NO���y�.�mg�">�8���7�!��c]�wD�b�lqr����S�i�=����5�}D]��Oh���*�3��AGN;�B{ln{ǆ!�r�L��T����!�C�Jv��CSp8�Waː�?�r�&��K#a�~!-�wA�ֺ�6)����{:j	�Y��'�&��F�=�PH��/]}a֗ {ךF@�W0̲�s����e4�|��d��ɨ��u��u����p�����uq0�N�	>T��5����ZNE��������~Q��~���]�)���T!�G��v����j4p�����ܻ)�j��x5���RU����P����1K���,I��k����'
�7C����6�]ۨ�J,���g�>�,L�Ofe� �?��Sa^�m%��=m�.Zߍ�h1��n�Q�;)��P�~���/�NL�����q$^�s=���ᄓG����^w��Z���a,�:�����P��sw9A�� �u�-?��B|F���w:��OѹJ'�����/�� Y�:���bn�]�<��<~~]ni�I�Pvb_��W��,���:=|'Ċ$HݤME������^y�Im(SU���<#G`�|��KKϦ�px$�C<�i��*����AXj���cwaZ��fy��el�<9��nI����d��*e
�'MM:6�6�zBL&����X��d�������U������Q��V�KLo�2�����0�Y�]��� ��ĹD�&ݤ���6�r�z��"с��Lp.���aZ��H�i,��(�Ii����}��?�i�?ɽ��rq�^祥Ŗ(�8G��ǖ��K��1-��ijc\���z+k3M<I��wԭ�4�#���Z�ك�U���J�?�)�c�����4l{j[
��'Bܫ�9k$��4%�sI������
.7����K���� ���N��������r������vϠ*E)�A޳ﲘ��
��cۂ��.d�la+똴�U����Z�?�&��4U�]Z���ᚤP�to�^'e��
|���n4=o=܏bm��~���G+!Cj8xr)�f�;4.�DI@*kZQ�e��c�@�~2���Vc��ρ�[MB/��TG�Y�-s�n��l
d�v��&��1��BEaU~6��Q{<��h�+���c-β��z-�k�M��!�y����pL����R��ԯ�!H[�����TAw�ԃ+���ګ�ǮC�`�[tj[�p	M%J1�Cy�E�?On�fC����P3�X����˩�J֋�R�,�B�m(��D�4�������⺊S�1Uؖ��~��պM��@W���X=��aBݖd
�����l����QHz�1��Ӷ�u8S_�]K���V��%��,�S��X9+���L�67��}eTxӼ-��������}�<�W��1��{��'`�5}#9 @����^-\'��ɺ��7M�_���[a�gLz�:�Cjp�LfuEP[%�7w��&7^��(���!2��?02���ʼY����W���f����
�m�>��լ��,�����Q-72o�Ǟ��,(�/3,���aÒN�9��E���sa4m�dy3Y�tF������S�}���	���Rdçx���:�j�c�M0����4S�(э��~��Iqؒ�G�/�a"%�(�T�r�,�����,�V�D����2���I뻤F*#��[-�b�M�oB=�}N+��L朔VY7�dv�΀���ۜ&_��i����?^���
��AZ9������^��"��ќJ�|m�m�j2m��Z'W��Xu�h��a-y9��[r����.��_&��X"�!��"�qy��%��I|��94 ��̈́J4	�B���(ʚֿߘIqIJЕб��I�͑	�b���yx��b2�@]�y���S�0o���4�Gug���*��I��Q�F�碠���R���ɏ?w�6Ŏ���C�����A�̂�潭��$7�w��]�"&18b��'���/Ѣ�O@-��8�mKЫ����f�/�	*��:��'�o�,3�kr�|^�����˙ؗV>�=���R�p�����є��F~��6O���(�WR�g�俯��Q ��u�tNLĆbyEN��e;�|h�����)%��$��<	�J)���.��<I|�m&�+Ş���* L�TS��W+�^C�Z�k?��*�<�!|����3J�@�%��8�7�l8��Bd�k�ٱ�c�� �( ��2��
6��ˣ��T���ҤH��5(�˨_;e��.����og٣�s�R\� ��9�����F��������b�:��V]������hpɾ � �����67ԉO��)������?F����1�7����'Odû[f��O��Gg�HT#����:�7�g~�*~�����Ej�u�y����^��a�0*�7WF�*�����1W��m�����?F��e��.��m��۵~����7���w��#�;�Fʳi�p-�J��(�{����'}�! �>�S�ӿ?�LF�eF��D���7dR���%��F�����őV֝
��d_.�ɫDJe��J\��s�i�֎I{V��@�6Q����:,ih��'���}��T��xL��{����v�T�ky^���gn�A0ʅ�U����ܲ��P��Nr��1�����_�n� ����{��K�� ���}P.(�Y4�r�5Su�Z��/I.��M�����`W�4aa9���1���Ա�(Z������M����휈U?}����� ���/�����3-�$_[�\�G��$�0���/`�e�K�����ϵO����ݩ�N@�˹�!���"���7���uw\�̡V�����Y�� �6vW�zG�������~��������h�N�}��]�;�PT񑜰u _��
���x) ��o��r�+E��@#��/�X����q�Ѿ���n�����k~� ��X�VY$�J�Z ����^�|P��Pcތ���s ��H�NNX�X�Z�U%����_�
�v?ПXm�8��q#G�d��l��(�k��u�J���`Rҋ�I�=�vGٽ�Z����O��U�o�|�ؤ9�0��o���K�}6#ud�_�a;}`c'��u͔=��t)��~��p:.��;�&��l�%� mR*�=ƃ�&��u��2'�S����qtF�]WW������S��2������$8O�;��CB�
:�k_�x���K��9�c�, mn��q�X�"X�-��E�͛F����U%��*��8^�۶hՃ��yT^��8(|#&���xX��k�����k��kG�<��.m��VMPY��J��o}J��������h'L�m��::��Aa�0�L@�~:�
q��o�s)bh��}o#�lq�hjOy�����a��$�V|UfD	��a1n�<�����,������� ����9 ��Q"��p�
1=�����b�8���"�vt��َ�C�`Hcq�ʴ+e�!b&��%7hf�&Y����,�����j+��>�?�_�N��5ܦ������di�},+�C3��������3�~W\eV�)Y���E���i����_ s�wQ��>��|ŝ�t��"ֱu�yNoJ�PT�D�.�w�h[�H��L�<?x@aK��])H���mZ���3�l�mX�Q@��<�Lb���w���`�<�*�w��Ѡ�\
�u5j�$�� �+!��NTr#���}TQ�ٳ�bY��:":�x���B�[�[�z�x����n���_K�5!�.�n|ɽ�BV�0��@�<O5�'�Ȅ�Ɉ�߱#0���i�r 	ˋ`"���a��*��H�쩔�)>�A��@k�P�9N��2e�p�6h�z���{�!v���Sb�cs����|��|a{j��$�{fƳ�6z�NG�*�M(kW�p3��+V1�<�XT��=v�5<�h��\0>,;��2	P�Pݰ��g5��
ٛ�'�͝\/��avJ����vs����(Qp�Ϙ�K{K��
�W�k�@$ �n�_Qz'���Ļ�o��7�d�;�,��:|�P����Qd��#�myZ���w�G%)�E��/��S�[��Y�Sy�����|�77���Y�قsf+�q���'��l����hz{.*��~+/���r�� Lr�O/T��es�ߧ��{�!�;o�o�(��j��7lV��Iao��n�&��FF�:v�T�48ű7�e�"���S���B��)2�C̰>��k��9 BnnVB7�:Ǒ��t\E*qa��d�8���[r���&C���7E�qhɟ��,�^F�>�5!%�1���VdB
��x_�Zn��z[��k�o4�w4�Ǻ2_�5j�O�;8��=#u�"�\���f[k792�7��(�fQ�P��j�d�s�3~X�i��r$K2B��J�̥"��r�~׳\$3�˂g�@X�/l��2%��A-k�n*�����YG�B&��e��+kp <聯�u]
w贺�&yw裦�m�R�So֫ٲ��|迼n��n�2��թ�
Gs�*.FF��u�7|E��G��m��$ZуZq�p;�~+���t�k�Ƴ:ڨzLKy�Ib�ן|� ��3�ɲ.ș?Gf�PW��:Z�8q �@��(�/-2B]�=�1�K���� �
�^鞸�[.�'xR-*W��>�����(��\�?)�1Gj�́2�?Z���^}�&^m����ՠv1�d�=H|���s�zQ@ԉ��_$u��\-5�nB��71�,abR���ԧF|ZR��\��<Dsx%Mڀ�x��߃�ތ�_ߪ����J�.��.g�J�p	�m���R�{d�ˡ��@�16B ", �aX� ��L0�P��$}飡�M��?�#K�v����5����@|�H�����!�"�����FkR�X|�PY��&+q-r�Y�>�l���(��q�L6�\{��u�t��AlϬiA��1�^�f7�c5�r��2���������+��J��)p�~��y�)X��9�������玙X�NH�a^��j�Q�7+d�x�௢f2ۤ`+ݐ�ۜ	���`m��|�3.�����%a(�)Xj�w\z�R�{�kG��4���O����h���_�5m�3hi�)x�O��cO���s���6�
$����|[!�*����d;f_Y��L$:"Pi����X� GF/�T$�-�_n�M���TS�U�i���C/82�4Р��

d\���}L���5� }��K8@Y�ɋ��э�W�xߡ�4|7�/rB��|�XJON����/�Z�|�6�&�A��u4�_��8�g��ю�g��`���D61�F�;F��Id�`�����4�6	�/�-����
��7Τ��oq� �I������i��5���3Z�O�4�I�ެr�(�L�'`Qޏ��Q� �|p��Ե�y_�Ff�.͝��������<@�هӱX?>�Q�b~�STLG�_ �*�Dy,��������,��sZ���ԘÄ�졨͙	�y�O骼��sn-S���B�:�Ϯ"��:��
~�ڱ��g����w�<4��Z����<���J�PT�QB�HFC�\�����2�_r�q�D_���{����3�E��ӹ����r�ɲ�s���C0��/�o�lB���j�b��8�s�[��$<(`n2P/Ҍ,1l�+�<ޱC�S5�3��)�Z��i:��r�~��{Ilk�~�j�a"���3%eߨ׫{K�e����6����	�� �4uh�g�:�D��TW2QO0zm,���)#�}��l@N�[��gC0jF"��M�+��2�·pD��
Đ�����9w?MU�oՎF5I�5��r�k��m�� 
�t���Ғ�o^�O��@�l��E�8t��|w� ?�#7�0Q���j� ��~&Cd/�*��s�w4����ma��=\�F����ᖬw���P��,�����'�_�PJ�(ԵƩޮ3a���q�%6�׎�O�1�u�cj�ogTcY-�{��R�Z���f]v��������e�=��{���yiK_�Q��_�0(s}E��Y|�P�3k����^���\5gM�vӓ`��c��=2���7=��~�4	�[L�E�>~���Jͽ��zD.QY`V���@? ^k>�;�(Mg�QRdm��ܽLB���GN�x�A���L8�`4ZWTIoGSB�SS}S&����y���/���#}Qy�(��e6ò����83��`#��ک��z�Әƪ�������.�
����bo��qȹ����~���]r���	��,ڟ�,�0=jF8|�t�1�P��(pIu��J膦O�e
6��!����<���M̃�l}Zj�~��=�H����.�	-��v�����*�@�,�
~�j�x���k�?�z��N���`�_��%�$$\�o{"E�=�����]cA5����_m�ܙ�R�i!x	��FXҾ��yʆ�i�5�L/ރ����Z����A�BOFM�4�Y{'q�/������j�p��r�]�2�^��"һ��I��ncT1�����V�Mzh�����}�0���g�A��m�8�W03X�կ\����iԀ@���K���:��!��6
?bx�k�;F�E��,��g�T3���J�9�=�8^?/����y�����N���m��lɖC2(j��2��~��*��&InD�zt�>Jt�a^��Un����鵤TC��寰�A1�56����<
5��O�Zg:d/��s�j��|k��0��#d/!�_eF�wrjW�*!�8*�������J+�!\!Yٍ�.�~Q>�
K�`8�'�;��
Fm���Б��G%uC~�2@�)8��%y��{+澪��V~��h}?h���VI�V+Z���E pUaW4Sg�ĵ��H$�����jj�L����:�ӥN]hh��a�F!�'\=G��3�����3�{���:�U�����g���fK=rn@[�� g�#���syK�J;Н��E�_��1+���kZ��A[����	�Ш�tn�%*7q���7� �y����V[ƽ`I�Xs�g*�>y�8��gjټ%{%��6�B�P�d�L(��1�l���t�߽�S;9���i����3�5�J�����U�zCO)�����I1�P��G���x��p�.���Y9w!{M�6s�I�ʶ��#�&�4"ɀ"�R�U!/��Ő>,�崟O=1�Vz�rZ��eC�b�LX6Q���
HH��^�mB��;(�rd��T�]~=������%��G��[��'�^:�� e\����9E"8N�棍a�M���.f4�Ӌcb���m�f=�I}̦�G�}�{Li�i�����nd~��+u�rۆ���^�詧"��p:�(��o�|U�_b���\��-�V���7¯fx�O� �Kw�!t�I�$���m��?(��d,�#��O�
/mw����.'��?f��3|Q�n��7�^��]�oP��b���ѫ�C�� <�8�����*8uf�U�CJ��0����O��F��p6�%#�&Ù��R�)�B4�~S
�|�r���jʔ�&�Fm��&��5(@�^��*$�v�j��ߨ"(���M��J���ʯ����R��+=��(�� ��lS7@����ԍ���O�����H3ee���=nu��x�v��a8v�������\NYF�Y#$�m$�9d��\*�|P��DT�Вc�#��6���2�j��Sxѹ���=����(�o�Ҵ0�MBy�W#{�r3n39�c3!��� 1-溮�+�w��xc�|������_�:Zw)�֜&=���>$L���	��j�T�����mGx���������+��He�~�ɫU̵�2Т˪���1���(^��kV$�;;��	��b�\�QQ�s���.<#�#_��M���L�f��<R�~�P?��k	��T�sW�&��H=2]��Hrǻ�b��2Y���B\0H'��9��DA���Io�G�'F��"���i��0# ��{��w��3
����Y��\��(km���v�F&��89���AO��B3�� �F���������,$ce[�ђ�`�kЕb�8I��-��~Ԭ�{��x���8���n��Fcq��X�h�#���ҩ��{�i�U��\vu��Q�<�yKA��i3�P@. ����0����'��1h�f�*�L/�|<A��Q�D /�̃����,����j_a�����{P�{���~��v�������m91�yAT	����R�������1�y�������P�흁��}Q������T$��(O$��dC�v�9P^|kE�2��-��/� >b�<E<��5�X�������'�%�J���o�i�έ�>�>��S��#= ��h�n���}�n���N_�_��v3��?c�μD\� q�;�x~sI|P��T���'�E�p���`���I`}���k:��;�d�i�8��T�̹x,��H\>��Ϭ��������L
����V��*��u�0�]gXo���fs/o@�����o��f��БT�}�؉D�s�1T��bfy�DڲI��ڡ�������k���r�<��f���������(�>?��ŉ��!����p>���H=��i��KX��|�U��Sh(�'(zO��>����"=	*��1��!wV�L��JH�J}孪V^o<��>�0���~����	�gdez����';Pj�~��J1/Q�9���AB�;�q�����-�l���j/�
a��Iwi'U��] �54z�g��.��X�`�|��s�[���~JXN���m�*���Xk3�JweA�w�Aȕ���D���*����M?zڨe��EٚQ�j� �~ХR��
X���-��-x�	G���Ȉ�-�M�zw�5�0|}i��CL`�2���Y]�{��!��
"u&߄�3x�@���і�� � �ֆ���bؐ�,�7G�aLw[�@��h��4�X�����A٢]k��E��~U�i����{�ZZC�Jt�qO�Q4W*�?�vL���/H2AYYgN���UǦN���އjo�&s:�H=(@C*U��Th����m��I��!��,ـ�ѯmv1'�Б)�5�#�g5������ˬʵd�C��
4�Q��0��!P6{�.8Ɋ�L���爃�Gn~�F�,3��BO�2f椊Dm�虋l�t���˲-����g�v��M�rJJ�ܥ�>���xGRɈ�Ds�1�}Se�g^�b�>i�鷠��(���)y;jII��e�k��:9}�8_����N��"D&Z��$�Lp���G���ԗd�3�}^$~��E�� ���"�1DvL���B܏r`��LP�@(~����2\Co��%���G3Gy3u��]]c~��w�|UIl����o�`Cv˙A�}c��,��s��j\+/��x-�\�2oW�w�c\�����\�T�2~���s�]�fu���K���~�13dOBƐ��������A���!;x,�DRi�%�������_4CJ���'/Gzķ��='X���#�.���y��l���+Ӆ�z×��#��ߟ��(���p);g���R���..
�[��f4�-�'s'��L� �xvГ�`d�*"�Q4
��{T�����GrvW�U���;ER�e�o,J!�^C�4I�e�6J[�g�2��#,6��M�Q��mϣ�D�6�q�Bp�	�waT�Ѭn椔C��&�*�*�˂�[����q}��aC.�9iZ��K��kV($u9���C{�^9-�^غv#)6��V������JFf�8|��k�΋�р�|Їe�ߑ���e1���ĕb4������H���D�^V�A�XV���l
�x���ۚ�V 6�b�;9jb��G��U�������<�KA]�t�����CW]�V�����5+��ʎ\���v�����2�u�3B�5�,6�_��_��9�����jhu�dY:@Aյ��¼K�,��ZE���ٛ�}AGm�<v+,�z��ܽ���WC?v��+Rw_�V�\��"��-���^f9�Xލ��EF!�h���9[a�x������+�ɹ���{�S��vuL���r̞�G]�@�8�y��~]X�b�2��ߪoB��׌ەS�1��/�OC~�<%�q.ݰ{�|�L~U�Iq/�NVA�;��0V�mʚŷxM:�ؒ)���=�0��c����S�X6k6�ް�S�J+H@�g��Y

>��/N�'<t���Eh�Uf ��zܠL���/{�L�p�fFg�4���=��5�tC\��K;;��I����9�&R��~�=#�y�3��Xz5z�3�
N�.�}�b1y �kqX�H:�z��SU��f�[��Ag�h�-2E(�|x�k����~�AZ?�i�K�q�E���0��wz�!�/*P��:_��o�I����DwM`%��KP8π4�����72�$.Y�qw�W��@��{Q���LHNvc�&��2�^��y��cw������x��#��z{�Ȩ�Z��4�Sӥ®kc�Z3�. �v���Po�k�_�ِ�"F%(D\��D��8s]�V�?���^�ׅ_�Ⱥk��[�s\+���%C���˿R�� �+�(��i[4���k����� ���E6�u�[s8��s���>�U`��Z�h��N��U��Z����Y������3ȉ���L�0�Ja�������1e�5�W��Tz�Hk%��Vr��6OTZ�P�/�vC��"�s�-e]������E�υЂ�7	ge��m��V:�"�8�<�f��^�5��n�Q�u�^=ۥ���-�Ie�|p�%�A���F�3�Pĩ���5�>
u!�4l��.&+E�][��7u�%�<mr6`��!~���5���k����'��"a@(���е+�rifXt�2��l+�-��s�l��χ�ߧ�bj6F}��rLԿ0�7jQJoׯ>�PK�.�r�Ӻ Q�)�C�DEdY�\�MT:*�CJ�=�?а{�?Srf��J��#E"������Vb�|�c
�D�g�Zj�z�h������^�$_��p8��*����4 ����.��`)՘�T�e��9c=��Ȩ�6��X!����t�t�8ܤ*$VQ�U��6)��g���;D�K�3����h�|�N��e�j��(�W�^eLg���j�ɒ�?>��O���9o���f��k����sĕǶ��oqArb�m���l		�U8��_�$��Wc�3 E,�B\[�J�ʤ�l���Z7|��"BUc������1����4��s�����K#|b$!Z+�DUB:nsF$a�d*�xct�1�F��!$ѣ��k=CF[O�o8�좈|�N��_��`��,Y`V��9m��+��`�ş(Oi1�ȫ�}n�/S��y��ó���+���ot���}J���� L�2���$����d�6N@S��wV�4$��b�"�G&���!Pg�'\r���t6��(X��� u�����%��p� �|B���Ңa�s&�p$��=s&�	��u>pg�A�۝:S�<F�9�	ĂEJ��n�пsr@�����`۩uM�b�%��c/Kr�8&���QF��gh�Ԃ8#o�#��P��o��ݨ"|,J�iH7�zD;���cl��c���s(5��� Y���rt�9Ui�����1����3t��)�׷�,BKA�	Y�@��f7<��V�9�`��bsL��\8<����]�ƀ��󏏸��^#,�U��x��J�ukӾzc��n���u�xbaW&��a�ضХ(%f����!B�o.�MP�]5e��/t��T;M3_�X�C~�2[�p�����Ɣ��L&,���b/�oৣ��Mĩ�F1�9�9y�F���a������,Nn���;)����&��Bn@���Ew�����+��M��}_QC�<��l`��˓���j�ʏx?�����;$jd���GH��3xIlx��Ug|�L��໺��~��ӌ����B�[U#�hoZ8�����[h_��Wރ�nsh4�����m���b����v�N�BQ#�҈xh�:[J�)��Q�EGf��i��<L�ƨVf�D�&�������[|���%J3(T��~�aRaS��#�LD1�<H$�Se6��Y�=g-E+�������awg���p˓R,�ʶ��'�p��w�lA�$i��\��v����&r��/a�cTڐ�Z���m�������7�J�L3�j�zR#|;E.���)4	��B%�Y:��W;���k�~��\��Kܬ[ ?���UT��yf�7�˛�qVk�PQ;�
w0��Q��q,X�I��neCYCE�6���76{�t�š��]�d�C�WEc�ݔ^ԡ9�^�h�+P��Zc%VݜlF�VN�OߟrT�M=j���fvQ�e���&���>~���Bu�,�F��`g���^U��~�_�8����8(��	��Fp��h�UP*�ǆB-���C- ����˱D�|x��d�u���o<�%��I@�(�m,��}��ě�CX
��Ǘg"��c:�"xUW�
����k� ���.ړ�d����
��l�+nz�+Z�I_l*N� RP;�7!��gh���# �j�;�ʈiGe�y\��P^5�����{%�5T|��*3�V����l����x��UM�ϛ��"���:������H�0�L������v$��5��煐����3څ��~��>�s��o�g؛ݹp��_j�8S��Uҏ�ھ�	�F�^l�y��qmT$�5R� ?�!<�'Jf{k�o����D��Cu0*�ICR��sa_����7:����	��3\�Z�P�.�W��a	�R����Ź!t_���M������/OWn5�x�m��s�k|�cAatn�`��.���D��e�S�0�a��G��e�7�3~��NÎ_^��W#��L�r�S�n��x	u�,�L\�*�@�8:vy��a�[�72�{�.�\+[w� �i�M�� ��rN�EC�Ӱ�s]��3#l�Y�4D��5�&�8�q6��ChI�2)B����f��c8�uC��H�ƚ�/z#8�Qܸ��dW�ѣ���^7}W�џ��4tdT�٦M�!�cCE����ʧQ9�ߏ|�ƪ������9}T�L�׌JI��*~�3~-�
�#��x*��mԇ
#��%��V�UIґt�P}���v�*��^b�yWź^�Xb��4����o9'm*�h� ���D[����*,��]�bu�f��g�ע�)�w��=���dẙQ7��0j���c���IοQ��[� D�=�b̛l�x,JI}R�
?UxK"u�*�sA�F.�ZT���|^�2X
�1��W!I�=u݋�����"�5a�D���V�7ц�{9]���X_�r|ܣ�f߻n̀i��=�K�F�>!y�Q��6ٜ��ia<�)�Q:��;�Yof˺�y�o�>�gO?X`�KQdl0!
���tk�^��J#�L��W {v����1E�~��]�5��<�Ҍ��>�ƶ�4C����*)V�0��)O�����:��w�8볱��,�%�?����8X�����|7edg�����S�'9�8�RR�ۑ�g� "�B�_�w�;"�_�g��z*��zџ��G�.����
J�{Y-�t���!{X��@�����ib���m�
U�}�M�����������z�	S���7�7��