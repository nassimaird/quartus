��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_�Xr��O�C/���.$;�����v���?tp�����х
��:��0La��}؄�6Y�Qџ�����n���_^Z���>�((3���&v)!��Y����ຓ��{����!���,؛6�h�:	c�6&�磬5��8�i�s{7R�-�>I]��-HN��F��x��ވ��޾�N��g�V������W���L8�e�b�m�C���� gy|��Z,F:��]b,���Rmb�PF�.� ��\�}���>��<E\�/a����aD��YRA��UI�%_�ڝ��k��0�޺�C��qM����r.��S�>LUp9�gqg��⤩6	����-a vJ:~X�!)
B�a�s��č�V�D\���h���@8B[9q�
d1��M@��� ��p�t�\��]���Q-C SƔ;v�{�iK)O	��q������!!G�xOdjR���F�X����:��Y�~W�҃͟�Ab)��f+n�3��ꪎ���gE��<�[C�Z�I�8|� ��֚NӦ�DBA�uD��WɃ����%�!���b�顨�.�����ɦe��2�lEM����(��ڡ�2��ӘU��XMdC/~Z�]Vְ����dA��'��r�q6n2<=a�T��fMD0ӿ�L��7�A~�R�1�isB��.�shO�<� �d�'XSyQ/���55��2�$ߘ�6fOE�Eʽ\�>oO{�����eӶ�o�钐��7AU�j�o�.e��u��!\��.OK"Tq��ƞ6r._�B���|��e����甦�.�`�R���K'?;�A�*��l�%
�D8�iKR��݆�%����,ǚw��N�eÁ��4����=;��?'�u5��ƹd��
y�~�	c����"֟0����-aC�g|!w��i�q�)F�?G�fRlT��w�s"^lD�a��řK�m[����:����
�v]���r��t����S�55����}}!����|Z�t����ǉ]����5񴹏��W����"���:�cU�����N"M����3�[�n�\��>wO�H��z�n����F�[��q�y�JX��=�Gܢ���=<C_�{��d����U�OfϤ2A��5�>"<��������}���pU:![48�8�'�<�{F���q�w=����jYOl�?�4��^t1W:���k�����'��A+�|M��Y��%c/~�:v]��z"@k]=�gׯ���	���3��er!�v�vNt�4�]k-�(��k��f���ئ���|-#C*�-�y����
ݨvxg��8n�χ��L�z{���s�g�V&;;��[�XKq+}J�f���s\��2ƶƪ�'iY{Th�+�#�ZoV����t2�k��e�)Y\�����B$^׎	STLƉ�,��CT����^:'ӘAN��P���Xd�t�6���w2y���-��To*ʣe��m���I��SA�h�SR��g1��rg(����p�tin��M�~��][PF���C=迅p@�Zxzt�����
[;{Hl�P:���&1�
�V��,�ɪ���̭r6�= ��ۘ͡���Ñ���:��h�1�i_2.]p����C��@Qj|ŗvȫ
S�tëk���(�9=���)P����{��T)�~H,E.�q���O��ԓ'2�.��7(SQ�=ͱ$^g�E�%��y!� �(e4��Hi{���g4�jy��B��!�� �7�y�(J�81���X�]�`�����WF6�uz���~_+"���qsn������|VG���|���1�w��F$��ɦ�(�C�՛����B�2i�yBPA{�1_��nY� %�^������H���:��祐 s�~$�u
#�:|3A���*R�y��Z&��pń��`��~`
�++s�U�8HX`��	W �a9��V�bF�Sq\S������Uu�U]�Kw*sd����v/Glx��s�!��e��\�1�X�D�J�B�4[���$�$e��Yf~�%�N����� ����
���c�@��� ��v�:��u��ƶ�lF�ЙaB0�'�_����lx�=N+d��w�'�������V!H�v�>�hT��"����76C�Z����ի� ��m�;�����516��R�'4�6�����-j�-ი$��sG��O��sl@�v�d���w
i�H3DFR�{��񾄏8��p�!gy��A�	������6���q^c�����.zH݉نR(è �����_>B�,
u�?�[������hL�:G�߇Ϛ6m���	�ƪ
��Q`T��;�vN޸y�Mq���7�l����!.�{��3��C�#�d�2���1��9�C=%�ǉG���%�z���n�z��b3롹OY~1�v&��+��'�>C�=Ӗ+89{�b%GF�%J�4Đ|O��\.)�J��M>iI`�4�X�f��S���$�w|�'S��SF0���O�(�m9��s�k����*�ŗz�ܞ/��#��r�A,�*��͸���I�:wq�
e~��c�N�o���uKo�C7��Bb�:=��n�W<�C毌`��[#sLa�F�����J�W��MZ�%@C��.�r��լ>�4䝻�(YЀ�UR$w��F�j�p]ڎ2�F1������D��7�}'/�vѨ`π��6+X�l�vZl�N��cn�kcZ�RN�&�|��f����I9N��c;�)Ŭ���_U��!/:~}(o��J�b��Rw������a֭�M99�?D��U*Q�Nb�]�mo&øݟiS}�E@���E[jX��������G��?)m�h��\A��Lei�wl�ݝ�81˗t��?� �̩��r�*�18��Z�`�T�2���}�Dͷ�a Bg��zӷ�j�\7����W�+���2�RklM9�q��O\�pQ�.��Wv��>�~ɓ�V�2Q�{}@��o�؜B��觰��`��O^�b���Gs�_���h�2���]���+҇ܪS���QI�NE����wɥP� ��b�h�����|�O�q�.i�y������Ym)�r��T��J�hͳ��${ʧIO�,��`	���C����c�b�=��F�l��!�x*;���<��Y�q� ^(F	YpIt��TFdo�t{w�F�	@"�Q{�,Bo_��ź�7���^t�}X2?+`6;�ޙˍ^h��Kk�O��~������+���&T
7w�Îe'
��?x�x���!�L:� ���<ݏ0�)�a]	��H�Z�U��;׏:����:"ɨ�Lrc.�-뽚���n6WU7uZ������4��ݨ��	�Q��9r��r��L!���n�O�Qd$&��V
���D�&��m'ў;8�O�� ��XLp(BX(pϕ��Y�<��G�+��zF8�`�"ƻ�{pگ?��w$E���ی�`!#�J)mE�;�j@R튤���vʒ���-~!oOS]A,�ߘD���n+�aǤa���Qj���>z;�*<$�����(U e3��l)��5q��bK��o���,)�G7�ص;�3io��螓���Cw�sۑO�ệYW �x�4¤g؊p��51RnsT�I���0�}*�Y��B6q~%�����6�S����fq,{��Z��fK�o-�V͏�!�(�`�?�xi'�'ԓO?v�.x6Q���N���f��`8Z�Q���FL-��몡9��3�gZ��[I��[Ѥ��)zC�Д�UZڑBޓ�PG]��>����Ύ0 ��S��q�7�7�����Rgq�?i)W�'y��`UVZ V�>m�|4>d�;k%�ݧEE{�3p;[���!�U���2�G�&���>ó����G�M��#q�$�c�ы�1��G A�kW���1�Ԛ��+��51� v�l����!4`��ci���A���ܣ �&��L�4w��:���,L�Yp� Ww9�3�
������O���բ�"$B��[Dg�w�Ol��GB��߿W
���-}+V����E�$J��:�>�(^\ŋ_�}6ź���`[����{��ҝ��/&Ķ���/�x�5%�)��Q)�E��K�1���\$n��"l[m-�ڔ� Q���:�Y�ʴ��F�܄:GBi�`���r�)�#Dǉa��GBj��~rq�7�� *�I��=#�8������� �+7 vK�DI0}��l�[���ޞ��VD�C��Rp(yr�Su;��ߏ��Nci[�><���@�O��%�C�p*�н R�3�'��k�qh��/9���Ǐm���[�M�2��`�'F��4�	������<�S����ɐ?�E�D�Dq�hq$���{��#�Q��SnO�q%:D��}�T���*@ԫ���LuLߏT�u
�� �)#���VWK����o�8������c"��c��?�����/��}��*��䓯p����Y�y�ywA���#���J�ۊ��>_�g�[�,As������J�Ҕ����@���X���!�K�g^����sP+���H4����9�&M��9���f\QrsK�-ho*��)�� C��S��)簧���7L:'A�%v��6�F�/�cu` [�T
�0�s�ɨ�����b�U���9��?��$,y{D�"
��\T5�r� U����3 ѳ�	����w�iqz#����t���y#�̥?��<]���JZl-�k���>iٌ�i@K������ Qci`��\� ���n,�.&���K�p[Ma��Ӝ){�^q3�����Z�v �Q�Õ���6)�ă���]�?]m�`M� ���ȍ��Y�9q��t��\�>l���y��	