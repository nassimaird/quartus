`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KKM+2AetSP7P/3IDJz+LIuFCeu5HgM1HRF3QW80TLTeV9Tz9RIj8yLIeuudJF8o1
UAFgq7pPXCA/GvuRRk9HOxVMjGT5+hTizQ3E97ge1jSHGwouZCs2iNw14MH8syse
6yFNmO+GJtX+5uho7rJFwvbFQbZ4CjO1sWiCFhFcNV0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5888)
VpanyHKjOcCrHBR8rG1HotaN7nV0GxADf91dZYApBI5w5k9e5syyp7C6EWAZAOwP
bHSdB04I/qyR8QqRAwuB7JWwFPawCn4F8Oxi3/jP6eL4w9i6sEQG0uMIV/xaN/N3
Ea29ek6IpXtMTydhF+rulEkOozZHYxb2y2YpihPU7AKGV5HJlCB2zAugzPPD5d93
iXZUjTOk1HVPc8+oSS4Mt6TdcuVRPHlfy/mi00Q9Uvt7yMYMFrvA0SHl1HFKcbk7
Nyrjw004m20VPN3iJNrkqJWJQJfy6fA0/fNX3gn8jKIqxiIPxYiLR7iwteZrOMXX
/F92xgz6/n80NnrNVFVG7XiJ6qcQgtA5QP2shYVslxF7i6mIsEYzIna3ap+Skjjx
DCKUByIWGYzFxUdNdVA91QQM7qL3OppXvQ3cIT0vlZorYrCrzcjhtsFDaY5fPuYR
2jLO/1Y+kQLaRlileZLVQeUT8CJ95zHexcGijJV0y+M7h+30GcxKI8Yg7yrwfBAH
9kNlUyh/8OZMRXr0eNAIyrnjr76Zq4gjXwS891BqinzjWzOmPjGQoD4H3Trlq6xb
O+YbdpgLt21PXaKXe4GCjQEu6e6jBB2HbACU9xaHPm7c56GFLRPLJlQWC2jIWCLL
a255nYXw22H56tvrQ+Gkrz60TzIzRzoElGeczKDHcPh3kvOAkc8cATwZ8TqH+dSn
vFJwAq5LAaA3SxOUKaYNaqMJAdCa3oVmljYoIcQu6n/rL53e+pIaMwpR/wuMGyaE
A3Bln/kXivcWu9DFtvKeja01RXrpu6dwKpYO5TFR5t9QPCV0yiB38/aKs52mugiZ
AuRde8qwPbaPuWr78RLyIfIWPSYzRHNYOSTh/uRJpMXuQAbQL1ZyYgDUffoPgejQ
8dvE6qq/jJxxFwM7bkVB/Cn4tSPrwYQM+AZQ6R2uFHkLlZcBfZZn+KsnNe6PW87V
86uqCdl3J5mCFXUBzRzYt3f5R29QC2D0dIRwJEi7S3y6EyllHfP2FA4P8FbRsRhw
Q7LIqsqVezDlhxfTCVg/C/y5NGqbWepmyrGy8uqSsRX9yVR5Q4poTAh3sHw0Ed1C
nNFlibddUphtVnVmwude8+Wr2ttQJYXEShqgv5/oWRzvT9GKwqF67v5EDEEzqFSq
CG+qSETupznWAPgS3ZSyHO1vPPlrWk1cPN4u0d5bqAJ4tk2qenCY8/Y2/o3sppey
1fsampYALUd55u34Vt2dyBe4WJCs7oFru9Vp3BsONM9znfNhDNnpuq431jCkQKD/
bnZxP5MuLx/1a7fa/78c6Xe3+d5uVFVCRRXD0++cZT68bnKd9SMJx6mSV9tFQubj
KRD95ROkcTZTJxTuvRb2mLBIpgi44E0UIHOBycZnI3EhLD9gjevA0XIc4ADiNylA
+WA1dEKPNNjImHSQZspwTW0gBmqaSAT90qu33u6qJ0yhsiryTy9hrFYPJJSV4a18
KP3Sj1lpn/lCzqGKLLNn4e+R9fKHHg6z2FjOlgCe3ef8hbHuc3bZfy4vy1CZn1VT
7wv6fcy+/z4LMc4D++PdGm9T61cEnzLGxsB4brRPcOm3ZHvCPePBSesAWKaAL5Ni
Zf91uP+wMeqvnSdq9Lzf04WVDKe6eqy95Fp0FkQmd+FgmT6xDIjEew1itTNOS91Y
piTVFHARJBX5OzqMPgzCGinPb9VrBscNcwtfwxbq3xLcQ0i6jmoixXGx2WX9ugU5
piY46q76ie1WJKub9CM1cHO1bTkgJzfMrQrdV5n6Rb94Gcq47WKvPeCSJLisK9As
F1p5BqiXnCX4lYvUSIr5cElk6mp5KK8Fdq78RedvbT72edK542bTIFxmIx9hJdhA
cy5zOvAuq9lAUwn7AQTN8RPgQRLwnP4ZNzjCMY6Kbvi1SupVwyaEWEvw9FChUvB/
bWGTMnAQwRYqiQIbNjHJOzxuFRFqgsBet8DmVRNcji/ZPEMXKF68CiIWyanmGO3/
eb5+9FKv7qJTtDnpKukHowYpIWuUit32zYw2IODLJxtfKUvXbOIJ0BqBQHcR4Iss
mLiTN+zXkJaW/6aFFguq27SX7CIUsQMz9SO4gx7LftFoWVgt936W191nhZoy1bXW
xgBhqj7DaQq0CZ36eCB0FHz8X7IXowSOh+SY/GddHng6bLkk0oqMbuCUpTYXgNog
Mqooee/+c7RVLUjBL0E13vJZ3N9X8I7kh8NDlSYea+qcqVjFYEhrHnbjK7LQo33f
gtmPgSE/oniaTCdDb4lIo+AVxwsjHkew1X/efJLpYbNUE7UATgPSyNX3uSGQ6oDH
flPU9PiYsPzi7yYq9GTplt/2ojaQEXOaVenJathYBC1hLFgUymkeVD3EpiDQTg3c
J3H2h+I75eeZeHsfvQePFYslaz5sQugpZnemep08fogerse7VyuyCE7rWKUrs/Wm
OA0ZLaoDEyr1jTkxe51XxwlQGXpePGrjIEiiaIsKPNBBoj0ik3CUN5wb94p5WsZf
KLwa7ImJgVl3ACOPaUSAydoiOZ2Hp7V7oQx5ct2dia1myWSWw49VxpjRqk3PcNRs
q21jIzjfPCQL0mpmto/3Os+0FZo+2dTYF5gxWsJpz5dCu7+Tof1sY9+t0LhJ1SCN
jAZx8ERgiqk/ODqw1gEMO5bmk3qZrszSa2yVhzJEe+B2rFatzvmDGPV980xQ78oP
UNe7jA5sHkrBNyi3W7cqU78BT49zpSz6s2DaftgFyqBvOlTwUD4hDW9NEUWKk9L/
hkOmwGbpcTZYDiTx4nrPXoZGqEV4QIMhZQraVQZgiarvWQ13jyLG1TOdZrvpHvzF
FyWxhN1YX5KaWNo1zfyT7GynLhW/704DlnARQ58WjCrvUW6YhaL1i6LeHxNwokV/
+0NM62yKbuLdB/Oi7TaT4pTQNm5mmlb4qQJQcwAQDJlLEs6rqKhoukRinQzPoU37
ga5NrbjMmW1xaRGOBVt2dVNuzErUfBOw5RM5FBendPmwizRWaM5L6SP8B9l5DeIj
qFDwvPM4O5RGBpThR6kNkr7IzGzgzSGP2l6XjwLuNVc3eJlPnLoOW94FTIVyLZHQ
cKC+V4OzUwejZr84VWoZHn6p9cHGpblzNAoYn/MBgRsF2J0VNUoKjh7I5Zx3CU0S
xGOF6/Ifx01h6+TapFJ6LjsXOZbZto6u/FL4iltoLQlWwBoTjV7PXl7NcG4P7OH1
iODrM/fFvDeJTlVLFiMYpr1tiwoiJ4O3noKINzY/nwZlEoUsYY2I3UpMm1U83H2O
vA5W/o1Ad6oCrJcdmV+e4h4tT/lVtb1gokvo2RWrSVMZz41QO9yA93cLvk+dNstV
bFs/dODEuaBx/vuv4OCG8Zq56TT1n+llSZb0qzN15pYucvcOd5etC9m4CxPTprvv
iqqsuVNsOA9A6Pu/aW2NLc/fxeke7a2Cc1obALo4LPVaOeyzwkrW6MuAm3vsRoVy
34mTjIjqmKqrNExh8ko5i8Oe8lxbv0FKLAK1nJzakYJSegx5a30b4UocKBVHhxNI
kzJ0Nem2hlR4Fd9Ci6nXVcEJEIoXM1JcIqYzeSYyzXs2TFOnnB7P1Jzvf0JIPpLT
7Lzr+feYYar+7re5UBwZ3zgDX4nV64HZgSZhkTZU9vFjt3pvogVPoJd0XqX7/RST
2FTD/BzAA/pFER9bxtXNRgsoxhW0g0IydJ7XjSGvGfACzkWz5OZu+8PIXw3lIGwm
k42FKitPv3t08lvbwll3Ri1mZEn/GK6+EUAeR55ldV1KHZeTutv8VliheFBtsWNP
oLIExQt95QtJAe1ya0ETpxR+kiGOr6MLzGZl+T08PAiZRxrcKpxgUi+qNKoRzlM/
v0eiiDj6y557xlLKdGYz/PrER8HmYFMrx5QUxyVaguwTTpttyZKOmBGJPw+YR8s7
s6Ia07wUpVidobJ/W0Jm5kwJ488yBDcpSbgA7QXfmEH3vtG9BmVIXh9HCWuLJCk2
HfYxoQlAHjlcG2EuMeFltV3eFMMI4Le4rbOnqrGxXoydQRAuROOfesxpVikiCSc6
iGOONh7lWmUdA6Lr51xaupoFUZCzJwBSUnOMhzmkl4Ks89sSt3Y420hwwNasiGbZ
tst7I5NV5FEN9B+JFusxNKW4H+IQfznvn3MPfSIDpibq4Pb4xL7jwI8fgsI1gg4S
4/5g3Bw0B4pzrvET7+C7H9Furi8LS5VUk5oq1y9P1sUlqjYfag47sX4UdLBeBK09
EchE8sbQW26algjjE+eBmHNbO28K6vWZsY6dK/ZQS6aLyMueMc/XkEx2FgPQ7Vcd
6ZGssB6G+GUDTozzHZcOMb0hGtNtxHxVQKEWtEWKzl3wWtJisy7JTiUgiJ24G3xs
vlEuaqTEiiLJhbr0X4CELhE9lVA6mtGIFjZjEn6yCtneUKkitCQvySc1MFzFOOzI
cOM0GiLciNOP5ziTlwTcS6j9nyompiIEuVQQZHapFmxMvM+0SyjPYWdky/UoKbK6
liiBoaIQgLHVys+M5wOmXJNG1Y4Cl2WINXBWsOLkJOU1ONHKaDGx0QZt665Fr0gA
k7wDfhrSTvnDAFB2onGhaoBKdtzl61f/a8q0qmqjyJw7Ix7Z/9jOYWDuAsKv+bAa
nvFhWGOCpOyIzW04O7i1k4gEVsr8xzZGqHAPrumzvRQQelsMvgKEro6vf74UQFhp
ANzs7fSuhqwseA0O5pvvpAoxz1Ph32z8WM4JSi29eX6t69FBhtB2Ox34E+reeo0l
lnZX72FGto0F5U6zXeWj0VFNGqQ676tab250rnvFw0IyNQms2+EtluqjYmxWgVPP
MFhYIxrpgRnOvMCpLaLi17rLP7twWq/JNRGM50mqAbfRgGKJxMlR7ocJAZ9KNwi9
uRmaWwTPfyjDex3Q1pkS1ymzLnFVxt479s5kIrhjtxBn7+DKjQ97zqR6Xj/1pZAk
RMJm5tkjQ4PbDIKKsuu4G5RC016HG0TqXl6xlFVc71JYuzxFmcIzpaoO7fuMAUCU
Oc+jax+MQs/s3d595rkMCegoUECrLiHWUcNcWiedvV/f3RZH5Jz8/U73GbpOoSah
gczF0Tn9J8f+dI6IAswudSP2UVikGXGk0XmFN4cOKgFSPPC1N2cvGv88XtYTYB1C
7HSVadUVbnGWj5uv1d1ylG3u5NbtPWhoG3A1urT+NW8gIUlqj5o3IrJ+CriaJyGj
2CfD5dBBJCXlLQUwGn1c//+iChQ3daXh2s0VmHf+mo4FyQVU/HpbPE9De0h3A4D2
xb82TL2Lpb/vDMumDUOiV/FKBDn/tn8KOUsXT9Y8A8T7b8Add0ki7awGMQM8AEOa
UL7QGLC4XJy0L3c1wy0+jRNzigPkgQUC2eFULPXa2/JAtn/6/0XllMYnca/HRKGn
BflcHKY5NpL48xJSP8Mbeq18NT/KpZm6Ua2EVPUCAJo8/TUMiZ6wEfcqXZA2iPLm
d5NDKXNxjJGHp4UUmVC4AlJzN2q/g8Ir0iekjGksOo2KOLkymkT+PkBqzyiwW9na
bt0+P21+53EscTeGXaQyHs82U8UG8aMBLvN/8A3gb/0XME+JMsip+hL3WxRYr0RS
DKm8U2DBEz85AYzVHv9QKDEqKPEHkvyZcNTb+Qg59g7KBO4ghB5zcpRUq5n07QUG
TLj/mziwFdL76B5v4boITC7sgp7OuGe6DupYWEJ11N8uCAPFa+FsDYPg4co6KnNT
EVGyco0Dn6QDRiGrqbaI73LDlSOCmmsdzNn9aH4S4DXhcERVEvUXNn+muDdDfHdb
Io61+szJ0CFD5svCqPMSmCxQOrDGBQtE+lzstlwYG4jsF1CjKR6lyenMIqLFuzlR
eB/QgAoqdCcgz0e+6o/mLzzg/eYkMZ/ORXhGjvqbnxiyuBnKPxK9ZIrUFiFYfCyd
Szg5PAyPg9AUHivZ8J65a6u/i8mYOHgn5uS9jFPEMnV0jYGrjWfuOErbXd3eYx6l
4aVZgm89nwOwqhMwB7CQQcdQHXBHuqzkaPAYe6KZTK07IxTIYX0jHT9TbNrKb8aI
ffJtc3RAbvcUiZdtZpmGZ9DnfeMnMkF5Pf1UZH+G3evpM2pE4vRgg001Fjhrvjs+
Zf//mXKSSOHuzf1WCB9ms1Jt1IltmyIb6m2YfKkEzfLYAWjc1AvCicCwuiERJE1X
WI1B0OMCsAomaLqh+p5n204mvaux3XtgbCu5p0A3QxERi+iGRQKiCkit82LBAUSa
sd3a1T3aweddFC/oVR2PDpFf5CIZRgLJ2+S0do3ZoQM3jFYfqVw9m2zaFutb3XU3
fWoM/VozvB8YG+b+HhHfVlrUdNHr6AY0YNDhRlIaMKSMvgPbJ8gKt25uaxjMhQ35
eVsx6xzyoF3MAfc0HoA3sFIGtJ+GIL4Y8G2v5zQajgfNpSPMqEnG3EBNAoI4MgtU
B8/Ewdf9QTj451WQKFaHRuHBpt0Fl/HZIrrvigTSr/pRasevBrmxy94Mr5OSmgal
XYAtFUHDjqUu6GgpuGikbuT59nUbRYhlE5s+v16ZQqiFBspa/1hScZ14mwSYzRd+
SH7rZO2w0sc9o1GEW5/VGL2Bv/ajI4ZousMk4DqQVevgZ2Cun2C6dvyrOmVpsMAx
fzrmicOM0C94sLfbdvTsRlKgPELektnvPhIVQ5MgrN5QfpjD4ErC57R5rX+FNBYS
UzLROyDP1Ytp1guWtL6dJJ4YBcsQ+n3UERv5iobUbZyWo99HLag+5GdFQbQp2Mgw
J/jrxMw0ZKW4OUZiegTi7mRIzyXHseoJZan8C5AhikaFx5TcgA6zCqvWHTZyrZqC
G+NhL9scpGUmq9kNUwD2rY1j0vDzlsmsuZiLeOZjCtFNXJ3x0GHKohp06LIesPNd
uRcZpiuCensb8vPbEhOHlvks8sx7YxRsCX3+5Uyjq7lT3I81l0UmHZY0DaOO6V5s
zik07AryTttQYBBjOgBVLAVnHJiQgHJ8i0AZTXgiti027YwfEl1DeVQqVDp9V2Kb
ij8X95xdcuE13F74xXG9sw1shVca1XmoAFcBTVc8GepeuC+eQnmEPpLfbbjum276
gj3GDdgZZA1T3ms4OXY08M7nfu8Lh68bf30Y9ufXFAyXvci+34MQp6PFuYob+Bzi
6lgsUMsjPCj5JSuFwOxEVKLzM7y2QZarHoK8zbrB1KMMbylCdAXOYkja1v4JUxnQ
4jYmVgFZjrgVuJFg66dUVrRW0nYcu8aXJVSEnkEkg/jcb8P9JpazEtMiyvuCqUVl
88IQfayDlADp4dknOcqM8K9WEsf1/tKgIrxQASadblKPUCjQ0DGwLvQgtYBeNZ35
Kx8iVVtnUKEI547aAqZ0uZA1HJhMN6kB131oy5ZjddbGlNoJeZYgvmrznPfkgRmP
E9v2zdBmcbgXre9S5JMBxCMz8LFCI2YxUNQM665AGf34X18clQWjGs1DmGUXCtNj
8MP2UGttoyfWW0FS5oBIQoYTXIPNgQsvDPkLaOc+QKtvrN3ucoFkbZ88jPwte+Yh
VUQsWMvLA3EvA8udc0wCCenNkAdEZT3BkBQlqIye4nJQfEzo6r4zSRcaPv0lY3CX
zlOl1tiGKh/fuQ4bM3Y9FEAYZTo0TRd1Z13w0iLT9wsm1oACBCyb3kH/bOdj2PoA
ZKYxJP5BIBkIWL8Ev/kKVxNkyrdlFyaOQ8PNeHwffHdkFd65tUEwEey0miHs5bU9
okVRy0sONb3EFjukC1k7H8wwz6BkcOFK8epjrLmTD1sARkH+SLNXL9+E318Z/H5j
cLALD5DnpIIY/uzjzE9b//xA/45oEMfOMkkC65uJTIK3fQXrDDUlprvY14UCizsa
XQnW+pFXYRgUkpCfDPL3iEl85a3Pcp6oHE7Yrczr2Mc=
`pragma protect end_protected
