// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
frAsrYHQQj/a41ncCu2jcg2BbdB1uK7sM+MiMPL5eXadlJ3zY5rxeE11Y+VP/WYBHqHSLxGx2Cll
6cFx55z8E4ORCIyn2usVePqhWFGgpzaXXnjNuxrAchfXNRDj0+6y/8ZyMShZrpndY2L9LgA1y+gO
JaWoDxjwp6TRBI7CfP1NkT+tToc9ohQZ+XsEcVgDkv0EdAL1nmmJQvS2mH1xdMYVGl3PWyL0R/b/
j2Rksqs7vPcLRYSLgxn1jcKpynHNlmA4/8OGut9qepTXTRTjJjkKILA3lUXyf2c4Dv4gGQ0yJW4R
mFpH4pM+zvGtwSZMyb/FHey/ntFPCZYFTQdp+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5552)
9AxRhn0vPFjqRU3Omcm816u/5EJZg0qROzpaXoL9Vscjtk6RHCkdTLTHemmfrFaluQCLQLE0IOXr
DwPP48xTJei/yfmuUG3YwEAoRN0byQ9WSJFnJAGc/7H1dJ1y+y+8XGfNwB7+PsQFsn2ioPVyPP7v
k7sIJsVBtNL4NHJnGfMwhb0e2CLxtua3QCTd43lhiUMqmgVwv6evHFx/2H0WqMtdq0ejHFUk8QIB
4SnwQMLtZt4PhE+voxaofeQ2y5up6wfBSypsVuheinZz86PlxUeRRQ9BxyfCfaK5mENhPNxN0aVC
A2wBI9SBfZr+X8y+Ia94+fQznmRjOouH+Waz3OB8rY2kqY/13UukCMeRBWSMv1h2NbhuhyQaB4NQ
NkId2jxVI5Qrw80kLvscnvzs+BjfWLvTLKLw3lTnS8FGxHeuDuorJ63i4FJtrTj5TQWUiEamCfNR
JBZNaW6Gns83aovhk4UHF1cgyv4Cxb6XlSf0qP/rakhGU6H3wrG1mmKnK4CSK0LgifAzbBxqb5Kt
HVwO2csBsXJAkPJqgitm7jK6H0wQvqUu7Bp3ZaaG40+f5zda0XILk19UXa3GuFgl9i1o3Rqu3rgt
YlvNKhxSagVQCkihWK8JWtWxCJZN6Jf1tIMAmPlNVzAyXPP6dYlNNUb0AREtJQcSxX1RdZN4c9Ia
D4naItREkEXqPE9jQYGinTEuUtgBSnT+zBQf8NG9ujd+S4D1cUKADn2Nv1qrowLPBN8OeELdg/X9
BiSuKGaYXbgn5a1z24Wx1CcR1pxvlYiTJRC4XCQOQUBi4eg7xlPb/p1I0QdjYCQmJBqkZapzly3J
3LuzItUDDk5Y84ncogA9J9/sOe0tBe9gQSVkqXHU4Hxu+G/sVWtv8eUe2sM/5Om62ohMX9/iTuvP
g1rxuWgOkeFhJW7xYNUKARtuq3mSzY5YCYFW9xymYiukiQprsX2OJxCyKUzlzlVhBOAgHx81VrB1
ARKoxSsCch0ThEluo4SsjwOCSuUsd2iIhLrbbsUmr4ZVP4g1qy7QdAwgT4li9tMq3gRl56ZrAAFL
8lTNSr0fZFdHvESrn3qMP/YQZyiM8oixtupmNYSFxk4UZKGzgb5JxHCag0Qgd/yJJYNP5Wt/W8GU
VAZ1X6tYrl8mqqgLj553lmJURJ+97sws9x68yv0xWwlPjzxY+I40hoPr+xfpzfQncOWZFDmdKjGw
Xak8XHD4ZHFHAmfMzstUhDaAC5cQ/US9qyJrtcZJd4beZMqOxO0e9APcGw/j8D+V38NA5j+wsY/I
N7KlOS0dFsL3r5dKhYVdX3j0gYA4GJLe4EAJVZWq5CS8ggFBelu0rFQMCxG2vBUt9UnY63aKGpgz
/BMXx1QzfQEIpdrYLa7C4Zo3AoN5PFffyqvVWfqNByQMd7lu0pSWkJV7OlrJKeABcCo085QXycIW
e8DfT/YPhPj9sR9LqOn2//epeIUXWHf11f/lR6Fq9s2lA2kArS12BD2HO4jbN+jPbRrGl/IdJMqL
+d9GKHY9ErDRVNJTuhu7a84R75uKarAWwYYnK2CRuX3dPZjVdSSGMU2hQznUYKD5a1We02nvO32t
8Nt6mjRo+iPL7Za6oK0g85Dz+fySYAc/Xh1jqRXVOMQ6edb825GHJ/Jdu4Yh9AqGCzgUuh+0y6TG
Phvr7i7eXJOgbG1KRhdca4/ry5da38wlszKo0S6C3PHHscr8cSBMJvwv5ivR+qBWRwDFZHN8Pimm
exlHqgIi20/rbzWIfABlU07F5nLFFa1WASYjsZrppM8vcBNrrDjEK0/9rF8l63R5FXtXCyRlhrjj
41SyOa1BqcZapW/VUgiNoWTC5QI0I0o/uwt/qtY56tqG+BBtxqIhiySUZqqcNJq2YksSrkFjhapk
zyloRwSkmJmp4K2IxfEM37FQ8boc0afsbOQdwrv7JaHOM2ba86BiV5jFwqnCOXYY90CDVQa8B23I
gho2OKQiubrSRhvGmsS5GGEvH8CxWNluWTbb4J5ao78fOB9MpNkhipqUFwq11dNRslRLdiL0Yyp1
5OpM00RWuS6N3QGkLR8bZxrqyb2baPsokT4AXp3eBSzM9+jtZ7WOPUxOhIAPElpu4if9v19yDL73
XtAWZZUs4g6e4m6/2ZoZ5cEa+JKb7fWbTXtxXYstu0G2zGihyzWK3LZEibMf/MreU1zaV2OT6VKT
52QQ5pwYC6iKEiPLApl+UnAiLVX9uGOk440YGW72xtRI+6hUumveZyIPGnj9/XCcJfGFg8UW1Mqi
h5jtnSxjIKS5gPQoV51UHMUQ0UfRzdCIimjtDuSush5WNlaKKC6wG2APm31tfSJajAxhgkv/4UR6
k/OeDlwBy41ka6CbblsJa4IG7QA3sfLq5Ho8eXAFSS8k31K7Iq+K5421d0fS8iKgrC3PTuYG/Gix
b0CnMjldU4dUdba8FKZkuPtQjDSXviTEye2ZDgZi5MrxVca4+3CwH1lD9VmVnLpgetIx2Si0wqZO
PNcyyWheb39veB7IqFYyBipYcjd86PfuuMa8nxl5tHajjPTr487OEq6tWpZ/GTUXiSP1JQfegghp
twumjfUWdm1AR1XzZO6gLlGTqdh6PftpHdateHBYwTgD2UoRYBCyHC4D6ww6goDE1R7EXby723vg
La8DNplD8dv0CNfRMszPvM9Vk8/Q3YuqUYuOmyTgVKK33JwNl+sKT+w51Auhc38cmukVOt7cMyok
DKdIN3ZBb6a/GbTQ7txt4c4S0NBOZQIsemp1gwu0Ovst40Wppbzj/M4WhnmwMQufWsXlMVeCo5X5
kT8wPpYZY/1n7ml0y01svmsC/9XsK4/qA1isc5db8Ucks2bg6qTC70oW8RbgwKfxeYmrKgasw5Cl
vDtjPD2Q/5k0ARid1LJpZ/X68Uk8oa/IrUbIyokllNZ6B5MmAFo5CAPiemTo0WMbxz0Oqs1GbJ0E
hYlxNywWcfNmwCRBHoSv+iH5NeuuEQHvcDPV219/yR0KdQMYVt5EdYRsGod1GpbVv0zUe0Av1r8i
Lk7kAqr9fNnmXeKDrtsjywxD2vc4uKTaKkI+fBzoRe7fjFx5kctmlSGk3BAxgHpQMgXpoz66DuQc
4ciaPXWXBaBejFWxFiiu91Al96FbQP64fU0INpzY0KzD7fNGPI5ckgamNXKl23rVR1f1eX3uG54o
EpKe2kOIIB+t/9yjx3HBHWjzejHFc+/o5IJmfV/7mH/a1CYFes6mCaj7VB+JYp6Ye0sHZnQzdbu5
kywdaMD60tpkaN9TqECv30yMyE22Qfm4bSfrwZe8/8a9dLEV8uio5Wovdd2Mi5QnDLrZFaupili8
r2Db8W3393pCf9g1cao3PrI3YP4EpS77DL+e8/y+BI1agzQeSqvaPFO0eUyY9TRpS34UMAL6/vW3
2YTFmdytpB5GeWzI9KjP4v9L9/vmgseLm0X1UaYxjht2YzEBfjeQvpGpx8l80/xbtyYajPRI3rXY
ekh66rw73RpIytZFBy9hgGht08uDcc/RAGbVN9cZNOcx57VzWCYoJcpFTtVhIV4M4h0NIQHYOnof
iCrUlubcWfO4kcr6EYAc/SNPFoj6cO2RWne7cWK7FepdljSwwdGnzy6+5jXT4uoKyHotIIObFlV2
ikie4VXtG6dcI6HbahuXG9rmcwgnBPONV3zXFF0BV4CTnRS7UFtbSpY4U0zQXyBUEIiFNArwcbqD
Eh1vgPzpFdP9x4KUlWAiiHUIJHy9P3RmoOJPHHVXRqeV3UUN8gB0dBY+8MXYA6Sr/6dJd4PwP+Z1
GZAvug3xzzgeMu8SaEjYAM/FCaJUO7JAVj8cxsexWZ7J0RSJQDIhnX/23OELRl35THY+zByQ8mnQ
yQRf3o8dL4RmDgG/wkEwnez7UFgIWg834jOsHC2IvTGK11xIYEZMvNc3JWV16gteE69jdwINNrZF
1VYZG9ovdU6CcshnQE6VZBD/+xsgYtLQ8eOTBLu8eZ0HjKm7UMQ8byFlS3tC7NQuG/y6pCCiy8Pc
LbpIo45+WWOj83X7S77GTdyyM1PL1ft/jATXv9TaBLjhQZT5dywh7f01q0znRo5V2MxmMc6fKriT
bbdW1TYrEc3agC2buwxaUSda9xPtKA1aKG5DJa66r4UMQisgImeK5/9oIsrNJEqY5p8zUgRTEm+4
HcuuKeauL5CVybqZo4nxqjXOxTZEHnPdMFbjZASrx4sdHmCrJHucJgbQn2ssxVGXxFljQkdmZfjR
iyStwodsu5ovyHCXzxPnFUCsbfxU+hHAyf/9MQsStx5rY9i7b5ux79dmYiiswuXxIoVrRKSbQCM9
JVuuWxBie06oyhaMxv1W/B4f7iYbGtzP6Pz6Mtce+SrhgJtMA/wuTUaSvttOMwmNLAIe6aiJA2t3
u+YVRlccEfK1kjvb1CHQe/goygs5JaP3vCmko+WHAosSmO2jyOpzKYMSoD+VbKSmK0OFNxg05sLD
H4z1LFMyx7KbX1dX9uB4VMNWpFeEXFVcA0M6W+a3vh6jOJiQ7Fyu28L3AY7PLXh94Q4CTsjJlP+T
ZoFyAG7KXpOyrftMGboyBY0dieAXyPqBtNklgZI1KIB2N2k8AR7yhemoG0VwfIH74vq4egnZ5CaK
1K/iyNoD1o12j2SbYsFIfy+Y20ZYKVHDjxhNIq05Hls9LwB36VTit7zw4n2pAikCXxMW8jzEJ9Dt
xfnayhxCezHjm/qNK29uV7Hp1OANveNkEx9HLpsV0krEA0YICg4Thp54SVTYtyEHt6ClSXhBSG9T
2M1vIYpO24IezTDuK26XhiMgLUviJm2qrQISA3kBGvoV2d1RawPdPP+MgnJ4t/lHDdtvRmN9Z/SS
+KFIdLoaodYxy4ZXr0Gy0Q7VO+n+5UBR4MlXwyPFWemRnMvS2i+UygJuC8CUAp6mTMzmHqbxPa6n
0WZCpOG4IFol3jGrFjFIV2KXw2wuhu/agLPPKvQejNB8tNLCrorENiEm/guTeU2SKk/JW1HMk60X
WeMHzf/AbQQGTlFqNNMKDdv7GCCYKGBkJxxObKdvFaNscXD8U7KwI4DQl3BmTlZB59y+7Meh79w5
Vv+Wim+j2I0g19/YPpkCmypViCzY3DnKaVhAumGD5nVeIVQ94gRa78p0d2MGto6MCzAiPJk3jmDR
Qm6E6wL9ZcFCzhWEXwCmnWbEOaU3w4gD1eDp7uBrDOdaeiT1WdyjeUpzI4JUhaHE3jEsvKT9FbCN
nl12P/Ke1DUC7skeIJh0U/Xc/hDq6N685WECaWAhp3+XG21mI90c1GbQIwQqbgB/I9AW1PzEVMZN
OzbY0lUENlJcI6tlQU37G7Zbg4D+4BuC4fM7FKSP/WQs9Sv77LqOvdEodl+6BhHHDlU19EHZbp/E
C/3QcXpFUVHjKPVnENGPy34FIM35DbnU2FoDKYgJXfvooQ5YFlUpZ8kfMZSh8Oetz/yfx8gMrqwz
0WUdijGFSjqfpkjUsHHoThFrBmbs381cTpSJZmP2/jAlFq8h3gi7QznhHDz/hAD4Z7fyatjongw9
qXdmLOBUVOXIhk9b3S/GajBnKtvx0ClNYpg4GvMp5j16tLTBvvg8RxcY3xwsh2LrToUPp7l8DNgI
wfXylqThKatcXyQad08XbCRn70E3H2B7tuhOlnW8LoP/qLMpzoNjgFXw/FSFe0yJe3e9aUhWMMnh
a9XS3YLCZ7wPJ0L0tWXi6ngqV6+WWF5xPuY14szdpW+zXjdAGqsIgtBy4Zqi/gsl2qgEQEMKbxix
PdaPoZi2Z7sNhcn+l+w1D9Z63r7xVPbDOFKgwcQeL7R33pEDa7n4MNpno/EOESqCIY2Th48Dpa6K
vtiv0qRpJV0I7u/NJ8spLdIBgAhzon1/bGnDBUO9RC2CBDPO9kuV25/DxFDWSsJ/FUkXcphL5tJo
010mRUJWfSYgeUwJSIG+OAGCiIsxq1fsCBA8ibnDDiq3G9Zbdb9jE1Gr/aIHT459x951PN5atJEU
MhjTKUBM9PKLoREtnNfzSO763bufpN4y8vMQoQpoaFgKalwd73pkXpKZ5pgjJR/Ay29jl+PjB0oy
efJD1n7IafsQBX6qH8pneHkE5xYrCe+EDCXSk4s6hB5EV1O4on4/aQyJ94t2SA8j5vGnYyvQe7t0
quBYYnzE027T4K2yUuWR2u51mY5h0NQyMB3QtdDCHm6xViq3AoqJXGruP8xEW/524pOOZgcSgTQG
EZbFivGE85BQGiAEkF5T7YIBaOwU/+Orb4rgJzk9TlQHIWBIqoNe4J52BYqd0sZeiK80QYaW6YKS
i0Gn2DJ0ka9PboPQ4PBa3baW7YRKk8sPQM3oYDCu+DWyGqj33kcR9mZoD8WWeau5/JATSoo1QUHM
Mckn396AjIiKI5iSQ/oXSJ0Lq6rh7ezuCaH5tTbbk7WX3SqLFR7WD37uNGtupR2oxtQBrPo2a5Av
gpKPGqW1SStDxgjYAiTdgdWFVyob+Ezt1lxQklY29k8IzXmj1UObJpL+RxTt9LnhKH2Pcu0hDuuo
QfvLbx2p75kaQM9yKLb06E8O0JQeQL8CQJR9caSopCxxiFKCfLnFN56qRZ/rrRNxw4LjakSLNNRQ
LUywWy/vqr63GDiKLNa3MBV9fx0mNVRAWINfmCRQImrXKQrAOsSf0ioa+5oUUt1bEAaqV3VZQeFp
6Zo/k/iVLtOgLWhNWTDfzdoUweP/QQ8yf9QiJH2bhy/99VjIJimJpXk+RXrmfyKlVunfzd6xS/x5
pQqtcvE4hTUdAr5tvizvtP1IVJJy73B1LMwrjSLc6KfKVb/+jPGvjxRQdchjifhU8+RrizyRAtix
lm0clMzgQYzVuDyoYUsm1CdMnQk/NkFpeuQuublRddVvKPvY+ESoXRWBG93lt4ZLKJmqYtKe832v
0/zqYanoFwSwYmYoyis0m9K8zhucao2X2D6wmtYkL/eEUOrE2lv2r4xSElBt+gPFcFrmxsYDrDin
itoZ2m+weYf7SOnxei6bce1Lz2hr+e+flsYIHy1MOEieM1qd2gjmNbeX8D3EBzC9mmfJ6cEXU8oR
86uoOse2dsCVq0lYY3c63947pgRNsfEztJ647C1+ZzC4oO9xtCAgKDtApULT/03FdljQh1h/Y3X8
9ppC/8OsRcsFZJX+CEx0311pNgCfUec7X9v9EEZEKy7bJFijSs2bqvcAHue4FgjV5v+L1dq3b7v/
kLYWXHKZK4JzXxZe9sOspMjL2y7Jny3mRWhBg6clTPO6FPWu/nO0jZ6l9QMf9EreO6r48E5HF4EA
dBrrX2798iZ7+5wnX54QC33eLxxXEah7afDAv28AnhaY4nQSvFgng+DGwVnJLP2m+Kpe3TIe6tNC
xHYzLB2ddf2ejWOviLcvFsxQsMjlgME=
`pragma protect end_protected
