// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LFHbEr2djhdkRk4AiUYv4ajfiy+fF+8vjVn1Kz92qOk2tqz6EvmjR38K5A8lNGHmnKPRXULquQU0
fftPUGWYrsFGfz06x1hoLC4i094eAuokNsKyCHVJuxYUeocetpXg1aCOfRJV9lTlMUOmDf/tkg/w
AOV6tnA0GF1AWfE2uYy8zajbysBb4pUEYr03KPNUpnEhAnWBW/L+7YFYCCNZYR/zZCwGLyCGzRX6
Uu9a225ihEOyxt8zQPar4ZMbg5W7EdB4HPlVo6cMtymmgrpj1wnw8yWZkZoOEfQLH+KGUQIvP+vS
DWFnguSVC4KEVQt2XQd+1Y1jxSPhluvjBHvPZA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 18256)
AiOyH6aJpQhwNNIzjfzdnpHl7xzEbIYvI3xhedLdIAQGJGAujIvW1gOVOnwovAk9qPgkEyux6HKq
J1vp23Bu3EDb0BmMLmdGbeUmVEeN1uHoqp+jInvjL2ttPltbtZzxZHa9tJfXrFuT5RPHHgz7KWtt
fS3dE2zHwaQSESt+qQZvDL7qXn/yvjGRVTjy7BbwUmewyvWe4eoYPKNqz0RlQ3VwQjN4eCBpHLut
4PjCb551YeK8RkVustu4mu/pVNlmpaqmFVn/xMPRweYO6vtq37uKHNK0Op4BiPV2z0n75zrltwkd
UcocVVFZPC3iNDUkpYOAtZxwB0aXyMx1YXk+MzZjpGrlLzVHC0hKPAe8OgHXtFDnrrHwPRWfiX4S
R3uvqCbYqP2Dr+BwuP74ECUdF7e6dNVYdPLHVguYBz0Va9oK2AcHrILX09LVShfCwn3s+x8awfrN
sqkWDJB9+FKulfItbjAlDEMyZa/uB73yhEFwBBmh3HAUCr+nC+NEeI03AVU3YJQFxv9i+Ei/0n7p
iPSvVdVZwRoPpvGOo3+yTlj8lXOKlm42T9BEB3ZfSNg/DkwSGRxmJR5k94fnd0wbpu2I/N2fBAOA
kS3B7PX175mvEyb6201+e+MOUwGGa4prSKIUQh2jCaEjvA5n/wgJ11+nK5a2lTG2ftHNMAboJIqw
T0RPx9lZxYXd8xYsRjVmvo4SoDCFPMahJAkQh4Jgff1nxuw6mW/3saRS0wmXD3gAJ1HdMLQWPik5
OqbJ2uogJb/H+bI7V7ZJ8/rqikhOTqmRtAEiArcJu4Ug/mkeoIziKmrqT+MQXrXE1xoHkJpoyhhI
1O75eFS2uSD7NrKXkW4Ear0rNvQb2sECF15mJ/jlBDCCv7fNzpYn0lSOsmBO9uA3wgJZpvzt45mZ
HmQ/9tL9YRBZvfv0uaixmgTFdrmLD7AAvvSfUPtwlYNz2nbvMqxPEnIk9Yph5gTyI3WB3I/EDohf
OTjXxVBiaU2ghtzwLIfQKY45jY9HIE2hv5BJ1o+aKA0anzoithHxw4H33IjqXi6OR0POBRVf5t+M
BiVzz+26Pccei3+c1e2bT/wSpq72CyoenSOoaAhPGSTvPAeHFJlAbPNB31kuc5sUUTrnLEJ0bByB
ZbBEd6hhSG+hnGLvoOjh05E/aGWPNSJmrSWhKHGj7ZObTDTvXTWj+GIoNcqwkZujQc6LJA+zF7e4
2ZwJXyYZWDjmfzPx9XP8FDk7vnJZSgv1UIWHyqVXnIgyb0u52bAgb2qms4TSKaq40dp5MeFRV6VY
tUUwVsvUdFCQmbrtomUkdbLTEA5RzL/dBWe05Wsr6XYHJDgAPhKN22A0eSaVOj+yriN0/LKajXaE
b4zihf7HsQFaHC1FhxxowH46K9C+KiVJqUByAvodLf50NwBOb1SDsVbmmfbOMdJHeCNnJcD+NpVd
S3fE/9rlNl2HJxs8W4LYZp7Hq71Wot4UYLVFgU7RvbJYVmY80kccrGpq7By8I/pHA4aL0V94aHbv
HYLYEsIHCyO3TZnGYxhtu9JxQJKIeRTJ0mGt8h0kk3XXGJcjpL8ENguIwDGtahjW/hLUJjj5gSF0
csqFOp5M2YKEkvlqpqr1TXJOermaiY4N1r6UZkAb6g4VFV7Fa5yebgNEHvuiSQeDe70oIS6w7HlM
xRQMxFREirG1ByeTIZIYBjn4CudTyotSsFqR9N69MeanF3uNZ4z4sMc78jS3CfuyaTrAKruAbh//
yd0kejtO5VUEMqr3URlAQ+VUEoxuzNjlhXU81fvl7kkwUc4dSPyMCP0ZmOMs995vlAAEjx1OkRxE
fv/szRmytU8XEI6pWqivw2l8ELyDLMbDxLRThtfkic2Mcpr/ovKC+QebOrFFiNjeMyCoUBYkPrUE
zfx90EIiFBCw3BpbmcLvR0Wax1xt3zxg/VONtFSfaFc7Tphbq/fNjf/qXkTfvXftvr680Usydbtv
vXDJg8VySwkMwVmAzWmARhmcn85/KmURC8PXSj9GS1WLUFeV+MgnbdTShRbbMqsuJzi55S2OBF/l
N0nvmV/h3AUkA3SspcF1G8YKh8eC7DY1GLliGOkWuHiJvq8vK4Ycu3W1/XBV9v/MilbcLijasRsf
IBrWu+80EV8bICM3zfLvma/iV7hZ+RxAjtCtNmZjGQrG1ijLeD3Jk5arRsYHGGM3oab6jR8EJFOl
8sYTZkPTKmgrcwpgkuzWXA2i+8Yy5BzBaf8chWc2aG6t1PADBHAgVBdr2KzVFIG9WpWPBZ4S0hSg
4p4Hi9Ihx+xcxZxac03Njiij6Tz5mV6m5s4Abzu+ViGWcLg0TYYE6P0GcCTeicjDMunXa1Yi2ngy
7y6SXL2iojRLiC0dx4dD4HRoiIqrqEkhIoo1q9fC40TeYeNnM3h71j/qqIrZr9A/AAH1yL/nRRKG
UBPkkWPjUI4Gqq+qiZnZzOBxtUAlWNYgZY2vE5cEAItX7UgWUTvY960pbGsTjOkQazZWwMcHeyOV
tiwNtojD38FfSOz+fm7AhQ5Y1ibLmFdP0DL4QiaQiRL3h+Nc1uRwhWboXlTFzMw9zCTxsKrOkqVt
zpFgx9W4yTEkjZIBI8dx5az2AUqQM9gvL0oYCiaZeTwAvJQu/oIAGXZ4o/hPdCzRRTT1zxtSNyPY
v5GQPXGRdqsugcWDcGqnZyL/JEXrz8DqZrpX3AHE8VwGRVMsqr5Y6011B3BFjKvxXuJBPtjjCg5C
vGbqe5UE29PzkuX0hFy4rTXtPZSHmEM169lGfB1DaOv9dg532lwwc7EcEOlRNZFbu1sgkIHGBYIa
vm6IfxS4AwJ11HgqBRQtwdt0JTLQeNWp/R9uLnFXwTXa7ICIlU3v1+e13SXWRfUQ0li41fgRFyRM
vojvEysTmC3UXZR7XU56zCtBWH7LsdAhu/2bhJ9+PK/ZmK6X+4Dh6yJrhfqaHhfv1etq3I8X/T3R
vIgPMyKXX45tbNp+lKlV8DBQz+sA0yR5QaQw8Jp/6/MDf+/UamIA89+Jdklk4vVf1MCFaTzPpD4+
NRQFhM2DA0s6EBfhk0IcO6Ujiph4jAltwMNGWmqsOjHqN4U8UNbUCYG1VHIJosra7CV2J35qGCaw
6Pz8BSLgZicIdW8G497K74kP0uxs75CTQCYJqouPe8+NtsXIWEgFFFiYiGRgGUd1E+2UiyBTPa1u
W451XnH5ucGQdhpVjsr45wC/MSvjeUrb+qA2+dXsn3G6aqvnbtL84Hie+3cJq49LXncHaFcH0LKP
k1H8pQoUo8P6Np8h+3diZ9Abq/XDV9+30YMzC952O76wPC2hCJi1CsVOS7fAU5n7NmrCOG4I/w4d
8GU+91dzZgQb+1mCjBFKzPBpjZHSHgSTfiPuByXij3tOJSgnKyegGnvpkTIhF+lHz+chih2mq1ZK
On89MAcPqkUAS2ygKHWja6FiqKmvWjjx9hoc07u/FF4Eq0HLOvTRFZZNXuH/ZOAdWjB4y6KGtnp2
C8xmFZlATPZhWBssIZgN6BdFwJ3ySu+NG9nPM8BbOrUGZrq7eVJ8jjYQ31uFE7Umn1x5dAdInUM3
qFW7COH5RcicyQe1X6Je+vCv9xqOy6ejsv9KisVrFQTMPRtU0M5ByDfPCDPNQhgpzwEhhqzsX9yT
SYaKE2BXNNw8tb1WuXh2Pwf8qTeDo/ujQMPeucFcY8KhwqQkLOMF7vgUFVJha2h+ISv2UKncDxMg
cfVWh/aQb5AIQo1jFYWW2TpDKKC7BZFjxe1XE1vq/gp6VnseF7E+VcCwmGI3kymyUL58af/EsuuZ
WuX0D4ek8arRf1EK/1eb/0hM0Zvn+c5UjWIqNLPaq99VeSWt/vzZMhAUD0ecDrphMKvOq57AbPFY
mptt52mR9RO+2Pc/kAwJUVM1wTG3DIbTf7P/Ke7Z76W4ZQzzDkEOcA2fpVepUzVs1NB+4OVZ9LRi
cgjBeMPNFt+ms5V6n7eIv7bwUPZOvauzAX/jC7LRYR5EPc8K3btkPdDS/wgrjWrFk3PPgm7Km2fp
pECnle+RH8BLUNuXPwgZ737GNhrnkyfqr/RAllCIXqzAltr9hg0EbZf8KhdDRbQRYe64Gq6of3wB
G+hOc4FY6fSVO0ZDKijxPSkzkDWljOQpBukF0rit/4OXG8Ynv3GiHBzBI62R7WO/obZIuEA2ubHL
foAxiB5tEuaYXe513XhHEypIN6BMGmvdmfY3mZ4iXKnWO2lZyYy8VT0riqXq3k4/wx6LeAJV9FV1
IWcDJYp62lMldqqz7xv0NMrHLQlsIgZa6F/0S9SfYSwYGlze23AZwUA88pYeMK2XYlUzfRpJTqX9
/nR1W7cohG6jXp9JdUYqbgvutE74lwrW7mQ8ADhkOsMytDp8vwxoMnX8PqAaaDRLxSFlGm0e5nDg
DQW0okWxmUSY1GeSUq2CGK3M+POdvBe0NF/WMOaCIkFQrfxDzH1A8To1UGf86emhS7mRBHKkAjyb
EB0hOBl/TAvQIfRg3S/o1vmoLRyRxHwsqxNbNCqv64EfO4vwz3IDPDhibSJ1V9KRafeXk/OaAEEt
8B0G7oC/uHf6ru/HSiqD+6kM4T/m6ZHCjPZ3mtbOWMvLL1hHuuD+nzWpZ7dRVneQghGXfFaDXDK4
B/haXvhMw9aKFCAfHKpf7JI5j0p/gFUReImKArkaqqNPE86ppVty2jIJWCl7Ty9Vb1XBnUfcLxWL
ap2Gk2TmeG0jS5Y7t3C2raUTGsBS7qJEYxXgOcI+E1/pqKqhnmwQKEvyYeRyfcahhoVgPsVnhqb5
aOCDD5hohYcUw3sEz6yPiKU8N7eH+VkoOQCmtlxNO/zy2hy67OvtwoSrrqOaW4QxJmq0dIjNFuPb
TDpHgW82wolORESA2qZ30q7p25wpP702bXozHZkzIx4gjn0/i+FOEkP5PrGlys/Brk9QVvpTMkLD
qQnR6ydIcvFq3pr4zuRl777zDh8Q7rR2xdc7qRB5S9XiEaxigXn8qGzEBoWhT5MW4JRhnETnVktr
3fErtPhxSWo8sYLGYUv5YR1i3nwdCHasxcBEQtWlLW8YK0LyoXmfBS9Kk6+5GP/4aOH0mQkdmtiy
w2n+v5JSNn/+hBKXfTJlQN1VJm4hLZh9ULl3K/k+vsHOezdm915jUJ4+9+35ma0VIB4WXaF8oYFK
CxbmAf9Mc4hIJD+tmAlhRyd/bttUtwNSl/uUq6CiX7dcKhhNBkeDzS6nn97HZBWCuAYl6A66P5u6
fbBRUq+H8Jyi+a2bc8/zGxpgiFKNQr7ehw6/YB++7LREGXgkCz6RcVG4yCTpH/zRQliYAbJMKbNX
vyHxtJEyIkojMeaLmPj0DQfNELRNAbIfaMwY7G+DbvWQwsKGShUg8h5eOOPFD1oDO0XOpUGREtwy
YvLglDCBik1hWmxh/3tsERYZVOtvQxYIqjS+os3+kcjMKnxIWWmMVdTnv/hEiVPmWfmmtUnMhQ+2
Oxz638Lvg0jwYnuhrEADBwPVp2AQemZrFcUIdaSpjtWPTP3UA+W9C1dbrn7IGuDdJohAh0kojuGw
PADE2b5BnG4j+MEqvinb12RyxG7r9Tty+zQ8VYCK/x99K7Nyjiba3qOv/oQTfp1WRC4awcOe3V/g
uDmj40cYaGoOpSUHvGtfkuMDTvM7S/wPXHM6bLu6Vi7pi7VWLF8D5nnBuFWb2l3pUiyOatlnfm+r
oohXjkYZO7nlr1053a3sLSCUxPmPFIgUX0a8ofHBSTY47ak7n2Tl9y4izxGha1ScwuEf5PEoDnY2
JncVAmmb6b+WDTqp0/5a+9jDgmzUperba6yediZpW+5RDBA+oIg99lUaYOVY0uy2r2qO8rqDw5tp
09OAQm1GaIlkcH2pzGux5jY3UVYCMSD4tycUVpP7m8bszlUIh2zgg6KxzygvVkC+uqlOpX79QYk4
1qrVuojKX51PUru6AGNCGS1cGB7kHIVYHtL4ttskPg7QfdQaV0Kf+19/ggshRNdqJSsUhZpVIrOF
M8YCPuf0RtH0AwTmtyjlwuVkTCayCt3cj84AYu9vjdpbsjqhr1+SJ6TLvF16aUgIYDdyErgiZWrS
4p1rTCpxK0xQNn4TlLMcTpW6AddlVJYHosN7KtupGaTCysJcMXBR9J8LCZeSXcXOUOsm0hCIgAQv
Hf1QO5mHdN6mErQPpuZML1I2vDXS9ClBFJelqGG+PvNDAlifJRS81cjue9+2uyLMSMNrALWIOXn9
RV7dvCwfCHrRw2mFjtq10ZSjMul4l89JwE5fUzYjgEMSZHwoR4yXtHgLZCiB2JBQp1mlcGH7WxZt
XWAiKGkCdTtQlGTKQRo/I+OQZgOwLTBxYKbRrjCiGBTM8FCz7dVcHgYM7NIRgxEZyK66aTbhk54Z
FEDr9VhAxUl5hPwDLlQDP/SLC21pWOxbjtkMtE6h419YhpuWOcPXWsvQtDTiLXXxDIbw6WHdLXT4
0u9tAk/6x7P9Tw/8yPwQLlpAxNLdRJ7nlF8oPnjeAtzY5eqEi66Beg7tQgjFHFhEPMokw7JBPrfW
HS/XyURzf+te3VfQTSCb+btMiOn2skKH+zvEdVLUgrMWDFJie58wkwKQUU7I1zuWEHAtf5JikUSi
3DyojfZxq6wKdi8Vr5H0AJT8n4S4WLthd2hNxnHg08Vmu3eQPsqZZnKOWn3wVvCvsFRoFD8vRhq+
29cD4A8fwmd/XNCBA06BYwTBvEx/wBKFGDbXB9ONSebNd3oUrDfOs/5cOUjoFWRq7OHD18lKzna6
sM4l4jDohhiBrCC6L3SrpgnmdKiy/AAjC2XicAniDVZSeTFPfkkHdj7jDsE0VXB/XC2+PxitenmP
Qk7ZuKc5bm5DWBoZt2U31Bl1pTy9QROMUvUzkAlBqOm535A4T3T/pHT8clJ12Yaj9RYw7/5NzdkR
TUxvJLcNFXgL/W2f5NMZxdrltW3V0PLndRhxAn55hYpDuK/73ppyYYLAwBNMrY9Oxqs5suAu45b2
aqGssno64DqMeJTtGIyOslGic/ky6DgGZTkq3xQCQ/tMLBSkx0yf4NYbyfGC9LY+33FeG6n04BJ6
Ts0hXWEh+np5diLvd400AUs16nlWWApfz7KB9EYN5WE6U2GqgC65+YpO89/jqCSdc17Mac0P501D
lYRTXwzQ9ZvGSRJ9s7sWvHi2GFLwdBxMbyBO2QUfpvV9Krw3373RYQmk99xJjGosJDdtHQELsl0p
0Q27M18D9mc1RjucLmMgtYF9wVIGGUcKOSigD3KwwLIaChICLK1b/towXKXgvfi0I+iBPjpL87P5
lrSGa2Z/DPXetqk4alSOBKiVqJfMgO+YdnLDtvD5iBLQxUgoU19+hMoHhPj65D6egGi1JTAxsJ8M
u/67bAcMcCHhuAON6pvf16uAL9wNTvDl/ITwJg+YNUmR7K1rtTD3QuoN8FnTrgxyewR445WzVAL/
lLaPrkKvRl5siltUGy/TWjxAAAHg4F7siX0LoRU/n5WZKDIl2n5eTHYmlrDgs8dP5rjG6UH99zaA
Yhs5lxZ2wRT4jfGjU+asp5b1+X+WtjtTUDAJHveoUCs79RmCJp2/0+KBnSTOG0h9GAIy7rKGjIWq
9ygp+RIsjXmDHEOeaenJaAIcXYIFXs/QKGwHzg6F6ps7163SA8oSU3+pSW+JDb1wtCfPwliZdsua
7OKDNBkEfekKqb+rqyoG9mVCwLQOKyfCPvRPsEs0luwgK+Td0yB3okU7t43gJmkfNkD2nMVvxXhv
u9dtIV/RywsGSZuk4spC1oqR6IYpCvBG3b45zIM620K+c2Bs3jp3K6cwOqWXcw8/eILqRl+ibH5o
KX1KnnOYJMqhaQVKuL/R/OXcHGgTFdxR0tXofdInPZLUCAhI4xf+lzN9YDL+QoTPgg4gyKLX+Gg6
StCvS0ZBVQ4/n2CwsqWs8udMMn+pmSAWY02gFOUZcz9nBiafpgjyQNqrt+xdfe2gs3jfVzJHKxrU
Qqtv+B3eNXOWvba1/Jxfh/2tvLad6jnQRmn1n4g/32MMHlspwxX2LqauN5O1E9ZnjPeoEuTd2Yqc
bze4VSV0hl896DQBF4GpGeFhPo9FppKwspKCXRc8UHPnLRG2EAOJaiuloOv54gIeOdZXN5ED31Vf
1l7vf4HHfzihIteYovbv8KQCVinWeYhgGhqxM8cj4KNxBl/aTxpsTTFQvlyhsqN4CLwHlCnQKHIF
mEpFSZwlE+6vq+/yw17GvjEbbC3WSkOuN5kDqRl94Ztw52+3GoONGpitUwVgnNsc07sgdqRqunSf
yhvirl6MLhrPR/oLDFCeSB/TV4f3+TQRmLBrPOMQf69PsLRLE/pzKjoHYI5zo9smpNQISGQp4DXJ
PU4Ka0TvZGQ5fVR2HGXDAXfEudMcJgb6POfZSrMXe+iv0tSgFysAT79VUWl/PudV/9qj4XdiDbqf
YRRQU+zyBunuZpWjD8ek1Z6HTn/rOCYKLFX4x1gChkIcK9f0Z14TZx+eNResRYZEOMGc/kB7vI+o
ioz0DJCxqhEo9KDmcYJ4dC8T8Ihs1nhducG6Q3PhKmQdm2+6miZPTxiaUwy3FQ/ZNr4SQ702DfEm
0bAZR29YAJyfuueos69UrcvL8i6US+4rjrX5dPuDPrhLDhitBzU1BXZFKm9EoKsjiMPWCOGsXL3y
1Pzmhs4/E/pudCyldHld2cC7orWjdgOq7JbGaNTKOnQ1Y2LeHwzlJQxFI/kgvNaT8Tu3TTnP/Yxz
vuGOhKnZvixnDumtUKZIrWc7NfAVW06obS9b3hzfeo6NXfLXMUL6OTDQ9MIKd99+6/I4LfhynJ2m
me7dxO3n5Rc3nRxb2og4ziYgmv131MQ9HmG3WPX+czbXs8hbMIyJC1fdbg/YXy4EtQDev7AY1D5t
H1P9pmyvpVi/UDtZ7cpq2N98kIfBaQ/+ZisItqn/1flQWbKzk7hYMQqUXGW2GBwFYzAjsVnPinKw
AsfSLeGt269lbER9EdQyE2VeW3i1wZiNnL5d13bX5jbIE+WqLjnWvqkfiiYwSCkLHM8tN+o6aSf4
1SaAj5nBHno2kqZHNcY5tryPEx4uZZBIbhARGGhPlckLtXVvj3BD7tIyB3GMFDa8xPqmTeppjdrW
mINI5Elxs7y2eD0WkfjdDVcQ7C969FdvMMg86tJiy+QkwIMTMuFriNSPbJIkgizlkZ9x7wwuVmxW
kUNbkI/EQz2/BWGlgVDb6mvozxJMTWnJtsK/STyOgGOKc0klhMwhmPYQO41q/LfIjayb0LevQlCB
+B3pb4kU+polH5ulLx28c+DEz7SqkUo9kUgHbrFVNu9hxhqHtBF3MTbES7zPprrfvSpKUHMKJHOT
0j6lJ3SHVBlTIpHVT2aWdSqcSuTqlSJl0Ya9dVx7wDdspLLWoi4mXbkm1XgGXSBwrmeaPAW9GtQr
oxiGBthXPjyyfhapn/J+8p+Ig5UN4aB8jjb5QIOHbVI5izyCz3LzZfaxcWRrb/3ALmQoGvchfYwA
LUov4Y4FpxGQwBzTJIHg/g2I1uIB5WpK1kCP21pxGsBgDR/qU24SB4uw+JCPzaaP2kkfwAP5gK3j
DLJfjOQmN81U4NU2PnWA/IVdzmayMs+7hTr1qjMJHg/hs3e6/v9w3GukTbsURva9WXbTwPM1PH1u
lHS39VIIlOQQCduJdkoo3W+Ac9/VESp+1ofIgwc93k2VULf9FIEFqILKKRo34N8QE0r8cVMjPstg
NKjprj4mVgRGsIo+u/rby94CCcq+phGydgz9J8jc+AB0DN12aFKAHcsPLqLZ2H43W8hNuSHWif0w
wQkKvgoqRQOnye81lPYTuRm1+aLnwMgzSI5iGRzszl41OvfXEKmlQZ+g8RTeaHw7WgjKyJvmJODa
2zYAkTb15LPgytxr6y1qW9Lt3v1Rvl50YV/t7MoSrP4AgyQG2X1yR82fSFZgmoyccIAW191YR4gH
MCkdndYfjYCLTJnNKBHvYkBYWIux7m8yNgIsNUt2lzm5AN3Udjvu12FAlt1gIM8QWZrAH/uxuHX4
t9G2GANRLaET0a7JlYQ/QNwasMQEHa306UEQUBAMbveHne9ycnNySZ/eDpW0pzpKsTE0s06aWral
HmfmNjtJrjqSiSwCyM/vEWj8OkIPcxM1OfCX/eJkhWWupXy3988ve3CpD+J9E4S1V0ZVfeaE15Zt
9csMKaJDfKZJ98FGUiHx4Itrzf2OMoqtselKi7s6H1maBTi6HcyA6hfBzHQgcyVld3XlHyc8f7e/
MX5SzL0gg4a23mkzD3LkkgJmDz5eG7CNdvOeItUJ3GUQ31AZcqzCG4L5ln91VLLOPOsK8emx8ZGg
IiPtqNTu1J+iKZpNhzCIeaXEkZP/qYmWXRRYZr5T9kHVGeDd1u3H9z5P/dZG54WZkZmmC7Kww/IR
6sR5P+hQPyhBh+RI6bS992fiEf6AB0v8uUxn/fszGP8LEHeueJlKbpEDPsEGgSh6ZFIYNckO3vDA
cDGVglUrpCT5Gmc3uKD2GWylp7+FomiThJldYIFXrbcrOmRQ/cwCyrbP4INwFaLoe4xpQ/PmLMYt
pNW3kHlHoashUS63NWaCEhCxw1CoUi/porkrISsRNf82XCCI4h1vv2r+hiGHAuGZAXOQuJwlhsWO
aTbTZom1qIhE1Tqxol+qbzYTBZWHodmXfY4At5dtA4kLfLIvNRXiv1OVAeY6YYitsBQOygpBPus3
ySO2QbNSDa8cEuEv2pZLRW2JqCGvC8nmZN2ubBCQ3zEv7b+CJG4ZAz2+zIj59kXBk6yFLfMoBIYH
OQ50hZKQGSOP+KoO2d4t3MPKmxiD7tkwrIODwMMSHK+blOEH0SxJEupW3UxlQ3+8YGKKjs5SCoD5
7Ojv6zBjOj9yJ5HUNyzFHoGmCNeCy236qLIzenjldQh28xUZ/DJhao91xgGJXT7+ZJ/v3f8C7jx7
BD9yx2QrbkEMozTduXRk0PcTd5evegSzQlhSJXl46FhCLZ81V85JHQTU9O0qCKl45hFqYBxth9ti
6uMXvjc1eU+gNU8zFfCgdxYgLFzVEd2xsV6pNqiJUJoumwE6coS7zpW5Aff8/ZIjCyHYRTPOw2sx
IAG8VNduFcvC4amMhmdTHnUaWW5NNGMA2/b/7xO2J+Ji9/xxSWj84O5dYX2re08KRwyY+kebEG2i
38xNhGbl3sCiurnGzfKWckujewdEtYOJqQ+f4U1wcJ+8uv+dW0/XKDBiaLv194vb/8RiSR177FUw
tKnav32mJi3UDjmQUWiKw29LIn6/nC53ZDDwMxFWkjNIwdSgpz6Ob0Bsina9/jngTUUXMzAJ/oZY
izJHiYCusk8ItqEXihIbHS6MF4KrSf4NgaHckv2qbls8P6wu8qsMMKuGdw0DTOfUorwdkBlgSK8D
ezjUKNrlZiLAWayO8hzGXUcpEmaoRiv9F+fSiNC7imPHCzfbN84ZzHHpi9+CULGPnl3a4ja42sNI
EARNJXoIAvgYgcTfoXOGVfuaIOw34GQaW7tvvdt1XGZh8xak63ohqSF02ekeRg6pUcAa9y6rbsk4
fhu2IDFvBabSeyFkOowH1nnWUNLPMmNUxUSPliZKR0p3OMr+DvecMiHeuNLeO7cGTnFnndzWCHtk
WRVu/fPdXSF1wYBX69T6DIMmP0cxsxZNG6W11xj1jD3spKZ4mTOAZ/nvvsus3ysFypOGNEAm4J9h
WU6m/rbok2dUOTKacRv5EmOhPSDeu1phfDegd+ob4BDVkCKdfhbt7n1MZUDPcOcUA+kM+GccqeP4
G3MTPRksWxzN7eCmf1RdUG0aNFFknlUlUGNqBE/wmS8Ducz4osCML5QgPiqgi+Lu4ud2fzrCD/v+
yOzKEBMepi6zrhEB9I6D7uLgqmH60aBaG/PHqy0rp8KXUslkKGTfnPtlmU9y7vmo0tkHqCFhKMx1
ttd9l4oWCJrRcJJCswpPAXKBKQO5CzjIXPaDl3Nsl+QNlYM6FGsPAMXl+ClbxRH0J8Zp9U6fvV87
MloY0uDHngjqY0PZ1fz3JLK+aTrFUembXXniKjeU32mU1p+4jRBrNqv5eSTKxHMNz42NsnzGK0DT
sU/gcMPzBVjO0hYfN4KaTBNcUb/YOY84odkEuGULEK+uJM8XoA1HFdsUy3yGUbehst23JAJJGTFw
8MN1GB6x1txSbrMouGAlIZ0mzrJV/xwzeiAyHtjQVIHBEX0sXCstskQi/SjN2gSuEjlyZthbXXQc
j18SWlJs+k7PGejjvaQS8H8Vl8O9o9KMuhUN/yVw26r150xGrsYAKdJ+2JHMAiJEohjk8YRNLwfs
vPf0cu2Cs2L9s43MGQ0PmEtG/PeYJSBqtD7xwDcYjdVosWrucC9iVpBbX2R40rd2QCcKHJkoLD8C
PWnQEQTSagq4nemsrzWPQcMYcFpL621xamfI1BhNnS1XQxcfWf5OcKV1/DpRxofJvhycZtccOzTD
b/j6WqmVt4dIUEQ6kmXL/tNouuvHeM5H1ue147U4iQfOOBgAZUFi0s5yETqW0W76lfTN1y02ossE
q9k5jcjLDafmWJYpjh9B6p8edioT4N/zCeuc2gr1KilimvH2IuI0zfmGPcqp18wxUIPUIXVsUobY
6VpbZEQwRXU8q5AfXcQ+RF2BJvoAzLtIMA14F73SRy9AnIZAht+tIvfyXz8MqEcVeFyyV+8rVV3Y
deH32g8a1pR6CJTgL62rmwZkA+SqROU7popwaQEqtMps+TG7GCVHAGlznkhwQWayARxGcecpMcpw
Zn+tUmqZvmmYxY5aemn4H81d7irdYf273KgfJxA2/Kk0vCvyRbsAspfLgQHL/Lk5JXbXFVVxlRt+
VcW5tjZh3+0JQL1KMw+LlQ2OnTFYq2J6ZaKpMq+Dx8BiHDNkjWjKfwFsCw+ciqGSKDU/4jckzijr
YonWTD7SjansAUmPsVwpeKKoFEgb1/qAWklSMWE63ORibri1IZdkBZNaIBTJGa1u44Qgra/eWXTj
5MUhTJmQaZx/JDSCQ4nPngZq9D11gMsWrMwnxq0qzRfEAdWMVgpsgXLQKXTBAQW+58LjDP3sWPra
/y3I5dVfxM1mZiTxEwaomOuWN8qK/EeUaj8MWopNrxySs4a2sSwOF+hwuf4v7nH+aMUokpFDisgz
FBas4lqwafE6HLXL0wHnwUearHydfDFTTu3kKWFwN2PAy9vafNpDLMm7izbSBB9t3WXQRYZwCrG9
hVjsFxNkPnPBC5eOEgAatG5gy+wgfM6Ogp5m0oTwO7BvM4iaNvemOIykdNuUqPvmdBuK1uFmHBqS
Sck9PYinEPwtWml3UiFTO3mju4Z7SFHcg0WxXONtI1ccHzQYV9z192cMsFRg0Be+/UV/WK50kxgs
9a9q6RfZGo7FVUkh3LC6osPextLY/08N48kjL4yAIpvJZIVR1Xu4yA7uAi5dEBZJdEPxMChsxuGt
rgZ6mQPYtjcKRqCXIDkeKfSJCzRVCAokreHtwmh/RIEKKfXcETv1Nj7W4SWtdFHr5Lif6segBC2j
nCASc092KIw1G0nwtnQcF+rZ4deJtNAlOTLpXzfmVmJwxCJPphOqEAGWtxoG4k0LDz31pzk+Rz5B
JNXcOYOGL2f/Dw+NnDV7lt8H/95cTMO/rEpckTQFaXOTne7B6rpHRgnMFXiD+AP4Km0pXjd2hmkG
SJnG1Bz0MR3PSIOPGsnWJ3dcubzLr29Vxqylsp+yB+XknCTJReXb2GdKi3oUcF0VsUntlyaG7o0v
0AJzXMNFt8OfIscTDSX1DH1hNnWsq33HRenVipA9LJ91YaP1cOvkmbyPXx9Sdv0ODwkfqpSszJyC
+Op2d2l6Tz2AJyHltNP6zZzFRIEGNa6AbWWIm8pflsge0VYca1USIPZDkEd6qWWGp0gGWUQELFAG
cwSvm/zwmOlg0Ak2DGbBL0OjR3GRXx3KPZy46oAIOIJvHfaM4f+Uo2PztAtBGSYv4yGYzJjEC+Tx
mFTnlNa/nPKyWhSt2gIjsDt0fabWrEUJBf5q0K7xdJZWNJBR95Lv+Gve1K/nnQZvZVqjXo/yl89T
0v4qJHiq8U4hV7wSnKnWtpYOIkCtOG2Si2laeNfAJO8f/U0mdKzUqBqHxg1LQvu2vpyHI0ZFp3mF
Mdm+ls2XGzhhkkUMi5KV2sCYMlDfblZ9ApJdMwK77bsmMbPF42w5NzuMzzi06KcTpsFCmYZDnNd3
VtC4jj0zU9H1yYBv5HQQ/JXzjZ7IsJGbHV+AjaH4oVGDg7H5u0TekkwRLcfBRbi2efwbk6j6yeU3
kLlVoFmXvvknQRfCLMK7rdAi3Sk0Ik6y5spifN8TGawfsnCfLAiJjWIri+5StsQ6BjkIND8WTD9I
ISJqnH1nZ+9HkigZggY5cliDlonxQRgmeyDJ7jX3vJD2gx6ExrvbmHizgLf4izdrULHJKkTrVDQj
iK4Utw0GiGdPVQpk4HnhghNi4WZrFyTJqvtJGlpbogwn7hTPzrhKD9VcBPaDCnA6d3KzfsbjEFLt
r5X9ZBWpHQip6U6PZty/nD6CTCQaAjxaEHR7H7zMfg4z22ATOnJJ8Q3+b828Slm323qQ6f4jmxQq
XEhMSmBRLdXTSIx+VpD3yqLUAXj7lUl/qZx48JL6/vcRe8Pc28k0w+3nXw2MWJKAOOs6ZuBgp4H3
N6yJ/LjSqA8496lWYgaES0qqq0MwNw7/rCRiVqWl9KLSx/QTwJHzuz5vFCGgComdNGHTQ/17nz5j
Y0Z+rrm9lPrx5gesmrEd+0uYy0+xLEMIEESXuoFxu98TGSi2DVZhwgW5uGwsh7mEFOIHGPgBqcPo
BTeyhLWUcQ7awsvP7U8tjW8/L/X64gpqT8RiGXCyPAOW7CKD0TjfF/WPDvwE2N0OJ/DsTiyXJfCi
S6emDztDyB58e7vm/afuF8sX3xZIDiquNq+1XyNLzj6/+WBndhUHEUM1SxP/8D1S+eFKQtju7/E2
yPbhr/dL5UQplHYNfU82FSvE+4oA23lhi8wR9Zcwd0zM6GcGRpsbmnSnQ+U+HPP59koCylZB1GcK
ejEJoRppuz97i7yjZrX7kI8yZ3oTLhVSYmd/suMQ3XZ2F6VQoEADi/z+vI+3L58GN37iyExl6PDq
vY1jknJtn7Ff0S5M5W+afVIKGctwxzZF4S9fDyxvE/sNui5GM9tGLnnBitnNgwBFP/JHj5aZclpg
neDbPl5GTQ9gVXcVk5uj/yAExvB235DhjBYVUhBJkEUkUHfhxsllzm4MzRqP4hX6qJl2TpI0Sk7z
/sUOAA2x0tra/b+Ho9hJquShm/ZuFiAqMykTs356dwJ6ztigDD1EI2kE9hXITr5y4heXzWHSB7R4
+0Y6NeL/RNa9jDVHy0M3sh94kmpVT8eOIynHa+i2ODMqGYlB8mOmjJLNR82zIGJ87xfvo03ccbJV
CNlE6uwh++WjI7jXxhlL1a1HMZxGvdx3gA+VHyhd6fnCVay4TFHsSVniTIJ9RxE6vJ6XsetOcWSp
T/3HIC19MWTbgve9f0rRov3+RF6myPWJeiYLfDdxvb+Br6/MnGUXeVkaJo1kzSMGLx5A9kWek7II
7mcyuxLHOOXCoRozWKxQIJf898DOG5wjBgcJ4BJS6UzrPKScixiA3CFPIxMg/+mQLEZT1ayUuszb
/zTF0yE7cw9+r1bHZlE1RlFFr5zef/wPSL7u9b9tAOhxxvpOAzt17uEJapHAAhPq3IXTKPfWjXNm
vIR+C/Ti8Jko2g3cxW8rvtwMPYy1eYAeYje/6x+wVEzkFDYh2n3FNJUhORMvo/nRVHTrB+VVZF8d
lLqbUkb2j1myDY/aKd8LtIQfN8BWKSQTMtJweupZ9xUzdBhx2XqZ6vHSJ5UhejlhxqUGeEE/Syc+
zGwLCdakIzCC2iEx4ODa/eyek+qAKDgQC8JclpgxVjwkmynbj1GU79xy34BP3ZVHkfuSJNArZAGv
tkCKpYkzvHSdODnznTMcX6u/06v09zHzv8RCxS9Kn5KonV4sF1tRa9sp1OYz9Qqxa0UGyUrPd6fm
SIeJCed2FqZqFi0zENgmEN5Pf96cjFKKBa9Idi1H1ioNLAMsJjpgIP3XgVnY1OI8bv7WUTDttLJI
pSveSxctCyVIk+eU3NwFzrJUEhpB2xUNlj4E2IZv+POCTG4uTxWkNBdZQ/9DU9Uezlz+ASSkctpx
p3UcjEUSRGglJKPbOs6KkPVPtqyKBp23aLuQkJD3xCkg7lHl+rIDO2KwQWsOL1czlJcVdP4qZiGE
tLTDwTHmBLi7QEz6+Wj9ZHDpBOBLaXWK+gXVTLGKQttAxkuYOUPdexZG25KzLZ6rkLuQtFl3Rzxn
/v4q/O4g82Bavg3OidMx2KFKa8aVD3K3X+TdHXLOyvVYTuAgvyeiA5rQA2rfvqvD+At89OqVnqCU
X57taHCaI2jJl5/kzokExtCRZLzf+x1tEVlUa9Yn0O/2ZDQ32mNxVr6z/fnz98IiRkTD2iKMNT9L
MUVxRoDeY764sF8MedC3flyszE0Xqk6CiGOeyxR6UhjzADNUKECh4kulLXdUnOvplC+oZz/mhZam
1lLRUAzaXWAgdcDPumsMrn/CXv0kXFumT8nLI2LVbdtuA3t2GhMLnCYaQkEKRIi5evN/huPkLxAZ
0Nivy0Df40P3/nNMjJj/uGKo1ILsRCs4vBgwBZl6w4wET1b1HWFoZXV0wa/SghHgkCshqAbsFO0S
KGvM1lgFxwNKv4EJQZRULSyrdiBibqGthbXe5ttBLBB6+wTsHNQEgAtKR5SQ29SV+qPhYI4/GXOk
3Zgkh3T1jKx8x0LfedwjXdmudmyd5WMRGPMDNJ7jRWA+COOHOFL0IUgxhWSpaWxU1w1YWmsMQVK1
lXO0K7O0uN+8vCMp+GqTmkSzlqsXJ3HJlUCbtkIBi8DLiU2F01kNO/nZXcYHtpOysnqIR6Pb5O0m
u8UpO9M/eZo8zi9ia+yzN1Y1ROpXkJEq6vKYg7y++YwIZngj5TlEUrDTAeEsu1FZu/jN4rwx9BCx
JIJWn1n1Jscx5Inxj/STGmoVrI1j+nbbj6d1x/UT0q8CaRzvLX2iDUYIIJ0r0LKhbxXVnwXRHOL0
bz2kn7cWjqELJ3yKKLXOHucC2Y1Rt3r/by1woryrBjo5i4BOXy3aI+veDXrAG6Nw9ujmrBop780N
CZRk8wSEjSCRjgofe8DyJR1xXvyWFjYi86mARU9RnP2USeCrPGVyupbWsi6+FGXfcjHvOOwjfk0b
KvXKWvazg/HPFbAzwDdnwW2vcOXnbUru3+DJImWwXHnhPevdyFCqrAG4st5KmPg6Kekh35Oq4VIT
leK1I0ht7yk+U6MwYmy5XIINgSDDlwXTolSq1vFGqlQWfZ/vsKc+IEWOipb2LULRGEBooYjE6HHJ
X2T6LoYt+7DzeaJamgdMGbE8IMUlOTpnXx9mqdcpSwrQE9iEpBsdxc5J/hursWd56pHcgi4JpxXB
1t3+bQP2Dtof7Df4/yhUI1TrqOZuLM6hkCeh+eP12cMFBezxcaT6xhG4RBuhudLE1Q1k471W3t1+
YY2lhI2n+4kgYSyFr9KVeG8oQcK1+x5lHwl8SgjGeyw7nn8ZxLYE1RXS3t3uA1L7DwM4SZX13Q81
v4hlTwzMkIqFiE5e3bI6Pq/w9i9Npf7TMlp1PpuGnZ1hS9teTKJ8Tw3aKhjLVCag+mbR35vrmsSI
AK+udKPs8CLOXuVR9Ru+t/kgZ8W6g3AeLF5KltpefavC4m/pnqOlALfDZCDAWEsWpQsp6NkligvW
c/XrLK0kco/qL15LcL7Q9kk1keiLozNWiZduDFVCjy91YRfYQ3KtzXAtvinrYz8tNCQwq9uKpqRn
Gu7CbuC+QBI2JU5UTo9JkqcIE3Fs6VqeTbyyL2QqKdpaRXPlwAtRWDGorHcrEdl9+GBLvn0FjnDO
hz6dzavUpi6oIqHGmn/jmx+pinJYLTAZ2iX80zpA6L6h+/6xAGZ6oHbFlEp/9hpfegSVwt77+Zqp
sjpLnqiXVMJao2OFGMpXUuzAAnO1scgJJQoXw6Cd+xwVSuYy8mtAXu/Z1r6KpfQ7WEUZB/vR2qGr
jjO/nIOh0iaDPJ8ux1xIANjTS/8vbSmdYHzdUtIiqATeza4f8aPlaiv2MCC4oPjCmrHBFPrCnUz0
/XpmKGL0YG0TgZqdkAyvKKSbuw398g8VKYVybZ9jH0W/34gd1b3mo9sQl6LaJUl9OIvkzWGiYVnH
70I5bnzPiXBtGxTcmv1WcAGR6pYJUp6sHR9jPgemipw1+moderpnE0w4kCg6X26K3i3QkeQSIiWl
x2BkrAdVXbl49rv/F8F9cvYh+XY9eI4OWKCXHtYaoCWrQHHlpRHhRAw6XrPIt33r0SWX2Zp4yRhs
Es+A8eU1VFP7ELP0exmJbb7MrJPNDMUFqAzJc4l5J3fvlhXj/MktM0NZXRXFf5fu0AXir8HkMgAH
uUfp/7uoKLLMuoDR7b5HSi2mehUpDFqMdPMmoC2pFahzA/JnDRBP2/GpRYN+3BEdIEqV5+wZl+H/
RI+EeVcYBdie4ije1SYGb36BEqOSDKo+DwHTrm+Ukzz5q3JFX94g81dZIqX303k1IO4c9/ccEVC8
oxiXFmrgDpsbThOBVY7893BjDyAA+sh+gu5bDdrH1LvmemoI8t1Oby+ZCVapk+8vm9STmyVyY8NR
omKzuR0gx74MVm9R3Es5yxkiaAifMIl80dg/g0QNqPehjd5xAsV1t2YRVAAwq+uvJGtQcxJKZBAu
zub8waGJBhfgEN2VFUeB0lNO1lhgbGNfl+XK5MVwMHeyEWrhimjSK5mFjl+hBDx7TfAwu7lu3iVE
cnaOHhdghwNbggKoKFqJP1DrZxWz8uhSPhPl19WjRI/JpannmkkQDH2Udd+MhSrZcfAuolSk826Q
TOdEmFw8oSs7KjAXI3mnuLhkAiUaZRRHlDNtG4Wo2qr2vVlX830iqghJK808fXPlVVUqJQozYHgv
9tOcMt1X1PPRKwv6LteLQVpuspzo7N1T7poq9KpRYAWbmmfgecAmmI04DA6lRl08ZG+QwFBqU1Co
u9Tsu24qMrjQNONaCJO562x1u1lFmt/vLxv1TvymmPRTVOeW7K9/FRCvel7eRmcJlbWR3Qvt2rdO
NkFjF3BlYx48dS4VZ1Gx8U1uj+Eqkje2W6JptcvfRLreiSdWOeQsMXPZWQX6f5MuUf49uAu531bw
yhmv17xl6jsWPu5/Ysh9eHH4f+AYsNWvy0KgAOw1A1MAQYWLeQRGfuH/lleKLzT8n88kNMQS0NAC
1VvoVokR5YR90XTt6tzDK8LQ0Diastx7WCtwkZLWgu/dFCEE9Nwp++SUqZO62ouo8Uh6RTRTiNQo
0SoeJRDxuaAQBiCQnjokoHbiI1GBZGLXs2QjvN55I6jI2yh90dPAjx2lSi/x9yd3EZokAfONM3gy
X0KAyDAd7hBLLXYog8zfyy0J2MRKxWE1sHZdW6mR8MqLRSciDMAInNivnap4QYySL0cmaK+4As4a
SFHorrwAbvioGw9Ovll+41/fGelipIYmeAAVEGqc1esmR3va/HLPZvDNAMs5rNDGYXKloHmK22vi
WGnD/IZ5G6Jm69tu/WuQCK+J9bPP8Ub/9FvIB4sFfzvE5d41NPVjcLxjplvkbUdFcY4wzY3R12of
SHHe/mTtW506yRk4SHcGrmPswWLJHsF3Sns1iCgYJzIHzkvLOh3eRrkbfO+nPwhvk/PpLS87t+D7
HRgOQ/pbrL91fxajt+6IKQfz9uUjrIMlaoDVdOcccnyhzLy57RLaEdET3Efxv7bquKfA782WDLA3
npIllIDestKU09XDrVfCiqMJPJR2GDKv9MeFNrToMSaiWmUhw7vrLbQ8tNY/KPw1fCtmAS1fZUrZ
JTDYQuFPyhat9gk1AAIyOi6EIKHGhf6qKnG/uCy5nnH/XuFBTnWELdbhBs16s2aAEXwtEe2woANR
BKZQQm7SKK2R5EBUrhX/YoNBiZkUvmA8jVRWk1FAykh0CKKTlCFVaigt6EunNQkRAEzle9UnXf4k
HOgdXakmQWdCK7qpomUBPrKi140+kr/yboPIPV6Y3xYREtlgQm/5iMIGQaO/s/9T4THPBNzX9+2D
99deLA5nM2ep5iy44EUXYKBxx6lhtGbZZ+2lAmQQz89ikVeL4XU5IIRLxE6DXEqp6+BATwoNd7p0
pr6OCaF/f2ruBv7JuukO6YqygzK+97uVK1TgkZRg2iHQoemCRTSTm/qVKMjHmdJzr+7AfRAznNjh
OwNj7b24n4t3lHHokyTmldiZakwYUBAKhTdp1iX9EIYOsHDqYznPxevlLmPYvw/2C+yaFobcV0sm
gdgFpuTPoMt28iYwyrnoJDJkx7bzsV9WluHLCiI13Ym5Kp5/yQyc/khVW6DN0n7KG+yzfl3/muEi
XR2UE3f8qX/wEpQ8R3XCnRKy7DTEVJJD06wCkG+w3i3BiGv6wntis/wUHvhFpxcLGf2Z6DrEnlLR
rmVKh3ZW65F0LoUm/7pYW6fIhDfJ7DmGnq2yDX+tei7/DeK9FRhCBin/q6BSXWZQ31XPYSCF6mOS
wAJwI2UfiaUukrgQex42/JGIbOfEVBgqjUXryN8J4ih9tpjBdFRIBGn1BPsUAXFsprZ1AzjzXpY8
0CVXtWXTka2ZkfUPvBrYhY63DNjbTL4Y//19ooS8cDwderS0YmAnJgmjcymBx1kZOS3I5a3H3J11
4Ys9En7M8hymZO1t7mEKMqBdfEZyS0H9vybnuIDMsiAHESVBkHvuq7oHUE5PvkMac/uMt+zPkJmS
Vu6DQL9QuF47R5tN+QXi/EmBF1JuNnYswD/PNBw2L0M5AmX4xpnRhy7mOASRn3acLXhXXbhuZan4
g26SwwdW/4PXBQ1syF28n8WWik31LVYQsKQ4PjoOPb1Y8OGqmtJOadJRauumtwKw9l8gvTU3QcsE
/dCZCjX5T8XkYabeHuz62Hm0lPKw+3gkPJ8j8+Lz+6hBmSD2+C5PnAtqgIsLZtUnWoW8igaEFlVr
ckFfY5LI+2jr1M2ieZdxnf0z3TCmFj7U19c+wuTqkD3uAupGMMdl0H6Hr200mrTVxw9bLkkYPRAa
G/TbBLv9qpHFwL1YTRr/wLmnS3ZU4dOhmlkQ8POfg+EchUCqx5DAE38Vo+Cn1pyHk/O8+BulOozX
FUg1/LLUA6e9E0meYyMVtZcyWs2m/CCtjt1yFNMv7P0redCr0leN7ENNDrlhrqpaLrQP8MQ8MVa3
kH5HlUKz1E6ZlFzsv6RvBbP2cAfXrRLEavlssFyNr00BMudIXKmFXFMJ1WjUvijiR6KW5J4yMfrU
QNrxAJ278zadmkKf7WmG6J6+eymD8NB9xVQNCxa6R/X4zu5fxtD5VHb9yGPhgrZx7+RTkoyk5+8z
ZncKHP9Np/XBRDerNdAQIl5TzYB0zBLOnMqp9koucV6gjWbsmWSGc9YPfLQV51fnq7/oFqnRtMe0
fZspw6MyLkZ1Oc4H9HybCIm6rtfKQe5KcNJXS2CF94rH+cGqkRUukG7L2jpkaJMv0lISRzULX4QA
i08icEf6wUYBuDaXrqWoKzQGGSjoM1wJbBdm9k4hOKCEain686n3mOkn7MPVJ71eb51aOHlwaN3M
RhTrxNrQXRzC3wHo7P7sALsGdFOElCGoOHWFqcpEQ0tX65xdp6HMNXsb2+HCkes7JOEU55ZhSciy
U3zm0T7we1vBbXA+OlXwfS32LJiInVRk/odZt2czAvfCXXW5fjLdGfmm1b89c/eTkjOFob163wR/
SVPDro/BgM5QGsvzk7w+qep+eGWlOwweSX8oUL/3UmIVo+EjxkmzqXdDNmKZaiK+Yv/XOc/9jMvr
jLtpT+8kr55DEu+c8tBsiIgpLm2Y9h3h50hwVBsa2bYtpB+R75BfDfwkE1WMCQdHva+sOrPnBXj3
GSXrA6GiK5U9Zzismu1Rv5dOe5CIKa8wPjfJp/gthMECXBpf+7+HgqRIO2Dn/JxIEPzJF6x/iLZU
474x6qCEWi2hVcf2ifYDI2SeMBdY7R+JtdOJwWebvra7Ut/thOe3D6ug9Hmbu0hrDUCRj4bJ30NU
d34SC9rLuvt1GVzpdFBSR81cTOn46aoWXOaCTp0htJ0aM5k2oUAZgRzWHG0vpmkWtzOrtbv8UGde
jqXpVp63AwV1bFV8ENZQd+bWL/jCKlbSssuc476OB1BcuyxEI4T3fUfKKIMvsjTKT8mKxuADnKWR
jJzYPRCfHbM5ZRzJlkx8AVKtBNvG4DnIyYfcY1jEU7pWqtiuWnuQdGVknnK9BxvypkrLT0TN+jL+
AbG9giGHVWGpj+hK9wmS6NEV4F+cyemwAvD7fdlhMrZamQqHOonw/wTEYOGrt59zHvPhi1on6vKg
iGQ+UwKCVxgiLrwHgpEBVEiEOHQbcjK30xQj5O7Nda0q4ec/hfST513w6br+W/zR9tFonvV8OXms
MlU9lXNRoEE6nfIepJVa7dnJRetr5t9Bzb2qIkBsMIBiuFW0P5RuZf9fyZ/WcGdGRIPT/elZSCIu
L1T8FS+BicEB44khdZuecMyYJBeqJ2fTNyyf2fdsk1aKoNTPzHjesFIYtXlh5EFIEOS/1kRoJdwe
CDd+51Lud/e76+cS8w0zGF7yVyZLLttx9nhn6HO6HSQsH8Ez2cWaRDtb4LxgW3FvVICxQYLCe4dr
nYyfqDeQlOUlbcRgsLKEgIEvIQdRES0okyxrq2RFI1tzGgBULbTPLFLPMZ+EJ+GT5mfxAWTo2sgp
k8om1SxftRQzQbR2mpMXCR9QAnL75sLg4TFa/G6rOrzhc/kr9iPXsByJ1R4MgZic2rRYrDR5qzpn
ayhW6SN2G2vbze9tguCeopCq+6acxWP+k7iMF+zQ67cmIlfylL93BfzGdKTtvUUvrbplpxQfqGqC
XEJXk8HYx20C9FkwJHYa73lJwon3VaC5HYhTqd9G5GdwHXA0aAGcrULgSfchuzfLWNyzxrD7IDAH
eJe9vATr3TtWjQnj4UONhZvHKW4MAtYXlQKLA2HNBCUvMfdRP6RCMS3yiPwqUPqAwy5EjtOb4/KQ
HbiGTLU+CMRDTpBMP7IATBqBuFcKpeLuGlwATkyp0iANA0m5F7LKwqYZd5+xLRuOh1IESuQXJnPP
+x98k8bM35JM0/8Mo0HH0EyRvLRDZiTqxnxNJBt5ElxpAp6PWtVdHfzBRxW8ehz+tMDLaM9chXaN
TocsCRJDl8RPKgby7Qov/TgctDQzbueQriE/+1QYLPCbn62hWZNELnx6oJAlJawbeEzpHuT9kjCe
pQqmiXkdEC0aNBueMMXNArpX2LSP/udtwJfhETrxal52dLDng680rrRLrtP7nX5lI2UwSNMQVZZ2
E0AyAqpDmoMKhiCqoJ0Xs/JcW0H5ueI6Dzte+m4gxDIYFEiii6dZiB9n+z30nx9vQ6V9La4cVNRC
5yAKqDKBh2Qzy79RYFvlBQM7+sWFl3KVuntnR1PfeXMcs9x9mydXStYFQxdJjPL/ldOisFJUH5ja
tHlkzd/wXfSdAOyLK5dI0f8DoJR/QPbJNbqA5yXOENwjk63GA41QOI6FEIhkx8JWiwHxBpCEmKPJ
efEbeHvoeu0cMg3UJkbxK1G1hgbZVl5Im7Zlmcn3GiZB3atdVq6ycj6Ub/AV8Pul4em7m2BJWmwI
OXN+kPE2jCjhQqRB1jXldiih23fLM9xS8zDu4dUn0ZtGqZgViyC4CqRtWb6Tu7EiGguVHo+FeaEz
2mmaiR5tobDUzC8KPpb0GWMY3ehLwvHPo5yNF9wv74Xf5EX+7//NqTOOpP7PPfc2HvdF+mExuotf
1HL9awyVMWspQaMbFL/lWOUnCuWmSLVONQVCkv7h5G1vQXvslzr8uY2Jf7dQIK0fE9kHCZlfRoqS
+Dqys9b5qKXXUN/O75Da6Xj/buWviEd5NjHcoD9yLXL/MQGO8ckBaTpjpgQDo0qp2VTOa1vJr7/m
oTE5Ex6elEAUJ0w/vrIVaNAzHLlBzHcxIPwiT2eOghOU2yitKrtE55KDH2eDUyIoO2t9MT1KKuvP
QROVNlNkF3lNjYm0x86Apf77pYy/bhSj6q8yyDc1jdtXBr6XaJYRFL9f1vY9dNxqQQlGzSS8QABm
1HsDra5zOMI1NgtLWXbO71E7hgVLSHS+1veW+uh30EATT1CWZijDefxYP738uuzWIEs0oP5Gx4oC
i1yjupEzeF31d4qqQ8SwZfsQiHcHmHKRTeNcYuGTfwg9M6LorhGtn4/+Km7N2taINF7YyVeTwEty
SEQi/AfAR0JzGoMpupmSkA==
`pragma protect end_protected
