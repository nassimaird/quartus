��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�Ja�g�2�2�*���H7j��
߀��?��3D�@�y�=N�h}�@Dj&>�s��I�3^������̈́_��\���JQt���fLɜ+΁^�߲�ma������Q��0@�y�c'��HW_�P���dJ�ok��'��`���mC�LDr{d��}��z�jg�)����(A��@V������w!)P:-!T���5������� �yB��'���C���OB볰��֟ԗ0�:�ew�h����FS\-�`��\?Z�wt�ǝ���v(���#v�0�km�� {)T������\�w�Vl-��,�`�ScP��?ϡ�d�0ZQ��a�ɓ�j�9��-
�>�������X�D1�M�Mɧ�%�~���}���&���(o#����Uv��?N�H��-㎻,Tp�K�`\^c�VK���a�.>��J��D�+�p��M�f���L*\�$_y� ����J��p���	��BWnq��x�]�a�qe�O�Y�R4��Q��s�H�]��oo����� Fe�lLE�h�UI�����1��I�"^?��f���>tњ6�x�zP�cϊ�}��'i۱��~�I�\yK���QAإ�ˇ�-1������]O
q?u�4C�x ��j�����ve��]&2�_�0%ӏ>�r+�dD��w����G�A��F�/_"�$��ӈ7�h3
�b�FFr��>y�-6�0�r��܊P����L��-�&���?}l���szg��Y'jϽU`�q������2[� Չd4MD���uTo�B���[�#}�����-z�E�<��k �'��
1��0�ۚ�e� E&_��zs�U��������+��C�B��GV�����@nѺ7Z7�+.��E|� ��<JpLD�k�MXm^Rl��� �y��Y�40�D��ď_ݑ4*�����;�~�߮A[��m�t��t ��V�]� RC<���k��wbLR>T�=�O����8 z^!��8���Y0Չ�a��~;[�N� �ܤu�7�/%l�]Ej�70'm!�u���[�F��(.i��S�>)�
7�h�8L�N��$،(�G�]��џ�:����wm���z�%�s�m��Ri��-�&�8%�T�f[���D�=K�gW��߷���~R4�4cb���dKJܤ4��u�!�꼀��B�N�A�[��?�\u��H�0�c��6���Nj�+kA�� x�$6b���H�Mu�w1��nH���5����L8��v7��D���4�x��U���$�B
�lɭ��DU��6�@*z����"+_��ݭ�u`��D��`Cb�N[�Rש�"�>��+5>I��}A��=L��sj8R��0�5t��Zn�����(u~�=�0 㲍�Q��}�qw�U�v��JX ���V��E��Gγ5�C�]3��<���>2G\-l��V�~�Hsw�CH:��փ礥S}�H�%-R'\�� (����S}��;��:�Bn�*sA�bӃ�r^�tDnyK�ٷ�vd:&�Q�+��W>��Vޟ��u�z;�¸8�(��1�hp��b��Q��[8����k?�y�Y�Z��[-'�_-��([������@��x�'��\�)�'���:�-Oè��̩/g�y����"K�݇�j�$���zd�A �)f���4���Ͷ �cq2q��s�&~8���W�KGժ�Ј�s�r��!��62�p�^���h�PV�G����y`�Є8�{���/�e|pB';��-�M���1j����'�����<�l ��i;iʙ(��l��ȗ���3]�I�I:�1X�({\���{<����jh"nr��lx��;	4��/�,)@<?Xꆇ��*�E5oZ�-�P=�?�bST|ցQ���E�Ivnb���ێ�	g��l㊯�l��)�e�y�l���%�����#}���Dn���á��i	~'�IE���}3����\w94�����ɹeV��l@/�y�T9.�F�%�5Y���y6�ֵ�/ڱi��q��Ξ�Q^��J& ���K' 3��ar��D��?�뽲M��b�e�˽�2䵀�
��9���v����V�2����_�B\E=��CD|����?t��>�l�n��4J�S~x�㗹�ҁ���  �g��L��1�PXAԤi�MI�Z9a�BmX�x����v����&1L\Jن�S>�~���M��u��9��E���/"͑�} �72pU��mh��0۟�|��3����'pd�f�`�����=��%sr��u���W�,��$�>�` N8����� %�ʢu�0��t/���q�� ��iZ���lW�s�p7�g���3E�j���������
���/-�ۓ�|�bYG��f���	���VA�����z�7�E�̾fl߳gӺ��٥*��=���p��?OT�f�6�̏��+��)�9iXҙ����ǟR|� q���z�u��I�g1�-�5f�۔ZXSrj�k4V�Rc���������h�>Y��N��J&��OxKu�C
q�ے��}����&|��Kf!c�Wu���jl�s����Մ�A��	�5j¶�R���v��q\~d���/��qg�5�%9��� ��g��-^�iiV�,^t��Hzr=ݮϑ �{�491M6E��%���Ҕ�<�k.���6bA�3�C����t��I���Rn`����j'����T��(�������y��cy�Wh�5&���K~�O��Y�0T���.
�d�����|n~��٣0GF0i֚�:'�w��bx:�L>�|�x�*#n�g�Ev�}fk9���oBH��>wq��D>����\�0�X����lbY�b"���E��J��Ê<�%�߂c�of�^��?k���ՉL4a_�t r���}W�d~�3=�݊��_P��}�l[Bhm�n�*ib��U$��_�����z��d��1�LsC��T�ZѶH��v�Vmpa}D��G��qG�˩������}�e^?B�3g�Ø�hQX��V��_�1�T��@�w`F ?��"gag��.+�kBhz����~�+�����ͯ���*iS��9.W��R�Q��p7�Y�3�T��ןѽ�7�A���V�K��]O|Gr�O���v�zy�����e\��)e/xb'ht�-�y'EZ ���_0�pڞ��Py��Z0L�O��KE+�����b$z��w������Tlpa�0�B*��r��?�T�W�����&���.����d��)W:pMxϱ�C���i��8��7�8Gɓ�*s���i���^�-����r(��k!�X#VjR3P*���% �Ҷ����?7�4l}���.M�ʙLӲ��Ht�h9��JMJ����羮�d����������G���Jy�C����(�6��i<�pg9���6s�9�d�m=�g\xl���jN M�WY�ӵΎ2З�Kا�b+�8�RQ��	����Go�$2	�v���(���CF����J4~&�^�d0y�^�<��G'�:��p�Q��>�G��*�n#�9?�Y��`�����*��; �VP�@�Q|:�1�/.�dy�$��^P��.PZ@`e��0t*
VM��
IZQ�:�g�U��̫�������P��|Z|/�k99�$�s\*#	*�Y�o��R�[��U����5;����]�?ܜ�m�4�v�P��]ZN�\��9#������#���EFۂeeK󗤻��6S�2R�s.�ht{�M ��8\�)��/�ܑ�m�+��,���'�)��Y'��huԉr!�+��2j����#��[�? Rf�i�Y�1�H���'ԝb ֌Z���eqwiD(��cǵ�w��r�d��ݼ��
�(��Q�Ѥ�(����tZt�_��!��y��3\�''��aN�X��P��uY�$ ��k���c�E����㑺-MCU��̿KZNhWUgV��:I��TD)7��8w�$��"�O�tKٿ�\�	l��_��wa�f#N��ѐ��҇=U��M6�������e6�cGã_�Wij�z!�+��6�l��YۥSh_�*�Ӛ����7�������ȍ�.,o�öd�K�NJ}�*>Ts �H�-fd������_b_���T��ZŴ���}��!��p�e�+���[�*e%V�K�}d�v��p9��)�C�N�ݛ�!���mr!6�S��E�(��Ȱ�P1`?�D�@�FU?�A��O$͊B@&��ϝ^,8`�KK�w%���k�$��w����*K��Y��Mw_��r���A�+_��?i���G>��ai�'7}�Q�}��O��C�.vK~�~p{�V�ʹf1HUI�+�a�F�d�1*��F��_O�֠e<��ͣ0v4O�6~��ţ����/��UIwo)��r����ɕ)s?=S�y��yA��B� t�w[���k�[�����J��[�W;�~���h
x_�t��xS�?ibC��A��@9��o�p�5��ݤ��U�)���4�{.=�<�7�����e~�fB(;�&	_���GWvf��aE	>�ᓟ#ZB; ��v�������.���W��ҀuԔ�7h��αW~�5�*�{���e����� ���8a��/�^Cx���'����ɔ/����4��������u�L�O;�>�8���������$ɯ�I��^�7[���Ml�Ey��<}U�|8����=	K�0IE���OU-�H-��8�����o�޲������u����k���P9�'ܜ�� �d'3����`����VtI�A�$��m#�ʗ�=���3ݰ%��0�K
�� �WgJ�D��_�욳��K��#[9��_�t�KN�x�Q
�(�6��4�j�����"��0u�[yšOdڢ��h�㱙D(n�W\�����~���U��խ��J� -B���Q�xa�<�<n�#�G��&����2���/����䰅���h	��G��D3�kбԴZ�¿ժ��h?1:'=�aoox���̧�*j�I�j��S�l�;�҅��?T��^�~*ָT��b���y2�]�b�X��� t�?�4K����XL��xK���i�r�k�>����DH��j��6-4U�m��я.�7� ��YN�n:��G1q�[�َ�;�HV&�8���˲��,~�LE���ګ�1��x�k���>٨�:�1��-LH2��~T�3�/�(�bZ�'�g:d��w%�9�9~����i�Z-�.��0H38e�t}wf�Lື0��,>�"�Î�V�N=8C<�<��i8�1��	Y�i�>R�[A�1�gh�=�b��X�*��>o�VB�����"c�i�_u^vM�:H&E�z�����~��N�B]�\�.���&J�fl�X4q 1)�C�� ���O�[�"\�[��
.�>������d���["��[��Ǒ��>w�c-R��j��c5·�=���n��J��9��I#4&f��%��<���2���!.-j�N�.�%�|m�$���j^�? ~e�uA坥�IITXyz��V�\1gC�����5z�!��]��_wY��u5YkQ n�r@�"l��b*V�����'�~�gg���S$5V@�z�k��/.�x.H���w�K3����Qa���	��]f}����,OA�}F�x�i�{�`g�%��k��Ƴ[����NgX�~�+ �Z�L_���@nȷj���G����66���L5}�����Q/j��938;N��_���q-�"��;w��~z�N�r,��!z���.�qp6��oM�<��p��Ɵ���~y@�M#FȖ�W��LL�&o�Z�8��X�����	�Ps �`V���;2T�����ָ{��06	`�Q��[bY��o��&N��}!4���]R�+3��c
�OlՍ����N3>s�v_8�F���������'�Q��K<9tӜ9�+�v[|%6��ݮ3k۩�D�?_Bp
2�,����{R6��W\�)���ԺЏ��gE�x�I!UU��WuW�+���.Z.��i �_��Ī{.��]CX*�#25e[�����$(^z}��x�9�����quԓ��kk���6�N���K�&ٙ��B�h�`,���&D���@�;=�?^�0�N#����#�]j����*h��q� �����[ˁ� �+���-��q�2�yCgA����[��膬7�7ex{T�c�p�+{��Eb��4�aC#Ԣ]lA�������$\�`�W�	���s7�_.��ݏ	�c�F !whh-b�NV�e���b��ڰ��1W?�o�Jx���mL6Q�3����3إ���3G�$�rW��������C\�Z�������DL�K�N9[U��	����:[��Z5�|ċ�0y�������� ��n8�&�3�����]?��R��A3CPu�D;T��m�D䬨k��Φ�jC�??1��x
��G�}���6�,Ҭ4�AP;�#F�������L��D���9��{�c��=dH�8v��"����hL����8�b�xw���+)