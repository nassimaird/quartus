`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DOUqK6UyjRDtGBPS/yzEyiQyIKbJauxjmJyLyTWykz0816hixz2ZBXq4xorXODm0
vqn4XbmOMcmiyfS/3YG2jTofk7YSv/mYIGhJ8nbMmFAj4lr0r9cpyZEPanzyO4X3
lYbX/Kqj2xK8ZcgkBBQXoIuFaGW7tCxm8PIlWToCNWY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18336)
sqK5d1IJEVfK3Lc7oFEui0eenw2gTv8y1uteg4W9oJVpYD6fzKTWOjBlKqsESmwH
JZksBXFFDuaOHkGG5b5ZWYhoMYyBHH0ZksOs5L1i7er+8N3Sy6g0iIXNO7lbuuRB
Z9YUjdEP+1umnumDFGaAh6Ajg+T6yNEuo9rBD6dZpH/cM4eWdQR9ADCozdjkPmRE
/7VU4wzcKEYI51SFbc9q3nV/jjzsx2AeoDGoJnESzZVbX6Fodkl3iVu5iwceeIWK
Mfbtn71Iih4MrramHwyRm8qanVgfgPBdsAzFfg73wF63PnyLjiAndTYTWdZfxUAc
muVb7Hb9JzhVjTyJOt4MmwxIcEpXnNAMZOMD+bX3YDOwhknJ55xhmO/6lGWTOknT
VZxip3YBGE45pWXbG1SPQRR0HY8QxNBn4io3gDZSDMslpZ08Ptp4ZYUUxeP1+DgR
aVnBXXEawQF/LxAO+XnHpKSWugzr2jlsyoPDAPDu4Ek+aVk7XiaCPiqV9zVfBmnq
anJZocr3vUwCNxe07kPNAOhI7uSm+P7Uk6AxFztRmQ7upYcWT1zE9uxWHxYOtsEU
9A/iLLNTAzPacsBxtyu+xmXYmMkDFZQAFty43nVyaTbyITIDG8eieBC06z0ma5bt
VIJFJpGrSibgGzogb7z+WS7wxf+qc1Bo+P/kTYXFEN8npR5OOvfwhkD3690K6UDh
alQuGJwG2tPCJ8drwoZrpDfZFpfg1PTafKC8exl68c8ZMNNkVDwLJvEI9zEJ/+Pk
79EwnUaSoY9d2RCTwYsFgLwwNJEg3NwTCid6Xpx9HQrFyvI9st7DFjl0yhWn12YH
XW/gYnuNJo82iqFRtqUZ3eywwkTu2Igs36kzmuezjn7+Ocfy6gSk1QR6m3biDjDZ
Vc8RVHZLwmuhelV6VuAE+0fUizlBsiWEibJKx1rUod6WTzBoH8oddO4HM1/P8nhR
UI/RW5RjBlFHn29DGEYbDCXCXkLEGzYnoDjhlTIgbdXgLdI2n3VtRGlQCLIA8fWs
Ki2Pqe3qjk0+RZtNJvmysKP2dpBdFJzzNUbXyh02WwDrfkHSOvSsjOid8e+fm30e
tksZwizfWaVUsQnszH172My8VwkSeIfL9+RddltcyR9O9zc42r9Am3RVfIJkEdbj
I05cc/L6ua71uILFNd5S0kS+tTOFDMDSOln9A3NkB7UuLmoZwNsnn1NmtkSabsxN
C/WhKeIClKsRdp1t5hJGGjFR+o2bUV1l6I4RVhl/fUGLwOwMHN24jcnNGcjMT/JT
B4fBKxHQaoqQrYduPGPZwnOi9U0vZSZqakS/pSBdkP6X3BFBh5f8GdFdR6VszN15
OFWWi0V11LO7sJJAKf6bNSLi/JGZnzYiWqoJSvLPpVWuRXWuFMU39hJvujPl1HL3
Uyv9NUr8wsFW/s4BZjZ3YTly94LfsXBrVI6Kl/EX5tu5pZKzn6qPRIGjcKgCL/MB
JQPCIjCzd9OwDKslrIZ4l69abxs5OzA+fQZB+JoI3TnCIXxHS/yjath0fPDM62MN
0PfBWDu91Lm7UfKwjFfPKwiUOVPLf4Cz83oGMZKQTQdLQYv2X92lDctvbA2Be+jF
um7vlpTuXBFaxk1AIP0QlO4op7p+FEeFZZig4tY4Ox3/6O8tBKkAWmzA1eUfgV87
ovM7w6o3mhKHYV+1xm0NlXG2TKYUAZBmTOpfyZqs4PP/HJPm1qt1JSv2hQHsqXnP
gKFSY15LvZMEV9uQIwCBvlNdMM3kFf5knnoSRajP0W99HgXoZ2f9qN/wsuhGW/lZ
2NRaw3C8O5iPYwFHJ5HIcneJTYcmlMW4aZ1T4TRVl7C9MaGLDVwbTeAqS/RXYiU+
pmSeoHocyVRJ3Wnw9p6pQNe02w+AlZJjnepKbmqaWZ8TikLo0YN+7C84qVVXT4MX
cpH5xBftA+RXVDqtzEL/PlsxxtU40yJ1Mj4bHOIFKQtAanLjCx/Ee3S3FL7kscyp
TT/p9+Hmz5+KtxEhois68P3TTf86v9qzkfDCs2auGE1v5ZL3EAxwCw6Kn0FJhIc9
KMG+koclHJv4VN10HEC3yjFWPPG3bMkfqYx1j3d69yRidQ9lNbNT9GaQ/Kx2r4fb
gA4k1Wwsw/7Up6Fkfnb/+pR2ZSNCleNGrYQiw6vXpY0nBqlLaaxHBIdrCSqTHooo
vjN0HgZAH2ptR5mG4BQmOC52GjjnEqy1MrAwTx9yaSa4wmEHjhhgmTCqQimI8X0T
mAjbtvPN8fbQFXtWXuD+gJYn4wP1dUvHAdxUjn3yto8Kwyr8JALzncgOWK9hMZ9b
WeiSo7RdIIkHBsd2S19TwaBsTQgM1E2F989RAguqV8+hjw8JllfB9N79Vf1VP+EO
kNcWb0V/N6H9liUZwbbhSEskSZOhveeNb5J4MJ4GstgphIfLn6klqlONJnVDAJEG
hi97TYkvgK3w+BXB8sZOdUck/IsKVVOxXmKPQOUpeNkkKFjrr8r21Mkhfnw+kADu
RHGyQFX51KmZpZULV4pBmr5ZYDZ5RALzjTT/HJEiOemFFL1G4rncYfMhOd/vNDg/
00zgwjA5MsoDNFAEl8kEMq2TF+s7bhn8FYMaC+bvqbcazBgPjTelPcSWnJ8X4aRg
A4CqMBNqI3YGhBYr25x0MDbuOdWbtK1c9pxttMomqu4KuDqIKwFq/WyoPMWv651H
8P9Wos4BXvYGvBy9nlCyrjNPx4sCyeMQhKn9180IipUj1RoOWjUymzYxdjvnm6F6
liycmHOQRZRAKqyK335+t0BzJbmIXr3z5IbPrUHrqgKzTqI+t2kOho7bxpMgDWBe
AZxTvtsRh4eaFqaNMj5cWQB5ZsA/WONBHUvdMJAMfFd4IyqUUzOWmi92GY8gYpsQ
znSELxJWzebJUDU7TKWi/rfsPa6FkUCT8zDAIbh3Lw0kuH/rR9ERcIen33Yh2oEc
rb1q3TaR+fwkPsSvR49DTAciCkev66xU7zI/9W3d54LDMl+eYTRAqkXZhgFnB/Ql
YrXT30JZjj3kyoJ2LKrgRhk1n9hWa1HNFWqNsXX6OiiYKoxWMl6FJwNoM1mjZYWv
1PdI/3v/EslcXzyU7RVW/SgFGktemQSua0NroYmvpjNhhjdam+DkMmWrQ/G1BcAA
lx73Awjdjy9plWjCqzuhEENDafWkoav2CkOa9TKpTV75z6U1EDhxJhHwtBuONCb6
JC10j5wFd2Hr7Y/eMB5vN53t2RbLizaLvtTYXGvs+THMFGpxK+p6ZfH5fBjg9DHO
ti6CXNkQsgdu7ciCQ70fhOpP09/KJVG5AjG3ayYQH7EWnAUBMsHXzl0VZp2443q0
LCDjzcEKasLcKBHayUk7aWxDodDg8WHJVDXeHGZRJNXEVYQYxnMgnq/rkZPn8LKU
T4gnJTOBPyyVucuWJLTwHGRY8s3j6ZmnBtS7CmYsXelZAmzmjfZ8iNqZABMD8jD6
642msyAHtJVmjOWUZEVKmJ46NP+38CP4FrZKJWNpvR1ozMVc8r/kOOLslBqTFf99
nhe+1PFdnezW6m6RzwCiv0J4OT73G9vxAOheGhcNm37SUpii4ehmjhGDTbVwZQg1
mWyh4+19CTVxH0LWWb5Qx7qJeGgJ3uEDcDSUxVXPAK4qYG7kmVCX6miyqSkgFhAK
84fkDAKnq/VCXQb31BkBc1sFj410y7vPJLVNFSrcr12ZqsJn0B/mAoYFA5pMQwHE
6Jt1RfX7Y8EYf5WsdM0E5m9fJ1xs46fgyjyU+IPGZ0j/3VKsxvIRA34YTpsPBKzc
m2DRv2VFyN2jMDyeiK7FIjpikNh57LxHvY/Kcu9S2EAhY1BrdyFUMo2zaBcFAzct
K7oXcI3cML/bLcN+beexvMe6IP3QfXoFOD6jWjjfFOdz0psoZ5Rc9QA02/z+4hFm
sOEaSNe3O/PVoksUEEuARcmTp6l2oJK9lPjvFxChiAHFukT0CPdhTVsO+NBpkdzH
WcWd6RNexN8IHux+2W8pu8lZvkbQRbGIYx2k14rpaCQrEy8GrWJN7auVRrNUv5EC
L+PxiKbrBODWiGqNwN5wFjclsumK6aIwNT7ttAU4JZVVDuvLTSyllCDLOv6lusM9
Q9RNowDqHedeAKy/PFMhXk6+qCGwXxbjIQUtfGQBw9oXW4ZF+RYvvk47aYGVuIXN
OAu1iVcvneNfvEVg+rvmzVrs7cQYVyVfmL2n3GnzOZR5KbiURH/Tp+suw6EfbPG3
HEWAQshBBBXwMmmA3AsXs0utA8MX3twqos44Yxba9hYLLH6dZhHqfcOjaiOn0amR
hGWNH8YC59TZNGTH2mCywn0ty6ZKpesfLXPmUQDRVJnsY0BUVtDFPX31t/EGnLnB
rQP2q6XgQlqZoX9+6miltasnP+nNIxwXETFhckl5JQaF/NUZt99SmKoB2hFFIwAD
LGnScY8m3xw6lQUsrCgBtuh/YQqJ7QC00GlwGYcV4aw2NROXBs0FUT3RmzH9/IM4
ukLyqCAIomGMkhjpOSQ0x6Xl7DnI77TsCZdS/byTwg9M4yidn+yjCpAaCA293bcc
u6hYZiGunK+VZaegMX9nA/C2XoMkDEacvH+tr/+ydYUE507hXtiIat1mYqFa85kf
zbHTkULtfixGDS8PPjxq0YN6hTtICSIB+vfU13D1a8XtPyHNMXlO20qCAP9dJ4cm
gzvwbJ/Uq0Ka6cQ0DtbNxiSo1ZnxByiP/a3pFbZn31f+f1q5Nlf2iuCe+tuuph0j
hNnF0oMNTMhYmJktYLt0ZxjnxKW8ZahrHmr+RbodJdXfqlLuqRZSPtEwLNkOOsoI
m+zL5YgFoYsCuPaKTJHHyCI2lB5lOBOVCAjwYI9EccKgm5svgalUtd1dCeSKhv8V
8kplbCeIZqa9uC0gYze7hPk/fz7Zb4UJ8k1uDIpDnjHF/+5wShxCp0FcJU4kbwrs
gi/J9ROS965hz1au03I4rVEgcAJcFO3EfbsH1tkDU2ZT2jhAQHgrFXndi5i4oPFu
S9xvSdDqkOrwFpeJgTlGVYjg58K7pl1d3SP9vzcHTOJJ8dDR16Tbcf6MDRpBnbOL
MI2NLTwrblVBi3lkDe4Wld8tCy6mx/7r5cVWS9QaAXTD3BIv1tfp2D6lkMQUKvdF
r/C47sEfcehJ9LMidOvSWeCeULGWoEDwm0kDbku54wlSiRVbnNacrphe3+BhK+ag
NJk/z000qlgwmfbmiZd5B8M8RMcw8v7oxklPqvgw95WDgQjHeJsRkP+urh9cWvdc
c+7wDOX+2ywrJgt4ldXcVmRRRy6sRS8JDU5edb/lGtMPebhITGFN8WcOLYaLjHas
Tqp0QO0u8vmHT4RnDMITMRHnyugh/48swf5Xk2+n9uBvT2heoNQn2kY4fOyilidG
jHxC7DhVR0B1coTV9QzfrjgSEXU5e0t9FTk4uJWPm+F9Uqfbo9uV09EQCH2B3/gS
f6qfEV0QyZYiy3HiZpla2bgKCGDbFvDVdlwpLPhj4d+R/eR+r3wIBEKZSbM8Cgrb
LHiY+g6K788CcQDUSqxFk3R3xPmR2/1UeXyV2TSykeuwjZ0lOTfEmk5Hzmt+XCpN
vX2C+6Ez0dRK3bhm9/vjxC1gLe1/bC6KNfbu47Kc6U8Rw6WdDnlNEcuS5Sp2fR3X
zys4BWIbBRJ8IhHiR6DWkakhxIUYankeFwMcvCONY5TtcaHSzFEvqGgdxkKwMw5X
GcWMlXkfkp8l72lPRcpSLW4ZNvCngj4dZTjILToAA2ZgJ6c4d55b0/6PfPVdvDSE
wg1MpuXPQp5pjwfrYljFtsP8ScdQuUKQ32H0sdevJY/KqT4V3qv+DdoWmSUVu8JC
6I7YzxtOqOAg4baCxklOo6NmY/PcqPExT2pv9Z2nAO74SiYS17+T0L9epGZtl59I
dJ6mBE8R1Qyp+Gg9l876wKtX41o1xIef62O/vGpBosTm2o0Em8UxyG8XXDrKItHG
mfwu/DtzJnp03rTtlmpnmbDGnsp0e7ssR72SLqfladqO7qdv1Lhl/0OooSRTVVHF
rkAVAlQ9EtktE35UU066Li1PaJfImjjJPIl7MrlULkaJkn94soYAavatvMCjGJvr
iyw2drER2TOso1qd/fU2Ngm4CvEcUFA6oecpyMLaV2DNKiXAzx+TztpJLcFjKQwc
ZqO0hLkH84etB2Aq33g3xfmbwTVCTESbk7gBwB6pv8Lj+eYMt1iCeW8O7S5dCZL2
iU8tfRJBnfrYwkr73vB2rxlVAWotphd/lcpjr2JSeQlNWx/zF5qQ5jY1Ll0hoV2j
d/Jxa7JtC68cEWy9XUSOBu1VI0Q914Yf7nWCywBt642Txgv+VqY/bQzP9AftKusz
goqITQ7cnqqGEj0KOUdkka0OUv9Q9bsPH5cYl2zDKoUuNfrsPe///EcXHPcFJyCb
MGxMwz5JtH4IsFTXHoxIjqyecdrDcP3NsfFg2+rQcX5FrdSQjJu4SNp40JXFJqpz
CN2XJcQGVCgz9aIKP23NxVkASo4Cw3OHtvi4ymcLI07BXwAlYdKS8SShrFbeuLd5
MIoAGhGmaWhclLqoPm2xm8Z8HyAUjmLpTJONGgnKQ+6k+zGZ/S4gHtNM5qZxJ7f6
q+JivPeJeB43GYRPTeGzI5YuYPO/HpplplTF018OsOGvVN6W1Ud2oW+Q70KteyNe
A7k6kh++lVd0nz7FDy0j3U52bE4uziDT8eKIlQFd9pcIRe0wfA0hqnb8jJZdiHUO
b/Q7JF+kvNImaRMcMlZunDBlMDv3WA8de5UJzvayRh8MUnSlzj6ks001OUISXfeV
z6FsbGy0hSiCrqO8QcSulPDNIBuGH3hShK8wPOA2rOXfwvnFSo6YrEZ/wNoRoy/6
MCWS6qyIqQ+MXLWGZU9wrNm7NN9FUjD/gI882vgUuHkN2LzwQYj2NxQ0rtKJd434
XTxVQ4JJcEN0zZ5sGoc+CAzx+nKfG2ZHaBoxyi2lO63unf5rA5vIqlz4clMnBsd+
9TY4OHWgDgn6rG8xtn85dvImPca+5sgW2n5WzGNb/dOCqQQA+1teESsel8ufRXEG
5xlAEIbBprrOaJZGlMHmPEwvcGYSbCpwq6Qy28z8KWIx8JmVUP5qYuG0wn5XprPP
C1+gLJ70Fv7d6SqEAFtPD+LRxIMIYKqQKNqsE+ZNlxfUOBPJwvc3DLCGzsRWsJe6
5lSDlKZk0wyubOFS91jlsFieykOJU0kIFEe/SIZR5VO/RnirMvLwTqqb3ohPZhET
Czgd9WwLAi+sEB5OvHoAQF3nKS8whKSsv32Pj0w8F7FpJtB2nJdo8EBRePYIbiOv
6foheSFML42uplX8FY+xevhDlTP0Bx/OYStgIpLj5uURnRfjkEVeEYbxHHGtPHJQ
dH6PMZc1/t/i1Phil4LP3nHYttsxLyHw7xqtPF36gY1sPrDgyu4Tuf2RwYg2YZpw
fMC6mT7kA//7KiDKNGO0jT54VtUdNsD6Dao9GvKPjARUX7FzOsxNeXrCJ78rE57z
Rcbuc8ua9weeQKKNJql6AMWzJMaZ6VGsB4NNBQUHKjDnFZUjH9h9FFhKVuNTV2ur
xE/jQ7ne6fCaQwSA++vX/YjmfPiZA9mbcIQXNcHxo5OnFykB0Yu43yHTiteglwO7
FMrxyfBb6yVJQtFTDZCWbwIAm1XSFgCgnY5gYe6h/oaqz9+fOIo44W5G3OdoF8wc
EwN1VHoCa3HeszKCXffbjWYM/H+B3++bIiAcQj64BpwgXTIOOsOvbvqkr3iNnUX+
8h8ql9zZXv7zXTkYG4G6hi1hrwUZcIf6VZC6sL2goPwtE9OIfXlm7jCL6hwlwspr
rC2XAiasYmI3ELuCrQnoOnH0H3n+GGE8eSQxoVXJSeqY2h20ENBBIXGRBNCC5Bc9
iquiYKlqgVnmpSCqu+rJtiLEGrd29Sg0XtBfcGHL3qCIPb+WPOHYmX2ABcD8E+XJ
yGQUXwWED0P96oT29wLlEmoBjEc/3Yb+QWqjb8q5+Oin/KK/O9ya/El/qtgi057c
qcMakLHUQa+d4+edWLD+oVcSppS49EPS7ched5iC74ovgALzCVEG2r2INGkOMM0F
6eQrfWi076S8StmilQwypiMaqGZQzL4sqWSLqOmBkblHly7HwhxRKO2IkxLhLlu7
eILPGN2FMGnEDV8fDkDlhLNOO1Z/T0vK28GdbKwEnpyAkRl0QcT9f6IUfrME4WrM
nlqlHW14ilPuSfOdKXGQn23xQIDECD+OThzWksts31B119ksGYYsGEsdweIT3HJ2
kgwenleKTDj2dBwo3C+IzVwKB80VDdfKmDrQKaoV3irPlmh/k3Q+6Sc4slYMoYjt
seKtbNkwhOL7NXlS9UOcX1ALwMMgLIVI/NjaY8Nenmv0Y34bo63B9rUy3soxJvX/
w/9ZPa+0G3ngAKT3BnHtR1OvwZldk8A38oMndlYkwjwW/hVTwe7gPGeo5fAjxym9
6S3Qzi/b7bdhwjxiiwWjZXE4imkVksoufcKUeekRpf0zAeeoe134k13OmG67UkMq
0tvs4G7fIYIcJ/FPhoA5unwFU+0bvLr/fI/OQUhcZfDK8oIck9exoif8oeZ+jyNx
nReZMftfcu6lAJksBAbVTKy1jCAKQ9sdK2ngmd2b5CslAhHEwrbNYsKeBiEQi3GF
FsH0l5UImq8Xpjswg2aVgObKUwHcsRvzeO8gCCZUjFCdgB8Faq3+Yca4Mu1zRo6B
hFvyA1PdeMZoPs3HYggPQG+fhmYY5MOiIwTnYi/qTiyZfAzj+l02+rgEsjJSnFyW
V/ADK7R9HzQkJ9qvJkBxXlUqRpCnfQ9wKDK9JsibBFFUe1RariOxTfrpu+zWMFM8
eB49nU/MG/A3o6T5sekUDQSqp8sYIzzy23xhkgUsakDLg3kA/gFYaxltEddvlQOR
jEDTLjdqkk+mikAjQpgrG5U0tCY8GZz1st5oaqxGL5leq6Hoh64BpTNxosY5eMse
lLpoGBE7zRy8fKLDn8JSIzeQJiiS2sE3Z8wBRs+35ZoJIRIXSoNkyVfc1kyTCQDp
Js/FnECBPgmJO8vbo9dhhwfqfUDrE7tsoG4AwKb4RoOimVdj2uUNGxO43S9GtUBE
AyGi9yZ9+pmN552jEDMlbD1FbCde/BTvh0G4DuQmL7HHLPLHCihlIVZPX7ho4MMe
dDraJtpQ0iNPiBcGAlTtX0UzSIoxJwvlLcYEK0NI5qGZqL8PbOfumwX3ScLns8z0
oi4ag7iDZX8HKF8YyqA78xszRlBHwUYBThGno3bSZih1UuSJIS84A8JGy70Ozgqj
yjaf+kFgGjgcFKcyfB9QiyNpwjKVMhTDQ9EUks/6AJSMQbKv1BgzZOEzLeWHc6LQ
v3rxyKkwj9FB5kbLWQu22H8kJqSONrLrM0WtTyvCFljAd/tM7svFHLE9otrXTQHh
Rf/ZitqJsE4zrwZMjo3Pc30RRwSH4QE5qmPoGixBHHKRu/IAsmuKgdqJszrNPs8s
yRs1KmCz4xzUdC3C5Kc7hLjlHnQf7wZDo+c1JyBgfZrLlRlhqJxI2PJ9L9vJl+2H
ccIdRN7rSfObQsxo+YGN/Ov1HxxYjzjuWvXqHPrhVnDqMq5dnV4FN/tYN8c3Vn/b
E3AMRCLPdhuImX3JQE6psBjzG7171VF3nSYDpWHK47i+chwurP7XVSeZGG0z9Skd
XQp4TGICW14aRwzt3wI3kakJlN0JOz2ABGdgbRqpbItZWXAhdjKt0uJVBILZTrFr
PTQLzi7fKaDwb5Qdz7B2V/XgWsA42YzpQtOZGrktVgzFAvNd8Z6gvq7kckvUI7Te
lRFx93xxfM+xM74d2vfxAFEv4n2YAeOq8r3ZJ9ljk6Ee0sjlEpU7ZpyOBBL1UXeU
VsKG/1edlwOEdAcxFryTozXSZYdLo4LU38Z535yz22ahaOtMNRuBq/e9dom0FvPx
0XO5zpac1SD3sUvr/5g5usPwPKjjGdaRpGIcUf9oTzjkqZod/xtJ+eL+WlpyL3zl
5NvYr0auDlbd2/XKKvJWenMd0HShGyOsR+mVfNkukxzPoB2qJesJYpbhqV9Oxf2j
cPak9n8wUEcL5JPuaDITI94C+O8xU4+S776OkblyEB6/PDLwuPrItThu07o8sVK6
QFMLt0fqaiRnNtNySRs4ierQo8xXsuCEuP/OmjBLu2BQDGoxaR2eBOqJB4CJ9Iiw
biFLsajDT4ksdDmCSaNBaC/v0/mrxqB6E/TFOqFjkf2aHexAZlxhsp9ggX5Vu/o7
okYaXTWIHgBD4u6QSSMHaSPRLc3vJUmILQLuS6U5zo84xGlRVAKpyvhwhCkDUylP
GiytikZCt+w/l8u/jsfOQFzKSENI6kQifvVUWKuNr/qOTuOh2W0AJiS8gstYIKh2
367bREBqyb4AOpGHWo5Fa7OeJFyIi3G+huR+p8PAz9nLwyUtix+pSBUPLmAlhU0i
WMsuVlKiYcSOi/N1lgA3gieeEc53PmPkZPGPdWBVQzkrqVldh8utjiD4f2psx864
j5xIj8W2EUNgkkEXY60RVRgdiwNkIFzYzhSkxQDE9RM/C3qIT2kOy9XVS2FDAJfo
aNBm7hjRrHOPjTGFAMTSuTidRm/ceGVEpuCKuwrtdrkYvgiRchE3GuT8BHdX/dQi
/ArJkU6mIjh/btKPCaLha6zbi4vMJ9cWtKS7syuo2ThnBjNcHZJ2/vbBXQddvtpn
MLHAjmJy+6C3Tb0Ts05eaMa8kaNxoS273BpxC9XIigxfxrU4RSESeXsTPRotG3Yr
D0ozdbB+tfseH9zbhvCjAVzPeXuCHTDC6SLPZk6qmDTMhtt+QXct7EciyTrQbLeb
ugKe1f0dFyaLdvXcL0ukOsWn5bO1t7yUbX3OfJ4YjvN/kivL2tUdzqOLm2iGdzFF
u44iZqomcoA42tc4uefKzrALYAPrP7HNZPogB/3qV/hGl5zA7YUZsyP44vFJ7air
V+tAfCR7Kkp3Ww04i3DA7HPPZiRR8bIaxpJ8xM2bxBmJNYmON+QPHa+S9OhEx1OW
h/EVuG/nyRfMUbE2HJ6vyJLKvhHX+i8QuuIgnHlPh29JVjGbaXVc30t7GdSljBMo
tnILdsgtQnW+/FQNVuCKCz0+gyNLY/KKQjKNBDBPBxDGMiKQ0UnH7u1IsHfssNhR
qKq4a5pvBWljaBOqEq0M/N+rCzikaIThAkUIOf9/59je3PE+74WdwhUsBC2FKCsJ
nZgC6qFN6HQZZxbF5GB2GJoyi2Ij/kjh/AflwpjZxV/0QEpW4E34wOdOjhpGt164
UJsR5B9v4p+lo3nU2dSq4hZuYSwxffKbeYh2Q+ci7oL/IO+qFxAlmU4PcpJ5N3tZ
8nRyQ6kEhw6N0O+4IiJSFpoQwV3RE97DLn1jmkizD6pVOTJHAABbHJlaK9EYYcK1
Jy1dLk5uugAlGDKO+oXWR8inM5t/OcukLvPy3x6/oMAE+Uy2CcAjOdmV9lXW4zTx
IdRcvUzFtTiUJVu+Yn63sj7VlLr5ql7Cz+4W2E2xMDezCh+leQCZEin9Y5UoMAJu
6PjZ4wNJHOlTYN9Ny5gP9+v4CRiYJHXpfwur0ERVijW+XdfJa29lK/a+0IDQcvMp
HsEo4uhPftkZ4x6uM+QBRJ1OTmHj9luWEE2W2VyZxKgcKs+jPvODyZffo/LyAPIz
HnoEMJ3PMxLWaPDUos7oC0az6W7sQZ0SOiSSlfsOAn8/gSCafGFKFSI0q9cIxAZQ
ETujyXseazUAn7E9Tqpkgno2ZG7qLGM/7FQHld0FZMrHNApmsVV2OZ4vgHbp4SsB
8NGs8WEB/ls+Q3AT4XqHX363HbfnvZItm0qX3hc9SHsqYx2cyDjRENlK4QAwFxj0
XSSfwE7nkUS80xtoF3wi0wxDRxVZI+Cq3kVfp+LuzQJDbtnX/zIot0Lfv9bhqNUe
YDFPibu0KctSdH2leLpcgWS7HOAD71hdVA4vfckIasz/cJ9E9jEGAybgw5wXPnrp
sDp0oQkZbPYHsV4yAUkjev0BekwZ5pHy1Hp94RT8lM+8J1aVe2iN4Ru+WWBtqPiu
DRzG5nWtNNIjkRp9o+zizUOmTWu/4bqZsLN7LFHaQLEtVbv5Ewcb947DT6GoIu0U
fQboN4yb2um2JfLPHJvmgYhTLVMWI1qorrWruk/4vYk1M4wUFKtwA6ZIDJoDUHsu
FunK++Hb6R69Of9GYQbeOy8RRcTIiEGqzhV4KWFK0R1LqqU67y+VkoqZ0LAgp0Mx
Wa125NdkM5B2Rz6ueNxZax6k3yDhdxMoUrv8U+r5RJfODRUIkgW/5QddKLR3ne91
g+WK7U0zCSCx0yF1cVe+PZXSwhf0Z6dR9drCfyYZs+VgdNkvK8otV0RmnwOwuQNI
vkllf5geoZNOX6E2isQuEKopGs1V311kvzE43AOG/Pq7DFSFiTPptzC4KOf1nyt9
lsgBonLWKfT2VBqjhlpM5VEgeyog2WZNASizHPWm32yrGh0kNfdX4dQsPj28HzQU
m1fuCVufGnPMACUu15qHa+h/w2+fih65mE6SNUF8FXUKaMqbTqkvIirp7WDxpymp
19ZxuHq9jW9/haEuBCLDVLW2bS0xtNGVfIo9VJttBISHZ8MUYresAjyZt+LY2LC2
N54sU6a2GQNKWjnn3ATLmdnszrasDjAIbQliTTDeklLv1oSYDJSCVPgb0XEXG5pF
ebV7hKKyul1n03Uj+gRKG2Zh2LR3Xlo4/Hdh4/7xwUKP4q4csSU+yAtcPnMJXjVc
aP6hxYuxEID2g1mUumKAIKOrKnaRyKCriR59GWyghwtmkatEy6M3lFm3VwcRa0nW
B3psQZ4k7AsZzTuwhL36x+rCojc1PsItSTCqyAnyRLtUt3jMgtGssvUnqIY9CGiu
0QpQf/oCaLJa2CQp4YAXdPSQrTT3AUkTh7dn7zlux8GOxFBNuJ5j4w5DSP6Me1X9
zjoOCkWSNLJvDIq9QvC/SbhIUIRRossHQf4uehMMNs2EE45dUe93ggWbbDf9zlnt
MCF1WEXkF9EzG3DSiVO16J2Yed9G7zuMmMAjUcbxoyLTPofv5zxylBEDq+C5HLym
fhYfR0HfBZbqlF+Z9Id7yyqmSbfAKut2J49jVL4xcvClFLNqQjFSbp2iZOKMcYBK
sYG/sRBpwSt5ftkyKu96SKN9mrmr2dv4vh7gFyxexvGiaI0F06yJmm+ofBirXRFq
TzjAIKPtf2tAv8IyZZOC0BJcbWi/TOsX8V/w/zt3V/INT6ZXE3EYRbzTgqaGLLiV
8UIrET5BRW6aDez8oMzFFvyKj6X0rYhdb5ApTxbod9LLqS89uF50R1exAzGeeqzN
PdreZ+iTvDoCsupw7BG0n2Ka7AG6mHI9H9Xr8iE5mgXzQwEeHgWMhgVcUFFrHlSn
PlTquQcL0QqJjTsf3PJt49rW0k/sAX/mL2lmKwm09DSmyPNk7HBlKn+VoUP0rlH7
/GHvIOK9W+5E2bJN7wuJiR6Ntf3UEhuXmTn3mvArwnrlbOmqKucoMabu0tgloCGJ
H8hvArPDuDHOIDlVvlKc3RVZnHZ+5fMizZNIFnK2KLwMnvU52eGHuLJKZ4RvazVj
JsDC/fB8DH7L5FRiStoxl1P7DtfCY7r0j2qj2NEb9osUvRRSudKukslVwNX/I2sh
AsjRcwB6ucETzwa2uhbM1EZjAvlrtjr/5xCVBvrQqun8/g3uuohJnwdNBLwipo+D
ygHFDxo17OHnCNBEwQ0H98cyNI0wGNLpe0v2XQpoEtdNkeuLgan9eVtsmB4+2lMj
8sR+EEpcz1f4baGKnKePhLR/zwRZSQd9GZwtM8FL0IGhlNT9pQje0Hm+X9gRJhUY
lBNB7gc6JTzBk+luDLt32XfNreZI2s4B7eVTBecG1TOJqQlbm3SAdFRfRm7mPVZn
hBHZnWMRD+oHeYDLog1jYUHh3qkcfa8EVR4EV3r1gSF8vQSRgknD8PJs27Mk2Kt6
JU0GOwaMi6y55YAaOnlg0KBNUuPn+IP4CGal2xrxb4o+w+30OgjnZNMDpXLb+M+M
kuyWXszt9tG+hvJ/jj4EsJyedBL18F0aGVMRRrtiuWriqQV6XxPvtW53zKirlHfc
i/3PEXzb+WSFd+QVh6D7JaI+jjH9f7ZHy+E8IL6lRKVpBJc63QVtyyL/iDbF2Yn3
II9wFgrZfZv+JSDsUdktI20h6hg2J2arQtCcef2DQsXsKt5dfecAPX2RNqBMbKu9
2JldLrqU0BIbs4EnnlIl2n9+hFxKQvSpJZ0l5J7XAXoI1pSP3qw0gENXgdORToa5
zGB1a2Dhy+MKLXxFzt7WeoZQAzVtD18yRDA1iqSmWGXrbey/ktPOvt0pX6RywtjE
wE6npTFGjD+B+mMLT5yowdn0/O30/hhTDG3Z7T4WTwd6ohBM8b7xbhWyIakffjBq
MwkywVlY9cwlxEwsbnz2rZRt7y7JxBliiO62sNhYv7qeuapLjkO4cjQhm9gwi5bz
hwkLPzECqe3OxCfDXNOmJO4lXcFqTOk0oWB9+kDYDZ8oa2gecNZ6LRwV9ELtsXNC
bteU/AWFQYWqHITU/nf4ondIp3W+zkOvN2WTol676Rp8Dx6nJ39eCCShnNQm9NCd
6VLxpZu5L++/bKX/+bKrLKJvBWRMgQRSpKeRgql4KZIKe/B2PTVZkTQ5GA62fO56
fbdMRsoCa7XXoPfitPN7r2nSNHut1IBSuRED9ivFsYP+MydnFwDfDNVyxjzTwDVM
CiHy8S7lSHRWEcwUtHtNyBCaLGzBjN/DmSA3J65wNcDTSYIhXlj/hdiA6ZcbFBuK
j4fuo5Yyw3w8FCf2tG3loVAbYDetR52/a9NM1I0Y6dsqo8EFMhE2SzkMhFE/8MNm
3Plu9CMTSUukHtk3ubnNxRYMKwTJ8ppZ6f4MTEVl0PX+Lyzzaj21ToG77kThqwTf
llsc//6CMFXf7i/CIPT61GxSOH86xP5J3XCREUs13/BOQPt2dM/KnpBm7aNEVKf8
pBywUdrOgwzY69FOBGvPqs6RXDE92NYAq7BAfg/1bs9T56PeHhiXnY9UZ1z8oBNx
qLPhJ2B/vN+3FIR6mfm6eqGph5y4xdetNd5Q7pk2xtNqdkgaf5ppNwG5RtTabMxW
DdtyIb2PCMBS9mFJVyIsYM2zD/QGX2XDKwmPGoccbxJWqugwICabgmQsojYmEoks
woB81Sv9g0lv+m/5vh6cVL/E+QLkqgOLv7VtOmjy07EnfhlSCS1Zd1e0dke7jBNT
CXpjEoCYerCN8/bksu28g/Pt8zrIsVzKIOIx21UtUfoL4ycNsRlpoK/Rpz5rmQ7Y
ZXZI7h/GQdvVIEkm6y7XoSx3X6HT1JJevC8y2R+JEgCU6p0tkUKpb9vAQ6C6QXZb
SzVER7qi5xpMMRW1rVSzZzx015qx/NqX5cp1Cnu80CqzA8hQQkOU5JD9TGWgx1/c
wwlonA2ME/ZPZReoyoEGN3wqGnxiQtNBvceFG4bjxs92yzMCNJkRvpfO69moYFkR
dv/HqpoXrquFY4vmfXam4VmfNPBvdsuRYNXdNGfjpUPQO555vSpCgIQvWvQwxAiq
bCfn2/6JrWFxjO1udpfu6ubA+HHD/FGS7PR+hSBuCe1/2/0Hy014Vsdjjh/XM1hM
GTb60QoPGBSdEgnf6F+Vsf4f7FN2pRASz1a7gBsPwcVpFRTf7gZQ/+Y6WcibMDfJ
prqU1m7GX7g6EQJy4VVlTJZxwJP0qOSV8iQIJK53uQxfo2Ufa5/uMAZLAaFJ9BxJ
yIWvtijq361rfx/x6Z3NE3CkDSVwG4lY+BraezMz6Q8K4BtNC0Z0PhOJP8cTVLu5
1Ai3Zw8C/zDdGutnx6CfbTk7zHpon+3BQykDCV8n7HAS8PmS/3QKUch+VkzrFizd
imQzfQV6o2LhIv+W4P6n0Fnjd4kFXnl8xaGNENskOs9noQITjHZA+Wh6ulIIeg0n
9mo42v2xOjdA/Ei8NggubKhWfNU4NVfhMti2x1uNwuxf51mFplPolULgxk49JOaS
qV5r01cUOtjVeebCxZz3++jzVrqgwklX7uNZSNdQClEVMiLf0zeYFlPnkMpAuhHQ
yU2hbeXQhx5vNRHIRGRlSJfNQ7kisu1Q2yTDws6KpfIzvy+HjlpQs/0p0Nva7KUF
StDWNkW6kn/TPqUw9Z5enK7S88jzkxN2Ny7isSWTC12VXj//ewPx64Gx1/tgIA5R
AwcmKDSF11mqNd579ktJ46q5uB252ehXO76lN3dtN5qcKVwyR3nRX9TXytPI97XY
EklWZB4Vlc8gMleM27Tims2f8BiawQuIhQDrT2FAUP0iHQWBBCYlKTpd+1j9Eeyq
SCHSOkyVvKlkM4cGM5ocL/t11PRdGlxY0IFG0oO4XHBDAlEsxlmec7MeCMTyA2WW
ZINApmaa2YlY3ok+3yrrS1/HD3uMesSlh052qNK5cY2atz/9IPjvrrr0z1wYq8fM
UADflQpFvur1g/c8laHLd0T0n5K6JiBPR8gsCKZBK7j5YRreyaK3hZHezxiXjCq5
Le7PdFaBIOQESjSgl+JSsG1iDN5UchjpB/wfHA/WbYuAGSCxlJH69WYBr730c5BK
YCv6DW91uv2pUp5SF2MphAwhA6fl/6IAL8OeIvooqzzHh1L6H5poIspBZOWN6wA8
m6gtMpjd3h6URP8NGxowd7RKxJSNe14x8mMn3ySNb5jIVP2dfKiUZY8yYuBo//Rr
dZrox5zqXG37FiNT4GPSKwvvq1tUv9X/qrdt0aDJ7QXtEZoqxHKJta29gHAOAi+a
/EulOgKOsVRpCai/o6rD9yLC+CmeT9EveXi8Bxs3yVLiMJJ6ONEp383kmSmnWB4U
JXJu3tvPOmKHzyBAnQEkiK6Bms8nVv4R6YavoPKnFyLYYzGIvn8KSpEGF2kQTvVH
mppB8O/n+qSUquVKZydcZQrFc0PkfPdhx9RlqFDopbWgr2sh6BmKECkHC4g72LXW
L5WPc/SyZRU6Sz9TmIJixCTwel9eTW5yiTghNNfmNij04POVd/CcIt54rqoOZYlM
38VCsYFPZcfC0goC2am5LLWM75g+BC8Mt3Z3lSta2i6JtGHReKj2xJLtd7QYVTUZ
e3MyLFILpqHphZ14lw3tXmHwsyCy8h/sEZr2ZM7LfVybUvfevDIGflUaD6/LNH0D
IARKQjuLF9lgvPqKYVMFZWaY5ipiblwzGjE7GwFX2Dm5nOJhE+912BFHMk8y4vu5
gBkClCPo2L+KwQxdLk4nGpGM+kMqeuT5mmQVMJDvO8oBgU1KtgYZpZ2/kCl2HH2m
jrWhODf1kzBslCAP4G7+/5rs2OLl13axWH1UoS/RnbuaN7rpdhunfwHEU/UoDOdp
PxdjxIk/Q3gqpEuvB6m/qNrZyFprs/p/aoMmFmP5YRSg0gHKjRzM4LvWOUs4/ZYx
VogRAcG6egyM3X3BqkKK/VmEUdyNsnLn2PUjnTIGQtOLgviwcDqhH4gF1TSyG5rG
PvCCWkMk875VKRhcvvinKGtCQwg63rWdaCZrmY9Y7JbiGjUPGX5famVto40aJLjK
gwAq2PUbuvlwfe/g7kBT0alkzH4XHW/0oX6drpioHYuWg6brwXw0IRrofjXH2D1r
tLjvIu/M6CMteuuQPNN7QlRVx3PEBwf3FtvEyRHNwXvzKq9VvXB/yKLUKkDeokge
/8QEzcYr6XCDzdj/Xjy2/nnj0pdrwAoterGOdxrcIMc6GgCn/jVtTRNTKB3Q5pOV
bzF95ukrCuyg6yJXFLHeZI46prkVS2d/kXPHHMwNuX/7JZWSDK3RMBemy/2Jc9B3
5dIuYs/eGEnbEF2EGEDIXDpCd3x3IR70wlknUzGZH+5I5QRrSVtsTcDcnOfOs/y4
U1simWjkZD+CYNV1cdNmQB7J+gx0U6E0KiiY3YrO95whMzp78/Nv63zJnNSZ0onz
UQqFBMwolyF1QBaXrnVoYgdTbKIUopxEzG+HHa6QYASH7cYdXuITUckQFB4tliJX
pbuapFWodCDko2E2VUfZ1AAJRCyPWDkcSlEdaxkk7AxLgHQKZnGrAzZt25LsbVHA
syR2alUR4KWwVraFOZiNa0iSQ184mb+EUyLUFX4uLubnQ6LpMZYhszjvqJeDVXAz
G44UVc6gBFQCSWoeshpVvfRdyQp7AiFtB1tkKo9z8X+5ubGiVTr7YE3eKovfmPBE
keqHkQ0Llxf2XS0EDTHvAdcEICmu/eEq1gAOaQ/xMvkn1nvD76tBg887ALQNP10y
bPRwXUVUX+UIn/9h8KQMzcEChXX064lIxCD0rtl7VFFH2WqnnhhzSnOtuzYXCrN1
mRs7C/yg98QpPo1JuuqDZPsBLuQet3VFm+je/Z9ji4bcgVytkHSZZXUBUJAs+D+r
cl1mVRTOai2Datfwy5JWVppa+msktkY1oBlDSOmNErNwmsoA10rWSMWC7Q2U4P+T
O1HLvKt6cnSqwQx2rFSnF/tyUMd/CWzhDRNf+F3kUnn9jLt25YwIPNtkTi3YqoAs
ymDbyUQ7vD+XElIGCXAU95WoTEAk2pimUV6RezKRA/m71MYKRiYIjWBrU8xtFc3d
1eAN4e+emsQNj5JXTDB1EgrgtkhxFlZMa1HXl0IpGPhurgCrU6F1jCbEY7CfI8lY
jsIu284Zd80MmPoa/DfuskRXxSSWUkD2ZyaerO7jQK5GG+JP1GYmd0Sj8A1njpq6
/Kp0KTFpNsabKRAKVKqDm8GghvdylDDE7QWehp6gCf+yCIyH2iaF5remrws4AVcg
sI1teGFzrriRh58Xpcv2I1dJj21rWiDX9p5KOBZlm0QkOaONScP+XZ+SCHNSV6Vx
2SPtl1ZQ9pPqyblql23MsdqcOBoyXWvXojgVSOYCd5svfx8gI2Ii2sjRkEB4FDgI
NRiTPPBYr8bVUsrkWt4NE0gHXAn7mudWFxo5W3KYKTxZ547xSmrpRfYd1cgeXHF2
KY/PAIudPK7sw9yiC6gCFVmLQIUQbJXcTL6yrzQ6aIptwJtqZQE1SPp5X0WHj8GG
9c6iwcDIXAfdP6ITe3n/gH+gQCEi3y3By56TLbjyBX1bGLeR48cZEwVUIpZcQptd
Wk0WAfxcL84pInVk+FqN5vvKLY7bc7J1ZvsTF2InGx77h8pfhAwOuydw+ZYPPo00
ddcm4OetgDIq2v8b5ncGIeatbCjcz2/WEGQMQSQIjOWOjm/iq+Q9dcTNuTk9gKD8
7J0NF8Lp/UTlSDAgMRudYov4TrnGx4km9GQ7q53LZfa7zf6+obtIeAqUuSHNlfMA
ilYf0lIGe8uQVQyl7HUE0qUyPQ1A+Dgjj9c5Ax3JWvKW+YKJBj7CpVXWPb++pgwj
1ODOZXG3wpk+BA0iUCbiVOCQ19IBFhoqOp5Phk5zSOpdZd/AR2rTWYSFDKqCl85s
jWSoiBIpiOD/3sy9MvI+l+nLTumtoqgwcHNyijY4IQEPLt5nwYsQRr6vRGbuBb2X
VTAyGeuQBMHRsbUcs8sTnzGEW9fj0eCPhif7K4thfSll9zn359LLclZ7aS319ARJ
GIr+hfWNtia1wKwEe/FhUNy6AoiBk9wXdaIMl/D0IPqNKfNFKwuo8oGf7jBK+1Ih
W5q87ILp/qfz+VRFjk+dJ1ezxfA2x5B145Cg+IjnfCli4Vr6pbTVZ4dZGz/hJ5wY
G9Qjta2tqlpjyTN99sMzKR5GALIpbVjI7j2ztKftdAlEvpZfdzS1NWBYi6CCyrPu
7ge1Z8+bjsEnz9fVrDIKL40f0KRWq4pscNTfJxj6xuU8i47LX0BxeSnI8yo/I2bD
CgzAfYe7JpoM6Bf+3cGC0cA63DAPoxG5aakRAkNbBbWtPEO2DJ/SqpQVJaeASMVl
Mz3dIS4xjAcxIaOHPkbkpyXUpN7s+fqCtpkdrX5YPFoSyJOSn4zONiccEV2+ueHc
7lcS9D0FXj4TLa8g5QXLeXAKQoroa0LNBXTz0xr5rZ8yu9pSjISzvi7sxV03z+SR
gyziafaBYJXdHpRrHl8+e/A5jO335CEnO6/gI40z6ZqT/AJg5K7+jEkqYD9ynUmY
q3iiPH0T8VSitZJnSqLH4/GIRu66cclZwgJV6Z6tPCZl24JhSUzRiUJhurMWpXZC
dZixy+HLxiXNsG+ESnFlx/Cde2hi9vkEFNsUKa90qZ4P8c+qVoMoTQx/cARhxn8R
SL1Z54XrVLr7PuQVUXZbomm81pKCzNuBOfSI0fw1AFPgUtnNeZjgHlUCA/iXNCnH
cQaPXK1xKL1f8v03CGVyQxjXpk+OEvNzY3SxmAhoKcDVvQIukygD24d5kfkP+Ux2
CAP+mZJdeALaUBIbcv7c7uFKLj74PmAERx3PBV/BwElqbeASnwvHBum7nhEwkHH2
h4CbziIdgpVoavabrN7Qr6kNu3OBVPSHHphYGBTY/T1e5A9kM+NyEbprLhFb5FnM
n7uBX/ihXfOiemgBt6MN3bjBKUk57Cas1CbzNp++TMncDg1ivkxde0NVr2YRNjUC
VjrD541P9c8haBsTOJFdkSWcKMJUr6GL5/MGZZinuvHhXEy7c0GFgxFYQrWE8hXa
dUv2Yak9cmNh6VtTD8EBxFhOtOTZC64KvqPOsdqpQXoeAws+h73nvcgyZja/Mgl/
yIRFmSo6Qzrh1HfxOSDGBAqRnIPMweknO6XXb/G+5/CevFfT2bFJ7ugXbuEJCr0x
KYmwoLN3qQRkJ9uEhe/AjvbIJSaMsjca22zbkpNNMuTLy5Ed4mQ/1VqN1wWUHuTH
sm+jSSNGo0UMaEMX2CZfMOKVqsfev1boO9GyBQ0YtgU37edL8J6/w+fezK8Q1pU+
/yb6nKJ4Um7i81Dh6PDCsvqvy6lLD46pmmZgi9tWSByTitbzECpNW47FRSCIrbpk
Caj2JQuK41XaInnLQ+8pqMTEA3Mues5HuZP3WKwJb7JagUvddZBxh2Q6LNH+Qm4Z
2pYOF8wdOX+xyU/lZgUBajkMdNY9Id9oEwLzaDY22RMDA957wWvoSBan4yDYdUXX
vYODbKB+mHwOICt28OTIgPWn7u453N9O54I+fcXMA+s+wkmwY10jjps29H/aBRWr
IRyFODN7ZbJdgeQKqkqqtzV3DLsXj0Ezl6mQqGoGLq0a7eO0rAtIjFdb4gKjiwsY
S9/Qdg+wiBkK3Vg7zt4n+uwa6LbfYRLTDLo2MFRUK1SXuCWfC0ndAtwILYWOz/sm
ZpCcq6vLly8k4vtTISghC2qlz+n/egP5l36PqKReXzsfAerO2Lp1BzdES7AqxWn7
qd6CvTQhHGWcPUDZgP1sYNBRZ6792ArH6+9lC+0qmrEhCmiaJK9SVQk+ZTP47RGN
IJkhI8tu7KM7vWM63vrhaX5/owZq1tvldtRz7pnI33b0YNXgy81Y+GsMbrC89aHC
1jPeb2OneB3FSzokJYSDfwJqBJ7uy+w+X4j7I+z62XJ90vfneUkQidNe/bMjGYMY
ZyZYoXf3oZEbjhmddHz4y93tGPLv4o8ZupwFlAQlSqrTWwuWSB5TJhY3UlAPs4JE
44Jso+XqRzAnr1qtYmj1t7geTPKz/6VMcPskLaCk9r6knyzgh+w7Stx9GLSXClQd
FWca1LsKfZ+OS4BuL6155UFQLxWts6JIjKPNqzY0xnWLTbLbAwhmFXtVx/1tSRad
yYrW0bXa3ZQFLUeMjAmcbKjJwkN35J7RKvI+m8szvMUO66Q0e/qvwAyVfcb25fBY
9WhdBb+w882BFgCB0Dq0qA3mMH8cK0Ajgs17EYXXlKwaEabq5GQrVVAGgHkl4GHt
oP2an1da2HIsACKRWSDSHZW92/V2YIXtjLTO+pVX4oxGH7xNajoNHKomIaREGMbR
K7MDe7XoeLi86YF8Ft39PRkp4xbc3Tk3cDn8407e13TygIu6QACsOshLdtCx8Lyd
732S+QvLseM5iJ7irn8Kh3vdDF9ZhVdPIaLFRC1++C4q7swcZ1Jd6SL65yT+vUyb
3kLpIJPR23qpZH7R+HGT40/Q399uQ+1r+Q6vLG7N3OFg5aTGfUvyXSDAQk8x6j5Q
xa+UcAkrf83njqBMuic4u78N2NOzo1+V06sbpxMQsQqw6/VhtMCPfpOFuhDiS5OX
YvwuHIfyLeDK+i5FqtcNos68WryoXMlsB098JBTS/HtVKzMW1Uh0uNZvGhhac4bP
PEgTiIXOGsmLQK4+94Mzp+fiGCX8VsqsxqaPYkB9b2tWKZQ0VlsPXJmJkprkSWvZ
D1rw0c2A7DQ1JzNxYKlH5vWqIo8GkhmJ3a6gjeRGAE4TOuHcqz5fgNiqn2l2fUMP
zrlQjxP95pz62A87SgAIcb08Zv6EP8QcCL3lcjzO39Asb7lyDn1rRsJjPwP1fE9K
qtL8r8RFg6Hl8fMH8SWOYYjAeKN+9I+Ic04+U+nHdZX2KnIgDjyljA3v58ezf/Bh
1vdxNlZWegDPg7EncVkJoEvhApKeXlP7TQWZs6ek7+f6ucmesqMt+F/N8O76A4fO
k//K0RlbkRJDhyLvc3yYDiL4HQjIn8snaucm94tvGYuzrxYvtT1Vm2SEyFS5TCEv
9FHawtxh1FuQsADpzPLfRl6Ff6p15zoGM80yLLmuMRkfn06rMmjpoX4eRWr/OzQY
R/nXzxnu42maxqqmr4kZaO8aXPTFj+KyCWmaBcKEDIPzMV4dOMUlqio7NpFC67Dh
f7zzG0wfXvRApfb8iVsfAwz/f/jpKMs/95XA7+SCjuAk/pMnVUZIB0wY2ZEDFh8b
2SBdCbwm+6StSscyGv74mMTxFMC2e2esnNo1al74jzREHycJ4+sxyNF4olXE5onS
XZjQo7wtq5mqQ3GC+jYUC+g/tCDSMXnGb8SMkOD/UVkzHSEQ5UrvDdKD3cdC66fB
9RITV4E4GhcuKWQ/8mnKd4AvHknpDtoq1PM1yLAnLIEmQGxKIkG54wdRjtd8Z7MB
wjN9Pkfv3DrA2u7UIWdYucG8yGu73Jlp4j6Y7MDdRIyi9PuH2oa7RQVoE+7lKCAP
BVBH4gpBBFpvyAWneFXcsj2CUFprNJ/gGF3PgBov+H+v3SIastYvJk35F5z46QR5
MVwpx2NB9K1EVXTUO3zNNoqMN5Vd8g25TTFMK+IFymNXyWtvKiZutMWVwRGhSRP4
+xDqMdPy9z5A2yl94BKibNqVjyJyM5f+1XdNToysKxBCUI0vkxJ+2eUOGZXeqqTf
Cmd3p9EfUmNhFhjLC7vU8PEflPrIg5cMo2me54Fa3LByTdfRcGIj9Yf436AfD/3F
552D0AMJdNqM5Ol8aIWYVV2hwu21AEmV7peLtgD3Frduln6dotIN7ZUh8383TZmS
U3/0F+VS8zy1BODCAgf7H6OGc/by5b+25+2tWo8rXUxS/G6YYPgDiHesoGmavw6c
5pfN1iv4t8YWnyITw3yhbOL/4qjeoxQxbTMueesdWSCmnl3DiWFOpuvMKB2ZDK6/
GR02x5DyL8hYaNA45/Yq13Fc6cy3EoDF8S/+veKNisxfP78P7xO89Syno2LyxLMp
1E0xJDYfsFjLumoWmL+EuP3PSHyGlvImrsQP4HjcxaOYP9lx8l8qORk44M0oVp67
dS6O4riZHJ6hS9KAHJ/lRl6guz3tvKcq6mkhHrntCI3XVaCRQ/mjKMb+3FcHx8Ns
hewN4gcr3lHusUpEujly3pk3eQvc4sP1+c+hFdE3NkBpI7KZkA+PVK+phu4hVh23
oafKLWsWLVrjxKlj9f5kI9GYwGEOjhqyCvvl8OabpJ9fWq0mqaSBCnskIk3CgLtN
N39NQ2MEMlGlyzVDm5/WZXrdxRFI11rFFvkuDLwXueIPjIPmeZpLHlJvwS8kPTRJ
XsH80MfjPyGV6xgbeGYbovxZxRTE6EKW2rxx2ziVqpyQQqx3T4BdqIqwcLk687wP
ZsG+4Qp6UwdkltFIEeKTDSP7XoJZf6ZOgCCozbBsDa3Qysx2oQOxuOaibow2GoKP
AyAfEm+rmMsdBAAy9ftW0Negp2K8lwa2CQJ/wgt1U2BcL7FHR3/w9uov23hl+iON
blY1N/ge6shkQwItlrgMmbRAbVjsGcfRjSPEogPV9vInD7UH4kg6X9p1WlTH5Icl
L0s2SuQ3MqwGie/AS8lfBS7hNeCmk2nVlQQXRQZBSn01N/ciICtI5idqQdiAZKHw
mpPjHfSpyK/G5Ny9ZBoqJIuksiPBPeI6pg15cKqs//4pwm/s8It2MwJSt9aLPgs0
7cIRnNt0ei1NyEIGIzacWSxhJcBc6Okl4HyD7oxWxX4c6gi6QLVw7Cb/C8VfGye7
3xPJ0snBVs8VSI+CyJgJKq3uPAHdJHPf9+FNfC7CsycX9i+exQAcKUBB8AUCbNNT
l/r8uIrJcCtYgB2TNXL+9BE2DUGq8/w/LDU3VtGLjUZGrKL2p+1oegIOXInjeDzG
faqTz06N2ikHQB6/iFmyIJmEpqlU+mBr5MuY1vf3huaQEst54DZ4n0lyE0VW2T6P
`pragma protect end_protected
