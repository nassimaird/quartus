��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�U���_I
y��������k%̜S���9('�X�@�'�X��m+��G������g��d�:]�<'� F��-!�k(�M�u�=X͝c���/���A�l�8��'?nZ�]�,�u�������k��ᚘYڏ㑠ڲ]��L���s��F�N��o3KK�+^_o;�_3B���'���f��jI��j��ŪD����8��3֓��p�O�P�hD�����ץtT��Wp��ZӰ]1�b��#�A�H��,�n�ʫ�I|�_T#{i;��5�$mX��b�"�(���<�B��p�J�O"R���Cr�7몈K����r��K��ΐ*W�`� �s���2q���k1wA#���k�b>����8��0~XӋ�ub����?�\;VQ��!�o�U��u_3��7��"�o r��-�ڙ �j��}��q�4(��jbu�h�b)h:������d!$_���E��FH� �%��?�V��o��[M#ߕ�>*8N�5DIba��lm[����������)w�3����#Gk��y��~�*�s3��£�9�eC��>��U���.S���u�_��D��1#�����\'��v���O!��M�,$�* dM��Me쎶��ʧ<��p�9:�`��[5�^�`�e#5{���% [��Dnî�]���3^&�'���l�z�t3�B�Y�ׅ����r��Rc���O;#��#B�j�R�&@3|N'h���Jޒ�1��j���%�
�on�{�����}��.|"�R���BSaN�!鎝�Te����o���ݬDNn����Fy����T�my�jH��z�,��(:��������`=�?0�%���I�;/��÷�ₚ?��U8�ay+�SQ1u&���� 'a
�B�J�Y�����M�DX�Z��jnހ�CI�gN����ȵt�kd��zΌQO�荳I��(G������7�dQ\�S��TbҶ��%��t��0��@�
'����v�8��-�`�|���V�����M�F��f�P�~��I��d~#x��z����.���L��?��D�7.N��n���U��gI��r0�T�[v�`r��B9g"#���JB̃= S�Q�<έ.�g8�n�f����a#Ӫ�Q�Q��� ��_#54\^� i��e��̷t�N�K'�[+%m��M�ee��MX
K�D�lMa���O�Oc�F�Q䥡"��%\�P3��i�����ByW%)C|�nőE����+��w���<�ŃmE)�}�V��� ��x��0$h������j�� �1���y�'�yԠ��iկ�TO/v���4���M峛t5�ЬÞ���ϖ���Y�j�P���G'�S��ǅ�px&�¾�����֭ۮx㰰O����j;�W��D�xuf�S�\��M�������w������2�PV�Z�?Z9�B��X{�OQ-��p����bX
?�A��t�gg	����	j�3�
��<���&$ZC�}�,�w8��-N�V�hWhU�d�#R�P�b���ނ��o�Z�C {,�_ڳD.��5]|�Ai|���C�t��ad֤�'D�#ZN5%�"���ӵ'E`@vg#�K3b��,_X8���C>��+��ä���5��E��Al���a��=�ʽ���Co��v�[ ��z'A)y٩��y"��۽p��LC���=�e��ڂky?�ŦS��*�H��yW\���y^C�y�{�S�ؗۤ,��Lf`�+�R�.��i0jF�����Xo��A���B���hI��O��C�`��>�_Q�wT,Q�\$MWd�u'��O��OŅk�a������r*U�%�s���ơ���-鼺������%�!�?���J<{4�u�&���_��J���j�Q�e�BH��~�e^P��h�T��q>���gD<�F�U(Kb�Ė�c��o�&���:��\���HB�P��"��q�Mpr��ۚ�k%i����'��,�h���.�Y�9����~c�+'����u�yHo}CW�L��Z�6������Vc.���y��+b2���ם����%�#��Љ��Z��=��l<m��|R�����aפn���WYB�����އExv��~�ټű6 �~���Et�s.i��As,�������w�ڠ�Œ�+�X/�H4s
yC��L�w:����>�{R�=��6�|��P8��wD�}�m��A��--?���"���\Lu��`YsȞ����&|Y�b�ֹ�/y�3��~��)<[Y<g�\�s˖�k%<M�l����@�5�p&�a�Q�Y�37@�LhTќ��T�i󖴬8�_xu���O}5��p~���twd6�EBڽ��Ֆ�mhܚ� ���o���ʖ�m��E��~U� *(Z��Vf�����S:x�oN|�H�U��w�"����tň��
?��B��<T�\Ϡ "���©���3�˽�b�v�����}ݕ�˼���p��ɖ�Ŋ7d�E��-�~մz�����\we歰>��8Z���]Ω�Z�=K�̣�LT�\��U��[߫(�5&Lؑm(��G�zh�%��
�]�w�uӢ���[O���[C(�vt?�矓�"aC�w����;�sNG��±��ϓ`��<��`��[��hEF�������`y�")��I�T��o�? �h���󭌼�*����{���;o�����e���n�<�ެ��bև��m}��!}Pz�+d���Di�w1���:\����g����VP4>)&|6E�5�"L�	�j4�c����;&yxW7��YDd�r����@+?��j�7�T=�g�>#2����i�i]�kM��Х��u��)�|~���ٗp2�J�ڍ��+b��=.�D�,e��Z��L����k*�MY�R�pʐ��G�g�����(�����7PB�<<%_g'o�pV�D�C���Ppڽŉ;��O]
���QiL�����N��x٫D[�K�ar˟򩲾��! eG;���Q����J*��7�W���KM]T�� ��}̶�n&��z��o¢\��f�O�z3u*�sɤ6T��WȂ
a�� ��\|OhaXD&}�G��� ���X!��e�Ͱ"8�H��<�, !��9��&9h)��m�2��(���O^�u�t�������Y�Iw{x�L�vR0z��P��Y��q .�{�v@hpW�pOYH.S[�g�ԵXU���i3�K ����ɾ\�~�$5���v�p�Xw��J��Hv~��r�=�G8&yw�a9�S�K���o��ȵP���0�G>�o��GMI1Q��D^���ˎa�0����祥��_;z�2?碽	��|�JO��@c��s�=�&~�TF+m?%xpV��N�V�;OV�g�M���f�<X�"/�It��cJ�vc����@{ix�jw1����	+Kѷ����U��.�}̋l��Q����E��;=�*��>��c���r漽���3�gxJ������s<�siMxÎ#��%�-p���dAp�.t�;5.L�Տc'K���A�&���p�\U[�)R'�G�h�;���B���f;�v�W$D�����)ȠD����h���������@a���!��Q���9�Q��ɣ�sF+��T�0��~ġ¦b�n�(�0�|2�u���y��"y*��i�.�䥲`^�}���|��\��9��>\����7�n&�&qq(���qg������b�R=�x�� y�D�ܴ�)PYV���DI�*���l���b�(�r���C�p�C@S��r7 d���7JM����q�O<��� �]��K�S�tR��w��h&�U%����9��	1��r�M13�{��-�<���u�i�uI ,2l��U���C\�z{���T��{*t� )��S7���GEQ�j���%�e���6R\O[;�eex^���|���HS��q��YU�dp���3�xk�K`{������]�F#��J16R�U)�\FP��F�,�$���#�e�b���X����/���n��$����� ��{�Ն�I.~��˺	X�L�8\���ou�­�LJ0L��mO=���lR�_1�>�ӂ�2��Y��0�P(�<Z���y�[�AA�hxo��e�%`N��a��,�&(�dOn�E��d�{������+ŀ?~Y���BC�����ݏ���z��O�!'�4����@��oN��zTG��;Jх։���!��Wz�ඦ�׊�z��K����,�A���Zry����o�ѥ��E�n7e:S��DbG/�Ǜ�]�[��CX�[�ò8����	�n��gGz'����E�]�%��X ����/��'�b�-?�Wǜ^�0�Ѷk2q��:J�	3e��>�;�s��*�^�I[S�xڑC`���2�j�C!�(����8x��ʲH�� �s_��S�~�!���}��jp6�M{p�P#Ǽ����굽��}�,�.�[E1��|>�Q��z�?+��5�We)��	Lߦ��\Т�}��+ ���s���LV�I��gK��y� �7�b�M�Ο1%�z����'�.L��f����M:�M7M��3��5��TٛZ�0�W
�z�������g�L�֍+}Ϥ>�/�w8�>�/"����^zOr���o�eو3��C��<����.S@��WF�ښm�v"l����e�m_�E����\���_��^p��K�ŷ�|�%F����^V�]�ڼm����h����������:������Ȑ+�c�p����/�g�i�������BFN$�rN�����H�˗[l?#. ��;�(�
HqK�n�l����ޱ�)�3�"���͛�6�����H��"�l֩�o!�<?J
�����5"���w�cXN5�`T�W�ņf�,X��5Y�������l==nY�� �k(H�Uw��x�*4�EO67�aMY$5Հ͐�?[:��q�!!�/*Y�b<h�u':����Ǯ��i�{@R=���&�D#�h \��,tԅa���TZ,��nH�c%�A-p�����7�	Bع�x��ݍYk=e�K�9q��[��縅0w`�Z���.��,�oD2����@Nv��S��E��Mr:�I�P��kr�4z8����:FlJʬOG�l���^�s�>	ȩ.�ƿ��N��Y�n�0l��?o���U���M��BH�*���h�)�#҈Xͤ�[���hn?�ؔ_5lqiUҽ�;���(�����V��3�X;��5��&ٶYn�$5p�*��f @�	�Sr;��[�B=�d�jE%���-*�x^�g�����({57(�T<������7�6��A1�{���y�^��	E�Ƣ(q`�����L5o�l��Vc;z$��c� ���t,/"˷�d��A?
�$���P�;3�?ɥ��]H"j��&Q��[�d�u�٧ϫ�]ݵA:6[� S�ꙗi�ۛYԮcY��Hk=�Bs����|3]l,U㧎l����������΢+��҂4�Y�\�㫇�]���u��5�Rr�Y\ %�&U$��jR�L��3H*t;]l��^�#Z��*��Qx��?����W��X�>Lcv�N/щ��kD��]�FѢ��sBN�v�K�J�^�H���,��_�b�8a���ء��Us#�K��(��ї�p᳑��ǘҍl) 
,5�*ˀ�cCZ�z���-��a��xͿن!`�`ү*C�>�	�9Pff�V��	�sh����9����)If�dx�yb��(�ϮANs���C�_g<n�Q��Pݛ�D���c��5��L�Njox�	j�������+�W����I�|�4� P�p�@u�"Iza?�*����&�H������ᆡ��	_(�)����K��Iޮpo-֝�Z�����E�"��O��a��$�#/>�co�3,���� }kI�!�Y>}���n��Eh�"!&������Orh�8��ƈ�ڄ	���mPp'|IJ��m,щ�_��q!��AI;I��&���ʹ�9�$|�䍰<��[s���QM����T8Ny n�	�?4�~xz\�P�DgWYS�b_�|I��0���(������]��o�m�B$�9��@�'6�ES�m'niF�n�iA�=+��#�&���*�|gE)�L0�ܒ�"}��o�%#E5ї���Z3iQW��gQ΃i�DzK����խ����z�O�@�?����Ux�z�gI	��:ٛ-�x�ִ��w{�Vͧ�Q���b��$Ѳe��~��,�aTRg��q�,t������v�æ���L��Y�u��g��(���dӏ���hh�
(F���Mu��4b��;�d��>}Bfe$�����/��mh��ϐ��l��Gi���x�z���
#�V�"�B�A;N�4�!)�|�x*K�O�_Emn�b%�Ҏ�����/�E���P�R���ƹ*_��a.fݧ�#�;�|@�؟b-� �ߒm���H�9�W�3� ��ub�M��w��7l�N�����6�:ϧؗ�k��͝8��/⊊��
7G�p�=��ݎ�M)����
�c^���͘T�;j�/TK�ݚ��#�()�� �Vk�����x�gq�9"���`ׂ�G����G�[��)���6��i��E�x������+�W�x��h��j$Hw�K��truQ���h�ƴ�<�'m	x2�Q*�t�'���S�Yߧ{�CD�`�*G�Ѣ�ÁI�r��ӄ���r�T�i�گ�P��%.w�a:���� ����^�8��ĐiB�wa�~�Slá{7 �Kh�*�K�B�p��˖XJB��y�'o�<~�{d�)�y llTĝf��#>H�t���ś�7�EwS^�?I���V����+4ʌ�� ��!�_g��,�p�x�|����4�-�K��1s�/�k�S%>j�?`�J�
�L��(�_>����Y��!��8���1Pϫ�H����3�^�����%�Ӱ(JK#�'����L\8
�f^� :*��IK�w�����ڹt ����NG�H�������V���&���B�X��!Ǩ�?���S� *�i,ķg�}�Y��\��M�J���Dr���yI�@3ze�X���������`Szg@!$<��98b�	����܏��M0�a�k�w"�|�������������f����m-�j(\}�q��T���_�5���ee����ǡ-v��&�?�3z���uL0w��c�� PK��&��S�W�xS�:����	��ɚ �	Amw[��9V�3B�M�����{na���ʯ��?��
������Yww{��\�bj��,�Cj�����UM�b����-*;eU�����$J
ݱ��xW�L����n!�U��������8ب@�WΗ��~T��Pؑ]4u?tQ�U���2�x��N��ʳ�𛔊�\|��=h%�]��S�ّ7r8��(��Ӈ�M>rDc��b�C��Kp���L���2 :0�\'Ĥ>ݶ�S�� �h�s�[�`�z��A˿*�n����d0�$*D;�%���_B���UP�R#hEc��F^�buL��kcz-��~�d(\���O%�W�6��7�=5O�b1Ea�-v)��Ϸ�˔��%�{��c�Ҫ($d�GeB4�n�f?-��x5C}3$�˭*L�%<�1�5�������~�(��fߠ�8 �"Rɗ���VH&�w��o��S�D��~�FY����Al����p�������,�R�����sڮ���!��;�z�Я�����"T�~���oA��u�������u�$$�����E�/�"S7��ocz6�G�{V�'���w+F]&�y�`qM�>��&ʆ7'�HaW�����#�m��]�耯?�bju/N ��⊧���Hd�j����c����&P�A~F��e����W�ȃ�/b�{À׭J�wvL���p�f	���o�x����s���g��)'T��I-�VM�-�\4ܶ]2�F�m
L�+ᕻ�c�	��A)2���m�����5a��G���9n��ݖz'F�.�b�x�v:���?��;�x��|��� �F������Τ�=��v�����T�!/����ӺH���U����n�� /@���(UZv�XPB ������t�������A���i��N����'p�̓H*�i���%c �$%{گb~�!���[���f ��q��^����{��>��+�ӎ̞������o��_v98�ܠ�?�������\�}�%��	vGU�ҩ���$�x7��1�=�6iz��W7��hb��=�0ka��=^���Q����������2�16��3��	�Қ���=�	���1�m�p�Y{H�iL6�?��2|5Z�� r��`-�ryi�X.��8V��Ao�:^�HY�F�EgQl!�cm��������sB�����F�ac�3p���&�Is�4�'A����߉fڞ	�}q�	kP�x�y�wq}�^�d\{B�SBD�}Ĭ���7�l��G���k�jԴ�ͩ*���2�YK�
�;j��ʝ@����r���?R�+���~@-y/�p����h'�f���_\c�l�\�,��W��n�^�sU	�R��n=y3܉F�g��Q�Q����vd��5Bn�;��d�A�����OI:�4��`Ԝ@�Ѹ��xAp�K ��9$�e&��t�d�;�z��#+��S!}�o���Dn�Pq�(2�{T��]�#�-qP��SW�> ��zF�0D��P4�^W*�A�k��t�.����%>Q��'^Ǚ
�2. %=���]�n��/�H*�a�'����ïƉ��G�+ �]�f �g�}�A)7��J�/e�|�q-��� ͇�x�و�%D�!��(3�*��,���EW�����ZesM��	�ղ��8`���F��^ˎ؉NAXd�ۭ�HY|Ik��g��3�;1?=���́�G'Gx�k�5��������^'�j=͌��`S'3(�Bł-��;ɞ`N��{=���_�����o�rт?��yG����9"�b8�L䱖�����m-���w�,-9_m��A,�w��7%�i��~���`�eք�hmx�6e>�+�S��c��XJ3��b�� �4�){43"��ɝ��M���d��ax�N�^�����HC����4u��d���� �u;�ۧ�J���:�)X�H��mJ���%�#/�	Na����z-���#���y+�K�l����д���N�K����Fj�,\[��=��>&��}2<ݣ؏�R�x�x"��Qd�w�3�#��,� ���An�l�"(��Q=Y�&Rr�	l��5��f���^#ż�� ħ"�B��pylľ4N�i>�0�z*�..
��>�Mt�k�+(֯�m�4C֯Su�a:p}[/�klt������֣Q��'i�2Lb��{��Z����_w:���7蜡�R�K4��!����R�Ɖg����%/H�zY����4y�:=d��}�Lܵ�IIF{o���qDE���ެ��?�����>TQ�Wä�����8��(�6�k�KKJ\q���*��C P����Y���|��v96�N�Z㑨sd��``�[Zo[�y��.���3q��G�nj$ᡤ��c� ���^�+
>/��Oc.!P,<��$�
�m�3Úz�l/tS��埿�3�M;�g�B���_[��2g��KXzhK���ȗ��ǯd��hô�b�R#�����CAa��O%^@�<�d3W�v�t~�b n�h�~�]��Z���({��ouȝ��~~�:�C�$h� ]�2��{��D���cI �b����^:�2��xp���u���`з=>