��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D���F�Vp��t��<'T�z��o�ބz��{�s�C�Dp��-)DC��l���%X)�by1���:6�/+TV[��i�b墟]d�:��Oa�#mK7����ZT�+�`��Up�ZZ�wC<H3�ؔeN�r��<-�^��p����b!�7����t��lG�pـ�\R�����Ǚ�0<�r�D~�X{D@�x�uF�
�iY�5c&@�ک��
�#M���)�N�w����S<g?7-�@�ٕ�[��p����lx��Z�d-$d�-��Sp9 +��5Qa�<~�V���1F����� �4�)���2��&{<����: �`0Q��2.	��CX���w��CH5rP�D�<�r���{\��h���a�ө�YDƧXI[�d_�pWA�������]�k��n1��>ͥ���^=F�5&v��I���J@^D7͞�E�$V+O��=�}���xܠڦ�E�����j#�q�|�'��)HJdV��R�_f[sWgL�����y)�"5�ۜC�{fᵍF��11$��g{Oc�&�"�]���
��A�k�S>MR���܅T3A%4�lO�L��.��_��Ɏ9��;ϙ����g�h�v�RipTIB��|`�\��q��0�!�Qײf�2f)ְ`~S��1~G����E�aW׼�4������k�*Q�~צ~��E}]��t���*x��_���4�*_z��-��ǕoP�}z����VFʶ����T� d�CP��5�D�me] v0�AӋ[;K���+�Ӧ�E�SjG��̪u!�3�t=d�t�7� \�����]\+�k��JH��[�=q C�� e�Ǭ�Ē�aA�o�mIǫ�`����}���W����kf�$����В�8o#�^(=C�؆��0h4�7�L<���Up"3/�'�<��Կ�`��$�d̃G\�>�4�#�mܡ��>!�����4P	���kt_�a.�"�?��{a��_�
`�J���^.W-��]��l�m߳VE����Q��:�+�Sd2��֦#Ĉ�CI�t�=�@��0����?u����q�����35��.l�Q�=mQ'.�ԯ`4$�[��E�|
ƴ�oFf��Xw��[5@2�� ތ��Xʟ2�Q/_	��o1v�ng�5X �cު�|sE� �{��\�=�2إ""��xF�'[r|��#�]0��H�������8�G��W �~$x�1�hﮢ��u}[Ո���غe�����1�f+�R$>!dT\>'+���=�%��a�,"�sǤ�a<Y9����e'=����_�pr�V���b5��g�8���6��oAW:[k��w���e��gڞ[0	��6E}g񲲞�k"�\�K1iPC"T;Mǘn)�<HY) B�����P�?�7�\x�!cP;I��U,��-����c�p������ܣ�~�7	�iF���a~�>驻�����A�
'��_�E����-�'=�X�L�r�t����(GP�ߠf-F���:�E_q���&Ӡ�l���N��'B0O�9�>t�)�2�3����Hp7L�pIU���P�(s��ŊA�0E�~6�N)�J���%�:˥:�FmR�>&y
\������/)!�9��d�Ģ��#'d>8�+5�x̓g����,�v�=����(��^�G��ۮ�tFn���a3��ۻ�C/���U~3BWޢ�g�*���B���>^�^�Yu���=W�*�K��� q�vl\#��]��"9ϢXIN�(����ߩ{p���A0�+5G8�]e�|E&Teǧ�k�{8I��ІV8\�����'�|��ݥ���oɃ�n�h�Xft�C�&�T^Ne �^[�c���o�ْ� ����3��*��y�q[!��5��Ԕ�a��o��#�ׇ���(mG��>G�٢w�b�c��La�mA,^ŷ�>0�V��hX���7%sg�Ba�Yġ�Z�e�I�DߞQ���[��9H��J��u�X�����bs�������A�%�K����	l��(m��+�h���*�t�I�x�XL߳I�,M*Sy�X[:��0�� �X�O�i%�����U��y���O0ڠ�Y�t}�^׳��	%\�W��v�g���6%"�o(1|beRQ`��}U��ݒ>���rm!��i~Kݦ�Vh������:vB�FZ��Q&��56H��A9�2B^+f���H]�����,¦Mh��H��?��6@-�i�ѭ4����f����h��j&e�)U� �<���T���+�?;���zT	7�;ZN�*wND"5����U��D�^��žIhܹ�3�,�Q�����wh�-6O#��N~��/�C�(,��r���R׽g��g�N^KB��5���@�ZWX_
��Ŝ�ͨ��';j�<���R^4f�U{~��r�t!�0�������Q�,�W.��(���_Ktz�mYs�+%lm�{s7��E�줨��?���!�5�+����x@��4�_�Y)CB�[(zU]���YV���fѣ�ќ5����}��i��=�Z�*A��W��#7�ݰ8P�W�w8�j��ꃡ�H�JH��P6���>I��MR��/y!��DaP8�V�W<�$�0��0FF|��a_�"�چ��x�>��oK�7���Q�9j��H��S7��,cgH4��㘵-^[\�k\`�h��3���`H�t��RD
M�u�h�ҧ)���H1)״̣I�����4Nzz��ɶ�*w}�@kx�٣ f;�UT.U|����q*wC�B}��k��Dț��qʱ햊j\��i���Ӯ�S }�՝���.�i.8˷�I��>�C9v*�~t,<�`!���e4��hQ!J��q�4����Z��ʛ�b�D;�*a������4k'�8�� 1��\((��q��s��`�#3��4��ϗ1~�t6���,d1�4���I9W�>n+"�E��%v��n#Z��n@vl��t�}����9�s���ݗ.��r���Wɧfˁc��w�\�#I�Ϗ��9�,��w����U�dC��PC,�`~�#x@�ɘ��(w�02��Я�)!���q���#����Z�-�m��E8E�/��
d[�,��L%Y�J�S{4�q��%>~���3�vv$$u�۷!m����W[h�޷�!-Js�	*�� �ܻ	����@�q�U���C8?�,��^nSD�D6�tB"�@7�	�E�A*G��b'7�r��Ad�����+��ހ��-�cՉ���'i����W T9V4���kِX��E��'�� ���X �T]}���U{��W�'&}*ܵ㠫|v�qO��CLh�p>f� B�v���o@4����)�2����D������T�����kĤQ��hγ�Kđ?�q����M�tJsc��sƒ���GWt���Q������@̪V���3�.�-�;��4�1}��=���˃�1�f7M
�P����e}m�9;q�F6��M֊�GK��d�(����*�Y��Z7��±ŝU�չ�$iqU7���F�����M��8W�M���>��&���<�?6^n A>��������rHfy�M�QzS��*;�B�ZP>��L,Y��%D֛x�p{U�)�t���m���j�`��>[ �ы�0��G��ӎ���ܻ���H�å�Oi��;623/����ѯ0dL����_Ϥ"į}�%�6�.���̑OI.���|>.�\KF�W�fro�fO8K�g�|K�x��%V��L��ȝ�=��ZL�T�*cR�Q/ ��q��	D3=�Iu`嗺��z���H1��P�k2ǋE߁|��$C5���.g��b���P.o8��)�o��\��yt�I���-~J���cW�0e}TR��mȍ*t�6l��H��.�{�-
�i,��{"����Ǚl<��M��h�V��fFg#x�Ȕ�<�_���[ӓi�����Y���ڨH#���#��权FL}�Clе���ۜ�p�Ϣ�Z�����ժ}u��9N�&7���;ҁ}���գLzǾ�ch:�������%Q��[��Z�������|@��7A�n�&*9�#�M,2����� �h�l?Ln����Л���ʄ�q�/���=��:�¤��S7�"���K=!iw\�t��OJ����϶3�)�J�d���Zq2m�|���3��?>>�|s��,����B)e��%+u<�3?v��_DS��"���F��c�@�Ӂ�E�Y[UK�gȱ�kVX��y7��"!�B|���9WT�5�ͮ�����#e�(�|�jے�(Q���d#�
��wba��r5Sr�`s=Q ���Pfx>�5�d(�J�tȱ"�Ӭ*=sa�¯P<�)3||zL�X�C;?�۽�o�.;�9�r-����}�T�����U���S'2�I2��1A�929&7�Rֲ|�C����p�:-�=�D����])_�W�+2Դ#(qˣ�A�g�.A�	�Lq���,N!���^�n�{���;�:��b��͵���[wK�K䕓���m_Q����dg���8�7�_��Hx�e�L�e(����
i@�Ϡx�1����Pz��H 6g$���ex�_��%4�Lg�����+�Н�(�=�pR���>4��[�z|�ƒ�P~����`�<򕏓�=mT�?�ѡ��g$t�%Jȿ1��-#7�� Qwȣ����ߍC0 v1�4_U�K1�W���F��N��o���
�;,�	\BGĎ��<W��> 7=G�d��8B:��i9�#��K�]V��6���g�E��W���5�� �C%A�N��L�M?DV����)-�
���,�N�s �<A��q_��.�C����HEO�ͤnC�&��hM��}p�Rr�K~����0@,A�R�p�+�n����={R85xBb6���p�.û�
\�~�0�� ����h��T�SĞh/�Z�d�<;�!�j��Ә�[��FH<�� r� ��eL^Ģ�\v���m^�tt �!���ְ����I����W��Q�6:أ^�QqȐG��Q��� �8E����ИH�d���pZ���~��M�s����f�s2+�H�ɀ.A���%�ը�l��6�?u��v��/���0� �7�]�xl��)ei�޹+�Xg9[��������Nk#J�������9�KS3;p�6�X��dQ���1`��5�(�1(˨Vn�6(v�z���N�L1�3wM��fɣ*�)IΥS�Y�P���_�z�sc+��Y�Q��������_��zEYr-���dZ��ޅ)�&�/ ��\{v��InN�
L����`\�c�Ǐ�o��͡��U�����i�����'��l��/�} J{!|���)?���o#���95|&So~���&����S;
�(yYpR�p���p�*+������+��ՆR�zE	��#t5�+����l��d��
R�g��v���t���R�:�����']�+e'+�Kf�6|_@�XQOD�hA�ִk��
(�Z:�S=#���[���u�+���/�:���'r��zK\
����Օ��[�s�`�!����t�yڢG��,�6ђ��s�z���,UV ���ڨ�2�\�*WR�Q�zor��F�n�(�,������b,�rH�~Re�c���-��ҒJ�+am7#�/��3�ͧz'>�9/�\�W�C��$<0�����Օ4���M��&.~�n(�X�ǺoI�Mƒ4C��J\��C�-̛ڌ ��k|� �R�a��*�9ك#�aAe�K������U�������b�zΣ����-�g��z���PR���K�zC��D�R\7}_��9Ԑ��%u�n@2�D��:@S�&�o�G�vG�C'�)e��҉��m���aAx�k�hH����(*�9Q���V�p.ʓ���$EC8�r2�� �xU���EH�-���<|����o��6ح�mP=1�h���X�&�Ja�"���j^|��q�U���+�jL�ڢ���DFD����C�� =�l��g�>PP�,%�:6�o��f{���ҳ!�sY������eE0��{0���l�엯
���4{��0�ݍF�	��u�Cy�����*�7x��;w4t���wqE�+�>ۮl�=���O�#�	�-����a���N�_�\£TCt*M	�饻6h�i�&BϏ
�'H��0�c ��k���uE1;��2;��ɑw$�=R��[��	?������b�����v��iM�>,~Էh��Q��lV��E���5�s��<3_�2aէ��C�T����e�~�ج�Z픐v��}ξm�4�-+��j+n�^2���'F�S�{	"��!��x�v%*�����f�/�Jރ�7�kK������z!l����Z{uO��@!<���B�u�W��vF��k>%�8�Bj����Y���h���3�9[h���I���5����x|$����@�� 5�e��<l\`�蜟AR?'��7��Z���VW�D�-�>-���Y_��B�����xc)ǓD���J��b'�KW�c�Y1L��T�Q2*�j���l��.]���I<?(�1bOp,�oL��"ql�_J�;2�"c";�=����(���Z
�_��Wq?$ �΃�*^���#�U�uG��9�����큲�������o��1ݶ�)���s�}N�㚥�bq{F���KYeԮ@�o_O/����Rh���Ɯ�����=T��z���2��E�s$�������`ű��>�lV#+�Z�İ��x�����w��rc��Y(�H��`s��=o���#ιp�5�C��h'V� ��2�?O0�qsv0��&v�+x2�<�8?�%3�����T�<CogB�g���HX���:��T���&R�8��M6L́������	0�mTL��iK��ȉZ��Y�5��ڣD�q��,�!��ySfaG���F1�]~�S=����C�������{Kǎ(��ڐU+�dU���9b%��ݰ��U��h)Ŧ�?��:��Xe���L��H1����p��!!��� � ��l�Ft�C*��y�~���q�J�xp����?c' �>!���%�����$WG�|T����48$[�!�����T�i� �!ʥ���dJo��k%�Q��|D��k��V��-���`�:�|�G�	��;�@��e�I� O$E������'��+}�ײ0D�.X�)H|
bՊ^�L����d���U@�~�N��B��xI���^S�̔�d8#�](���̃Y]��w
��v��7CkŨ
�����#e<����a�Ҙ�=#��C��"��lu�heP�M{ք]���Doc��0��y���1*p����b	vг�������ZW��O է�`�(��P!#�/��^�^�`��?�@�$QQ��NoŐ�D'Ix>?���~&�МZ{�@#肧S$��[-�M.�*��i�b�pYq���=!f+(�k)X�K�����J��&4�]�n-�q*Db)��o�UQh�]�R �u%�l@8��7�T�w�&,`uF���/�s7�h,���]��-h����D�_Dx\4gi��������َ��4� oo3K.aNDM&��Ax(4E��_��{w�Ay��fUgϦ��Z��%����;��~�P���Ó� 5��
	HG~X��\"v�����`UE����ۿb��O�<R�k7�J6m�ٱ :�"�5Ӳ(�=aZ����4d�����y���ɸ,a���� ��a��	k�d��%����c+�A������u�BKD �r}|�i��Cd<�o�0@\3(9mtt�lD��,�y�P�;�8F��|I����q�Η{�fƁ	����8����!�t�,���sN�D������IR)NA��F�-��r�Fk.Y������퇷K�Pu� ��.������9g�8�Y�YW�H���D+!s��_��}�$�{W�4hg<E|���n����4��܊�]�/�X�����K>p�5���;o��s)�˒�K:����",�)����(����q��h�J1�1H;��������A�a�D!�_��^Nߒ4�I��Q*^4#	�-&Ek�5��<Ոۖ��9جݖ���u#����N�_[�3��]$�I�����|�d*�oxor�@��/�i;/}�t	:�_k�ߏ�O)��"���Aޓ5��o�~u
�e�� k�62F��)����F��~ ��(k5ڹ�=�O$n~���9K3�]�N�H=��p���(���~�]٩�^��Wq(����ɔ9ZR��e�R3��՞�~��aL�̋����+@%�Z��[�V��/�r�ۙ�!�R@�����Ӆ���u�3��{�H4AU����'1�ihj���^Q'��j]����5�̰ky#4L�K���mH�Dt?s���V��s��]H�����4��ިC���/��[7j�S��.�V}�=<�W�쭋����u�i9������Ì1{J�;�<������z�$bm�n���W��,4Yz�P����FC.e�؊�U�kǥ=$q�:)D������Q���BeE��	I���h�Ip���VO^�Q�M<J}�7����Ԧ����9t}�r/���,���?� Ŗq���]s�cޘ\�C$�]p�
�J�ꖞ0͓'\���=}�]�҃#�l���}��[0�^q6����d�K ����;�i��Z�_뛵{q����n7�!�M�8d�Y�(q��b���9Avu��l�Ц|4"�~��q�{�B��>&������]�X�"F�;lWDJ��J�fb2Υ�eU�ک��N���j�+^\UF��h�)
��-�7�'�~���[h��6��A8m'��/��ҕl���A�d���&c@À���`9�G�=V����2��bW!�$>��`!?�%`n%�� .�������?��?�d������d5ڼʷ����W���cg�6j_(�1[YD6i��΅����b<m�b��|��Q���U�yW+��/�j��kY��Z�x���[ucm�c�be)���P��~�-��v�8�攂0*Q�����×ƅ�>����|+֔_v���=����8����"�� 5���ó8���>y@n5qW,��C"r(-ZR'��s*�B�`/͇/1$�`�,Ef�mA��9�p����F�x�9��_�c˳;��������^��� }���c%^<��R؏]p,��4�`R�l$�b�ӌ�O�f�q�X�}*x�M�%Y��� ���凎�s�`{^L��o����-�aU��jXR��jX�{$�J��\�N��A�&�I��+�ux��B�3>�Q_�D�?�Q�2�ē��7[Nca��R�4#^t���c��t%X`k<ߥ��	�.�(�1��c�p-�|)�֌�=>��G�u���Cix�U�%��a��)�j
���娧�:M��tIR�b)�������Ź���g� }�M�9����5�fۊ�ڌ�+."(
}�@�z���ܐ!2�v��c���|��5���Z�� 7��dv�F�Ϙ�T
�>
�L{	A#�}Ŏ����8FE���j�
z���rW� 2/F$F��
7�F��KWR�X^CL�?� �# <��w,��rbe��}�+�#���x�i�2�H���9,��"L*Z]��䌆T5�5���v�r���Jҵ�_j׹���z��ԼܒlBYk������ �a%�6�U$���\���e�����,�ޗ��'�Oƅ�}�+}���-C&�N�z6/P$���+Fi�j>���"��W$�n�d��
A7�:��Y����ji���'w�!��K���P�0��`#�صB;ݨ�2Aq���]dķ@%Ĕʢb/M��B'�:��o��3B�^Y\�:����ׁ9wp$�kʟ��Qt-UZS�ܗ�/E�#�G�,�`�ѢO�iѺg@^�e�ݭ�j9kC�OPk9w���N���"���>��(&�[�Y�"��0T;(}�vI[+���_af�w;w�ԣ�E��RVf0#��}yN��2��u ,�y��oOP1��������W�.��D�3��!�_�L�L� JE	��-��$W�ŵ�u�U�9ֶ���~����E�-s���2~w��l�.1�1�McN�2�"��9wQ<�B+W��ǨgO[��W���#u9��z3�6��{e�ҵiEt�9����������{���K0�a4;��¾5�X��C���%��K�Ѻ�ˍ�Z�D��۠7��!�=��3:�#ɓ��v�9��b͏y�(K_S��g��2f�b��Z�m%Q��,��}�)u���叨��b�c3.�G���,z���/i`
� t���� ���	����Dl���v35X�F�o��3����2�z�j�t�����
J�d?s�b����7����6q4���$�aO�<����{@Jc$V���^��k��]J Uz�:Z���"z`u�2U&�_ƶ�w����/��$	uSV?7d+�C��@��u��ڶ6�3T,pi�]�M����y�>l+bRH �B(2z3jW=	 �=�P�X*M�Q���O�ol_E�y���G��$��U�!h.��m�.�ݰ��lb�?JĂ�pE�:�$��W��zz�w���1�Nv���;{���i��I�W��LjQ��؅^�:�gӠyԃE�������G�"*J�^/Ur_i|�Nv�U���|��Uv����l͋6��p��/���N	��
�*�W��t�kW6�ij��.���6!�̻�f�rS֟4�Ղ����0��#�c��%��}�X[����O�!{b?�4�N1g�;�[P�������+��;l�Y��}ɻ^|���,�A~�}4,�u��+��谲� ��(#�{���\t%��[`�$�>@GB�wJ,�����_�a�y�?�2e�0$?�c5r�J�-��w8K���\t%+����q/f��i���#�T��wǶ\��Z����s�쾗�x"�v?;�
+�vE ?]+�`�.��?R�{��R]a�E�� EVk���]��y��z��9>�+�fо���e5�,�~%2;jRn�8ۚ���/����ޕ���w� W+�s����l?�S�mFO�F�؃���@��g3%yΩI�v�F3C�����V���鉹�1��
%m�y/�;�J��e*�y�sE���r#���u�]�Vu�J�C�#vCV�kx�B�� #�,�Q;��z<#�M��O�8>��6��YHòk*�U�/�!���H"!!�jn��ЋhJ�i��a���Y��5Ӡ��H1�
h-~�;~���+�E�����I:�n<�(�倢������p�6{V���<սb�r'8"4P��܏�|w�X���Wڼ�,�D���L\^'�^cu)-�|6.�ܢ��ݙ�6G�A.d�GS���sRx��nr�W��)b�'�]p*"����>��!@��	�<�h_?��5Q�x����8c��ݫC���U[��m̐��h��X����*�w��S���� �+�G�Lb�]<3�|�%n�8=ƒ���[�wv�7����G��}��(�&��£�C�d��ι4���p#ې�H�7+W�_M(����R�Bd\�g�-�S}6�@�-�2$
?_�4%[g:jl�5 �P���9ZASh��Qp�/V^pa����z�^����6��i�� ?��%y���Xy���ٜ��m/Q�:�W"�%� ��8��W�*g򟰭w��ᷞ�׭�+�d��c.�7��f!�Į�*y�f��w�pRC���s&�`E�W��(?v�~��U;v�8��@��(��CW��voV&��MnYs��ʵ��tr$#Z�\s��Hߪ�	��'��K�ǻN�������[}k�5y�L%o,F2��_՘u4+��ٚ�1����ϻK>g<<1Kb�|T�D�~���r�fg����=�'�R'D,���[�a�7�I��ܢ����ʘ����S4�54L����ֱ�_��渙�[)�-t��V�<dΙ�>��nȡ̞��1���B��h80N:<��b��Q8��{�
&��"F0��~�c!6����6����C���ͭ��N<c�'�;�@�T�sp��1�sF0/> ��a#"�*okio�
DgW��B��֔̚7�^Et$�'(��0zD#îa�Z!�8Q�f�FIO��e[�È@B�wޕ�;���;tb���$���*1�N	y�-%t�/^H�ղ۾��`�P��2 jW��F���/fMm�����B�v֔�Y¸1�$%�Kז֒o�,Ǹe��Mk��ҶϳX��2U,n���M��y%��)��q{#��GQ]���7� �� A�e����KM�GPm�h�e[��ФaHL!�&Y(��S��î(����dw���֘��ҕU��Nu$]�M����~�ޅB��F��]��x�����S\�9|��㾌)"�eo�+���G�cG2r�wnlj��D�O$'\�����޿O��Y��q(�����n�	6΋����>��u�����s	w`�*���I�7����+��*��	�|��8E츾�jc\��?r|�]�N���6�u�x���&yːzKB�����9��#����\z�y��T)	н�|D@�.� 9������)�T&��圾�m�T�ǜFZ���ާ���5����x$�n�x���#��LV�]Tt���3�S/�j����)F��ϕI�hC�zZޤ�����~����o�����g�z�����g�sq��4ʧ@P�.;d)�]|"lBzCY��Z�Ch>�?/sZt�;<`�f� o��8C]93n5~�gb��d�h��mI�0����5��rS$�&`��:&,Ͻ
�������%��u[+��-�	�G�a(J:'ԲO/�o�I�9a�ͥK���מ�J˒{���$�0;�*��Y<��֫FMǯ�9�y�.$�ֱ�#6�҇��jβv3Tc4��]�n�#����6(���J���N�c��~W���H��r��Gm��R���WR�Z�����ԇ�쒪tf�IN#�{$S7a!s�k�օq^z��5k��4�'��=����:&���&�	4���k�M�����i���Mn��y_����3�9��*�N9J[.�\�c���UnSw�L��[:�d+r�ዳm�Qb+�V ���T����s ����
G���#��6Y��rmB�b�ǔ�g��88����"gZ�۲"�J��t.$D��,��)�	��&��q�ȴbş����us$.��8Q�/�s���w���OJ���p��?��y�d-n��O@��/ֈ�T��Xg����P5y� ��>i>�"OIP�,�E���1X�'a�� Ӳ^:(�D�c�Hjé����a��/Wh�k���dP(�9Ã?�5��N�V�b]�"�->�������k�IN	�i'�mQ����|/P߾�y�:3H?�E�kw���+<Ȩ�j?9D-� 8���Y��7��`zU�{1���1��~�*�C�#W�Pc��I��Ȗ��h�����6HpP��?�e׎��`9x�f��%ޕ\����?|0WM?U����)������ �M�8^
��r����W't�{���*�\S]�-�v�E��h�Bi8���<��5��L�6�uXW�C)����ltϠ�� �H���#�`�$���XrQ7'��ŋ\��k�	+�xT���u�z{��K ''et�ץ�pRy1W�Q2m���zd��1}Y6���c���OɎ-$��9B3r�$��XS����Yk���:*6�I�C ���o�ʪ:s����v�s�%�ՠ����7�����\&t������g��A���mf����?�.`�]��⪻C_���� (�?��&ﻶ�� !N뚇��'a�ov,���~���c���H���<�f��G_���Hv����d�`>�ќ�������Mב�7�\S�����JY^$�rˤ��'�N�m�}9Ӷ��Y/J<R�ET�VMh�M����iǲY��3�	h��D\]��g��������Y��Բ�L�6O�<�$��3Ӛ�;(�X�¦�U=��˅���(��GO]��.2��#yj� ��]JW�s�l��������⭶��v_.��^A�eX�ΙWy��x��[��U�����/t>��ʋ%�	���'N��)�e�Qq�#$>�`�d��w]�%c���0��D��*��d�&8��C�T�����eV��H��nZo���H'�4���w���K����H�8�I�3��T=<�@r����JW�$�D�&Oggg�0e`��Յ�uD BF���CU��iaS�3� :w�p8�Q0S�q�{6�cS���C�t��PɈ{m�c�O��0yXʦ&:�P�$g�x��,e��z PE'�͡!E�2f�N��>�o<8~?ΰ6�w�<�p7	�&����e�yN��ʨ7|ǔ(��d?��� �e���&�,�q���+������⊀-N�)5����e������8c�N��Nei��X`Ԟx���1�՝�]����?�e{���n���p�>h�Y㣮����
���M���}����b�.3�=��7Xl��d����l������.����;Z�I*�N�'N&��m텼n!&�3t�#;���}׮P�iHFd*��\`x֊�dM�&��D�NRNO+�t��"���K��Rc��n��Yc�=7Ǖ�:�QT`��n"���*�_�Q�Z����z���8J��o8ڻ�;g��N�8R����@�h����2(�G� $5JqP��)���2O�T�����i����_�j��J똼�)�ۂD�G�E$d��MW��~�U s/��}i��/�T"\��B� ��鎔�L۸m�#��H�P. �&&{[�9ĝkMbY��]��v��ūW��*�F���Z��M�\0��;��#��'�<ǵ�X='҇�M��|���Iv<'��Gz1^��u.<�ax��H���ce����7�^���(4�_�{�>Oĥ�V��a�U���V��y
�"�<�"1)�hCd�rN�$���OB�;��J>��8��r����c�Q8�\�V=��S��K$�ġ��\z%���m3�����gbf|ɻR~��C(�V�\ں?�*���o��n��3�`��?���B|�E*�Cb���5T��sڄ�Lp'��	yb���1Aʢ0#1�[�ݎ�5Я�����j�M@0	kEĿ��<{�d�#��X�9CI�Q�9j3�|N�s�Q龇�9|��b7Y����v���?:�����Մ���gl*KU��pWyz,M=�3�x~�M�7��c�u8@"qe�V6�u=ո�}�����o����Ei�G��2sZг��u�C?^⛩\ѿ˳`4�7��B�F��Ϙ<�Y�,7js��,�!3�������m"^ш�`Y�n�f���1�ĺ�XvF�����)�Ђ����z��;�Ď{ɞ��;�_P��jnAD-�d��&R�|$ԃ��j[���!��xܜJ�?��p���u*ΧW�;ڻ=:j��ק�i_�����ݤ*�Ck�
B������Zs�%����Cڸ��$��KBV^��w�R�tV�g��""����k{Z����E�(W���)�g!#�}K�x��Q�~Ѫ=����d��E��z#ʊdt�� ��7�R���L���,����ܤ��J��_q��T�q��N�\��$�'1'5�r��7�� ���o4-�}��mq���5���kN>�d�����z+/6��XT��q4՛������ HaT�3�g}3�W<Smd{Q�ˁX��s�ߌ��e�֡#�Y����<�ɨ����Q���pV��b��erYv=k�v�8��<ݨfr��.������(�u����,�K��: 1�����WǳG�Ÿ��Kv�+�������O2|:�r�ZG�C��F(���"iL�P���y˫3Y��/�<8?�0�d|9c�[ΚC��Vz�2�Z>%��P4F�B�͹+�d���&����q�yLYq�mֵ�1�l�a��7�ޮA=���Q�����d�.�8���
� �1����n����\G3\L��3��+,[�{�q�\�Jӽ3�-����z�T:g�y��u̎J��VAO�K�g! �������F���R�b�+2e.�Ma�U��ς�{5|�7��wh����[hqR��c��3�U���X��'�qI nt�<c��-;��U�;�̟�����\ޗ�A'�%�����>S�q�&���4�7l~7�G ن����E�����r"� ���[�@��?dNU�yWC=�h�:����u���7^����A�t�G���3���q���� ���V�껺������f���rfY���-�p�p��K�k���:.����Gj(��y��E��3���^�e{�(����ණ�0�*�kC�j�u>�hJ�/Ho-2)ze���F;�]���O:���H�!�'��}�v�a]�]T�S�\j����D[�j�Y�D�&�A	O�V�u�)ũ VYqCډ�r1�h��G���9�ԱAjY1JB�������=��MN;���Z��F�%����5����p��f(ީ�\�
�o�\��]��,ĩ ��rS�(L����}�[��E��Bpy�[��T*�L��θ�5H��[�|�1x�P�iN}>�$��X&�-M!�b�W�q�Ď��'`z+|�
2�ۉO��(�z��z=���0{�&;�X��.��<+%�_��b���븋y�Au��4�����U�&l��K4��#vI=s$n��Lw�>[�f�+�����
���v���	@_M`��Laܽ��,#*�:�>U�'d��enZ�2�٫��в3%�Mү{�}P���ջ���ٌݏYLRM�D�)�,��L�w�]a�S�B���V�{}]n�`k�kra3qF��X8+0u�|ZPo�w�����OA�8<���#Ć ��;�TS�c=�A^�a�]Js�IP,�	����i>d���>�b����gV�6����~��Oؚ.t<_�W�+����$�e���SY}6��|c��k^��;�0��c�5���\� s�]
y JV��ss���^���0�[�-zg�E�'���%�$6����7�e���٧�8����R�
�[S+�t+�\O�	�i�q�jĈ�NA}����,I$,��f�Hv�;��7���uf����Y	�J�����o5!uUgȐ41��_u`�&K¬$�<:�Ӌ�3�ma���w�Z3k���Y�/a<�]ɐ���*����{�� :'2��y��G��R�FC�Z1��5�r��(x&V�W7)�K�X��J<�;�۴�=1�&�JF�(��L�%&�Yu3UH�����\��������^U���Iq�%B<��.���ǉ�@�k�N1�Z/I�^Ī���S>���>I$
��׽O4�g�?�
�cP�|H���^^^�}딀�c�0c#��z�e�#m�v� {�&%\1�im��x���k/�%��� * �"gL��M�)ʝ����m�+��]n2hf��s8��HE�������1;�چ���m��B[��`~��ɗ<~�1��*Cw��!��i��ka}E�WN��\���g>ս��l�I���o}>W��9o�5���h�܊�w��=��7�΢В��MY����=}�y�lA����I淪H��u�A!�&�?�}���,�6�^�U�r���6�ߝT�9���i�3�M��{j�5�L��ξo���o$��AdI�D��P���s\cR�O ��Fk��?b��W߾�|Vę��:U詘���g*:*����:�-�<lz�����FI����)~��� g�}�6�T:�j�P}sde������-}�GQGC�^1:��GZ0�w�Dv��C�ِ�č��t4�줎�\����d�m��PLK8Jp�V���[�)ZR����X�z��>��Kn��/�~��4X�����Z�8���_�RM�[K��yF�p�
��Ո��<�� �sa@�P���c�t�����q�����W�u�y����y����R)��MSh�� �S;՞���Wr
�1#D~"Ɨ�PW|�}�T ���Z��$ZN	���a������WH�uQ��&.�_$���?5��ݖÕz4o��)�1�xm����� Y�,�[1��u\Z�1���z�"�U�ޔ"�Zz�(��@)�#����y+ kJs�����K���Z��^;�ʶ!MK�4uz�{��DYV���"�ڔ˪��Γ`Y��;w�77��6��k�_��^T�F��0]��^�i���(�A:�zf����w���3o�Sr�.����{$X�Ḓ�!� d���%R��҆��29�J�����0j��H��m��T�$��;���"�c7"�)��^7�~�� G*��I��`���MB��O<��j�CQ���֌���D����8-�Y�4�&�]3C�;�^�5K��J7��Nzn���Y��|t�+�J��w�f����z\����u�z��䕩7	ry#�����5|;0���[ܪA��w����,A!���ʑ����!����n�&���,ڋ���J�����oRTgd�Hz(�E.����P��q����gtFva�mF����5v�!pxb���g���S��fX�'o��ie��A{Δ1]��N�p��G2G��j��`�3���i�a�������^����&!*ͧ-n#`:�ض�Y��ֵ��>�~����p2�&���!m�9�M}��S������ε�����<@Ī��K<ܧ�ͤ��=��4�3���tO�~9�T�B�[~��&! �W(l��ϓs9�RR��Z��R�۾x�X�a�R_�j�ցk��jȔ;�Md.�\�%rm�Eha�y�.�:���:��w+��v��-F�lf%+t!b��^ū����+Xd,�uU�"'��+X����5	�[|~�Y����Z�L�r�{�t2�������`o�����p����+ݶF�Y���[�ʹI�����Ճ��k��k�y�ʌ�qm��ԟK�?��L폘�C]%�?w��̑k�M??$�f��s�m���X;�'���7ȧ�����<�᧞&L���o�OZ���M�K<A�9�{���q�!\	��S�
0�z��>�HJr�>ѩzvt6��l奦S�G�ԟ���%�f��(2����R�:F�Tc����� ��c7Q��csP�	4ן�Ԟ��ЄD_6�F��ӚHZ�R�6�r�j+�;d!7q�"\�=��U8cV�F���k9!D�v��Sv?�l�"�!����Ȋ 饜.� �l�b��$h�x|��lf�	샒�s�'����qj+�y�d�fsCs��8�f���z����%�4�m� ���	��u�:�q�!$�sc��}�3�7�C�Јk ��DaBi��y�����8������C��{�5j̺��x��J$����qEO%g_������ĈIY��e�/���M�L����[¦e�,���^���_��x�h�5#僚��W�����#�x��Q,�K!�zY����^��ι�[�����6�n4�j�ȓ�(��;��M��4~53&e�1�;�Q	��I���vF_���A���i~$�P�����4�(���-(��
�<�^�����E�0�B�K���K�
� �b�;^IX���K*�_å��f��˃|���K֢����B�ѧ�9d�]X��w����m"�	>cѧ��a�>)�$YȼH�^g�/�X�ZW�`]����'�Ü�O����lq_�����c0�A&�^M��W��OV@\s�F��3&P���`�`�^�Ќw����ʮ���5��&�Ȩ}���
��-�չ�����-[�x����'�bЎ�wr_0t���C|ȱ�i�qW�����Hؾ^L>�Έ��]]�(����'쏻6��[�1�U,Bgk[^ x�)�Z��K�+�.\jG��n�N�N����kV�<�ը��ԴK������DG�tP2�+	����q1,
.�{FF�47��
�I�T�W��>��E���U[�*�q�H���|�ݺ�����%x�A��X�x����ފ�h|�@�wh���&)�doڴ��ħb��OfG�H-��WY�-��5d��� ������̮%�X�i	i��@D/��|d�͘WC�: _[0EVGs�m�}O�Ǝ�����~�LR��Ie0}�`5��G.��UЅ��_A*�x�f],EFuT~Ks�o
F�}�Iμa-ȯ���^N`p�i�Л�����}o�#i�b��p__�z�zE��\�z�����I����x�Gctx��(RX���	b��x !��}�J� f����S�����E�A�%ߨ��O�l�>˪�v�ݽ�����F;��G$�҅5%&�
[���;���'3JVc��Xu�	 ����X3�d���g�I�.Vˁ'sx�]�r��������jϐxAx�T����;i�8O�s����H���]�,:=�Pכ3"��zT��>|�("�������,MP���
�J+�7�u 2� ���w�eT�W�?7�u��8��.u�Ae���\�^	��m%�B�2�p�d	�.�����,bBr{��w߲�
��W�s���x��d�"ٮp���f��G��)��R��� ޞ�Of�M�I����=����@�A^<�;�[�|��$��ƛ� ƥ#�S�ŏׯ��/�k�����U�(����ȇHÉټS��Z����c]i@OE1�}��T����i��)�s
)?M��X��D�8��x���ZT��7O_���b"J1������c�(�]��"U`����~�9�HFFmB�;��A ��U1a��/S����L�<X\�C�F�)b���fM���@S<l�Ni�m�����!X��h��fq�޴B��Y�tp\�{j'=è�!�}|�LF�:V\�64^D.���{�Ѽ�0��y��s����K�Ȁ��G���fJ�	�JQX?Yi)p���ԵY4z3��!&R �c��2m-E��DCOK-�Gr��L,�Y;V}�ފo�����W;w�K���*��{� .�^�YWӝ���BH֓�Њf�J��5����iNel��%e�DW�C�A@~��Z�fyՌ4�$�v*�x,\S�Oz\��O���D/����=J�+ᾙ��3�G�YA�G���Q���i��QES~g��[���{�"G��u[Aˁ�0ě��町�ɖ�C*8u�ߑE�_E��0cwb/Nji���I8��!�r�.�y�l�A������ w�g��*�����b� ��<�*~�[���;|��	��ݽ�2��\������O|JL`OO0�-wr�k�V��&{H3�4)aC��5��Ji9��>B4'�ZL0�}6�7R`u�#�ݴ�8�ĤEK7/����e}��J���Nk {A����ȇ��B̎��v�	nY3O��f*�R)8�_7��M;7���m�I�zPG#"R������zە���i��w9ep���n�5ꍃ�V��c��l݉��D�,:���e���`�賩2�;��������2+�V�w*�Bs�2ޒվ��7����O�~-1�:������
�!R{9]�@Z"q���TٱD*�;v?2�5����H�<�nC���a�)�Ap�߱hџ�1h��yp��|��ʇ\��"TR� $�=�$$(�y���P�B�CM��hDT�Qa&Ե_����^�)��X鈴�b�~K��B���5�a
y5b���i�[/6�����r�K�@��x��zt�O�#��^�U���� � ���(7�Z��F�;A����0v�t�S*%�΅�}�mӲ��͠aɺG�?t>�3�*�*)r�Ԁ�+�z��tR����d�;8�x�ю-</��&�5d�<�yjRPkOj2���	����F��F�ҏ�'tc�b9�^@���G�����`�7X�6O�)�K�0^�բ����6@6T@Pق�1���)B�\F�L��$>�3��
�������J �$�[��Т�L���j�l9��Q��\������<����f�?�?l-]G�����C�a��b?r|l��<l#���!����,)]8̎��)��U����0�K�J>����K&� �Kײ[�����U8Z}�V[�:O����[W�7�88�4�Z�����EV�
�-�&�g�!Fm,(�ѭ�ה)-N+٤��D$�"63M�O�.γE�\
Mj�;��Y��a�i [
�0�yoO���ty(�8�D��U��Vk�[,�Um6�m�ʐQ(���逸�c���(��炅z�k���R�NoWF�I�U�m���T�B�(r(���u<i��&c���1�<�l;)�ѹ�<mH��y�E�\���p�t�VvX�o�!�FP�X��?�� C�3�'^��x��X�&sZQ �ؼ#�������v�K���z��Z��F��%��}u�)g�q'u���bx�����kwin\���U,��1���݇��O7��Xo*o2I��8i6r�.K_i����A`B���� ؇�΢p;��O���Y�N�t�,H���F6�r��G�݃�˪�!"��h��.�BL�(�HZ�&e�@R%A������K�[��h<Gp�b���c�1�~qz���E�u�-;��i/k�_�W��۱�[t���)j���\5TKm�j:ԻD�L�����P�?���&O�!@�y�������n?��k�C$)���=[rj	�˥�Lq�X���|��Ðгe�0�'B]?@��{OQɀ��e����U����Ԙb֟-H����y�NǁW�i?y0'�<ӿ���>�~����F��)�L���}O���r�9��<U�w�at�mK�P�t�@}�ftc$�[��YL�$�pDʜ�;�(P-���Ӕ�
0GF�����y�~��x�K�K�š�6�?�$�X�A5�,p.�=�R����6�@'��<Ő�Xk��ew>J��ɴ�h�7󚴰�tF)o����[�f�p�aguȋ��u�d��kr���.`�_��ǃ���Q��t l@���xj�x���c�s���֌*�\"��_��5JYIjgY6���C�q)�H��|�'	��C�r���4��k�]c�ŀ��k�Ĉ�ng��r0�./Z�����Oh�B ��Bn��0�qij�n�. �۵��k�;��S��R%�P:SU��^jZz��ִX�)!��a�����w�aL!{��),�E��)���w�����%�+�:�u��1F.zn9�)_�x,{	�m�ы7��Ez8Z�wD��+ oUcZu=o+B�3y?��7ZzX�J�9��+�@Y��`;�X��K	�ǜ��g���ZBe{��?!��
kx6��4�ͭ�AP��P��a�M�6��n�w�5A��Cq��X�X�m'����%&�Gs��TL����{����1_�	[G�x�p�.━�1�d��b���t�{��A>�T�������Ԡۄ� /�0w.��f�R��z�ݕ�"� �s�������u�D��!"������/�y*���Y��&�"?;�f'A٦7;�Gf�J�1�яr�d�>,�v;�?yT��毀6���lo���J��AF�Fd�q�P�,a�"
,)��R�P��n	�0�n���B鞒se���ٗL�y]�X���kٹ�_�޴/�ȴ:�y�N�̆��#��I����G@
�ݛ� ?8"_�� jW�JנC \NDk�德 �0�:E֟����i�l�R&�)֗}��1����\Պcm>�g���g�K�u�2{tJ�1�N��e)@|�JJ�4en�8�F� õ����C6��7�?L��<��*��������'t�kAe�o��#��Q��|��;G��G��ML����e���!�$!�����`]��X؍�E�,S�J�hD~�;J�W��R'�/*:�q���H�b�`�&<���ð���>&�2d�\��D��	�gO�-M�Z�7�the6��rP������(�I���y�ޮ^_�h��s<:��p����Myh����T�+����v��U.��ܳ�&�)��Ｆ4�Xc��i̜�����,\sl��@d=����q�y�KĠ�'���_Ԑ�vA�Rƌ��l[q�v��Α�F�"Հ8rA��Xi۱8F�������3ot�#�Q7%���� �A$�}_k���K���	�z��k%�������8S������W18F��D`��
3n�h�8�(��\�S�	%etd�Z�����[�3�V�1ネ��!Gl4R��76�R�"ˍ�S�D<�����4��'�K//���^�>�ͺѫ�dCI	5���Xh1<0��d%s�@+C��cX��>1�y̧�'} ������i��n~�凪��Yg�1�ƺCQxw`h@:@.X?���C=9}}�m�}3�QJ�Q7��( Q��e-Yi���҂�$|��"��!�u�]�����Ϟ�J�g��~c��ޛ�-�T���znNj�X�2�Q�ա���PD��zҨ^��� �k�?@�t�WH�����D)<�d������r�i� ^Q�[K�S��^S&�IM��h����#y虱��ыdi2�3=�rL��xh`/%]A�̙s7�#�?�VD���.d;���䈢'�^����*}8�" �H�O Qzr����=�<�r��ߓ�<�\|�NQ�X"��h#(ͼ����/�B*��d� T�϶e(�>=�˂sw�,�F9�A�Zb�-2h��d��[��sω��b8�;O��X�Ǩ�����p�E��^�X�����R�F��^�q7�L_"�_�3}s7R�c6ӎ��D��T��N:�0ېd��R�S�����F���`��)!���0-yJq�Fa�J��>�;鳧1�%$���U~7��Vl�1+�)b*�KS�5�9|�ȝE$�$Q������fH��q��N��e�Ad�V�#2	7��qE�[�����5�b�C�x��P:\�m5�w�9#t�A�բ�4=�����GŸ%�N�_5��m����W��cS��#/F�����2.l��*��;)�M�t� ��`�ۉ<|���뇷d=A���O�����)�k�T`8��\��
��y0O��"zXr_0�����J�Z�x�r�u�F��$�ZY�^�.���3� Kd�/0p|�T���z�L0�_�a�2/{���6F���z��
����}�ę��I
�RڡwR�/]Hr�'ގ^y�%�������A���x(���L{���oA^Bm�g�Z��cU�>E�S�'t�>3����`�>��LBʸ��WY@LA�Znv� �� �`Z�>��<9|p.�u�d�Z}���\'lG�gXk_1�ffX�bwa�C�~��+��9��,ȇM�ɸ��z`��1ޒ�MZOioP�X����3����8�^�k[�㣡勓SHО�fɰ�� ���� S	���F��x�s�]�Sp�t�Ǖ#����z��5.+ʁݥՕq�j��K�����,IF�q�m7�nȐ۾>�27�W��{(�S۟}vC��ٍ���;��a�(���k����%�{��>8
��j�~��2��yq[1N��'��Ys^��/���oM��<��Q+����&��X	�0oB�W�7��	�u2ׇ�Do]��+�YOn�Y���8+���3��I$�|���.{'
�v�Ô	����S�1Dme���bio5?Z�FK�����
	P5L^��{D�'�E��Q���W� �3���'�8��3�
�]��X�d���ņ�Z�	��@��ӱ	����^-+�����/��F���ZF�V{/�� ИnG7X����;-_��d�����+��	���C8j��ۇj�`Y�<vЮh�qk,�a�T�3�(xO+[�z���~�Eڛ�])|
8p��S�����v໯��2��A������c3��~���ay�+^�X���o�o�oJ2�_
����Fq*"ie�:�t鯗/�lxsH��o�*�\;_�.�t��<��G�ԉ����ӊ����D���6I~�@�z�L�P�[e�A�+_�д�9cXȩ%�Y�H�٣���5�L �)J�����YTĥ�!PJ)������qo�N����mx
NmnB�j�>=.' ���]4cOJ�G��yʍ�$������M���7/5���<�f�
����%������[;|���Aܗ��=Xm���ެ�*m;T3(O�3q1)	��dm���<pN=c8 �тj7ˌ�@>i��	R���V*��]3K���?{ j���}��@p
����}���NuT�����zi����`q�X`osϗ��߷Ҡۍ}�k��Rp���k��W�Qonaj4-�m��D��0�vY�C�??4����=��T+!��T����S?���v���K{
�)
c�6�a�(mU���6D���)���4Ti��d�n	�9��DlWyI�Q���6[u��U ��
��JCx_a� 	/�����0��A�X�!��ws�eRk�z�[��}a]�^.=zy� �dg���R�l�F�4���$1D��{	B��\��6�wf:ɔ0�	���|��w��D��[��x�5g�<o�i��~@%)P�>�7���в�u-Y[�?z21[2r��Ks���������ٖ=����Og�}%��fc���JF)o���Q��XW�r���ur��bF�?@��}��t#Qg�+x^�� ��m��eg�m�Ӆ��`>�`h��0�w	��^�}�^P��O��(�ь�tr	��ZD9�6%\�"����,03>+U�M�P=�u���fh�v����e-����ʘ!��&';��r~�;�XE����>>���]�S�U5�O��<w�d?0��G@Xr���\�rN��攨!���5�D�4.v����*W�Q�7�� '��(_~��(OR�

|L�����	��޹��f���[�W�` ��V#` �V�X]�Y ��E��:� �+.�fHN�!��*��ƞ�Do�;#���K�� �������@hV;��U�B�4q�����Q�ì*3'e�3ŶA,���|Y �Z ���!�yI](�`v��)�����Grk�_�Ə��9
���l��P��QiC��ʸX
��e__7�]0��M��MًM��B�S�k�it�ǉy�wٿ\�Y�������胄�VbB!��D�h#�%I�O@С]HS���a�Ku״x�
�m�6�D�Y4z��_���8�|��H��݁&��'K���s�A�1lJ�m��{��s�'�79����+?�*׾���?ޔOv�qX��t�n��?��O���˸q�҉iXD�F�41v���ۨ#�#��� �o�Eo���39�n��%�Qˊ;��&�\�k��U�T����Fu�q��x�9��z�~\!�c'Rޛ_�WT-g�ſ�x����:Y\D�W��*v%�ENV�ש�`Kى�(_���i5D�*���pVa*��
Q8	�k�Ue�K�X��ܻ��N{[.�[<��x�buƥJV�(�4�`B^-�c� c�m�/���5
F'o�{Ke�����mt�5���ZwSw�x���!�����F\Z2SR�| ���i1�&��+�\%L��ov�IR�9Ò鴀��X�>����/D�֨�3F�B���V%�k3�"H�(>#3Ǩ�~Y�e�d���C�v��a�2'�c���*E
��Nr��֔!S�2K��KR���+~'�~;y�a��g����M�,#�t�Ɲ�����HH���k_1<��) ��=uL�̙_V��s��HǨ��`֭�jWtb3��?��|Ѝ�I��yk�^��Yݲ\8��Uʗ6fډ�@��G��:�g�B�nb���v��K��� Ɨ�WF\�b�\��I���9�\� �JPMe�b.�W����������5˳�K�5ʜ�L��8�Ɉ0��H�Zr!�"��5u�!������>$��ݓ��Q+|�(�k�cfQ\���<���Cd��2�
�?�n�I�(Ȣ�ѥ�"������x�0�A���`I�`��;i��A[�{a�Sx0�,��E�s3p�(�°2[�b0Y�=C.C�HM�������X�-�5�#!�4B�v-��<	����p�B�`�S�Z�'k�����<EH��Ƹ��J�C�:��ߛ�G�<���V1���e��;��Y��B�f�{�e�x�P��ȺU�+v�t�����8Pr�y'���a���@�g��m>3ƲW4Bm�U�Z��r���,6����r�H��6��܉�l�����K棢ߵ{_��`V?6R@�?�l἞�B��udԊ^_�`ۚ^����.�ŏYN�͢����ڠ��<-���t[z��p
��xTu+7����s��4>�Ӻl��hx�!��h�Ye]w#�y����~�4\`D_@J����F �44g:�d�p*��g�H���%n	oe`��;�M6E��9��R�T%��X�x�9�3��A�,Kӹ��Kf^��*�@X�z��"&�7"wS⍐��ኁ'X#�G���l��0/���V��!�b�M����f�6��ɻ��is�o�_��UQWcF�v&���3d���-ʹ�?;L�y���o��A����/g�w����8�XR�?F��a�D��q=~�:�k��'����	���"���4��9XF̾�q�_���c�fA����y��ւ>4�(��������w��Ec�*?;���##zY�nlŌ����ʇh�vW��`�WQ��t.���lh�OvV�H��\���	�U[!�Wzs������Ø3_!�[a�ӥ�Z��n]\��zP�Ėb�;�|���Ψ��r� Y�>�߳�C���K$��h�q.Ε#L�a�8uj���-�	>� ���z��SR����,k��ϹYW����g(������G��q�M{�HC�'�C���Idx9��-�k�����B��h��K�����\H��p��F A�T/�.�Ê�:��BVX�U�Pn{�n��R�,�ӎ����3��~���8A�4��:s�@+����K�(C�G�c`K�����;�'�1�
�,�5O�挧x�P-W�m��iV"�����k�*��5Tx�j��FVl*}��(d��@:&h���cUGg̡d��|^����)�Xzz�k+]���5n�:EB	��T4���3��\!���Z����z�(h��l=*WUi� �yt���sj<�gFwf����q嚷�o�� �.Q�)Q#��z#�h2?���N�0���.o����P1\d
.���v��~?��o�/��#���#�I���������G���N!��5�Q�D�-M��KTX��"� L,�g`�@j�&_��M��s4��s_�]r*�\�K�Zd�Yc�d�J�Wے�L�x��
���q7x����[T@A���lF�U?"1/�YU�A�ݧ|p�-����=6m*C"RWH�0�YA�)�U�W���&1^�/�U0�Kg?I�av�p�8�k���.7�gY@��1"��箚9�j$����?�S.��	�-���h A�8��=$|^ގ^�'!�qʚ�(rc���Ǔ=��q3�]�v��NJ�eS����
����1r)�������=�G����zm�2-;��+�xw��ⴸ�UF�i�-�$z�HS�F���	zfB��٨�rV�fD}q���B�ﱶt�\Q�e���P�f�465mX�`�Y�lO�
;:N����d_�<x1�����.�֙T�C���$�}�ko�[�;�`����O�9� �NF8�'��9Е�k����/�fV-�3��W�6><�d&�%���CZ��[�yTi��M�8~� �'Yɧ-#����KF��1��`
��"��J�>��=�(���E�9~�����}&�Vس%w�)^["-ĕ'w؜'X�����!���1VB^ {���:>Z���4����B��0A	धZ�!
�]A�۵�� Ĉ@�����V�*�![�CfkGN�uA��?"n����}���}XΘ�g.���ә\>B���/$��m��ג&3�>�Y���4d�t<)����j����L����x{8����2��gי�eu�E��
�_[�Y�	f8��'��T�u�����#�1��>Ԣ���!��T@�}v3	�G�Mt���Ė��e�g�e�� �;C2+(E�Λ���N��R�Qaw�~���O���"IY���lM�k�ȩ�-I��ľꑦ�Ḣ&��F>��G���"�Q)_�f�-
 {�S�$N�(F���dY_t8s���3^+Ȣ���q8 ���TG��-�U��b2\?�zf�ěm���k�a@���������$zN�p*�P����GP��~ᥓ�p����}ĕu�@g�G��~��x�Ԅ$Di���w��TŇ�
'�T�t��P:�6ߔ�w��DA��l ��F�X�E�_r'���9̶{�����Hj�ĺD`՘�����%���0�R������EO�N
�U��X���}��NL*�SӳoD��'ð?�$��4t�'E͢��D7��RGX�ₐB�f�?�O3c5�����Ǒ��&�h:� ]�8���>v����j!x�\���畨V�'��ؐM��أ�X̑N(��o�.щ�B~K�����h�וTu-6��Z^k��w���"ד�08`e{�a͓)��`=��[.H�s��?F�<��Y=�kU�=}�S1<�9� �=�F�_��.�Oy��F/����x=����?�0�[H�`yL��9 �z��ӳ�������!P[ZS��[���fs>�=��+_�P -�R�3��z�N]�=r��T_��)��\%�A��u��<���율�!�����"�mVB��1�$(���e�7�N�bz�� f�l)��ZCZ(�h��6ħJ���8P��ũ�z�"����H>�I{΍YedǕ��
���w�<o~�1��
�������Y9{�)���Њ�Qy@��}�LL���t;I1Ĩ+�,>U	x�'G1N�:�C����a�M�����Q�x�� y�5�,�P~&�(t
�>`p=&�x�����:ϜL`�!Ӄ&F���#g$��{�V��H�#(�[�H^2���S��1�<z�4\�������2�oҳ��Jb7�4OmF��Rzii���;Y��!�6O
�Yw����Y��k����u�plL�͙�`��r�� ������k�^��Bͳ�8M�g �2oT�Z��n�#�gns����,أ�.��5�� dԯ��5��43WL���e�:��Wz��w1[n�KW (n|4��gu��aN��z�5CT$GX�C����n��:Bk:j�=������՛�(֜�.G���/�,�Sp�X$I��q{q�[��!e=������6)l搭���5��_����"�]%�����<�}��#�Z��p��9���mã��T����`�x��IIn~r�	�A�>��7��i?�ЬlA�X�tV��MP�B�t��7����60@|GG��7F�XS�^u��w����a�J��]z}�l�
�F`��$�.�bA�9t�jҸ�#�u��H���SW&��Yg3;ip/��k8o�k�::�ѐ��6�rM���k|~v�G{!Ő�����S��L��:S"��<���,#_	�*�B��u��#-�$o�A��A��Q&�O��%MYDO1�g�i/�+Z^n�;�Eq�=���v��,�����uB�B$��?���	�g/x�x;b[�ۙa�=�zk�?�Y�'M�%˱�����=hF�J��>1-�!�*���G��Qy����C&��>�*�p���sh����MQk��_X��i�lC|	����'�"P�V�FR�r@p�� D����A(��ۑ��=�l��2*�t�|a�!��|�_.GC~@�(E-��(�K���M���������3/\�����T���'��f]=+E��U̇�_�a;��ځ螔t$�n�[�(���,�ZJP��v�b_h�����wC��q�t���!��hiL�3G���ե�!(�ETU�,�j���	/��dI���&Z}^dH"�.��t[�D�ӹ݀��x�)�9)<jʷi0����{����qyl�e�s������Wz�-]xJ����ޓ��Vӗ�m,��@��
(P
�[�D�9�1J5��T,�f��gؤ��r�˻� ���YǛ�ad|�'��NK�r�����([;��G�T��>�@\Ť��;�]�Љ��;���x���T9Y�0���~r-^���&��(�+k7hoAA��a:�i߸�.�f)^�,�p(����Ux1�p�1�B��s(��l��+�:������H�B2;�j�f�!�5[��A���0*mX���u��������9�E���0p7�.��3��)�-�;/m�e�į���,d �O�:J)X
Lm6Xb�'��n�����I3R l)mJ�s>	oe;��<�IU���M6�2���kZyH��Q���J�GXL�2��j1�e�WӎTp�]�N�a�4�=��ع��j���W�d��Qb�8'����6�&�����4Ϙ�_U�o�j��^�d*(��۬������w���kޯ�|^(���}.�8����������WbJ��p�P��E�M��=����kO�
�4������Q,��$�cd!����X��'1�md�.l{W�c�k��I��Q��۾#ӌ[��2Q,�,�m�7NV�p];�_�Buc�%�ަ���m'�b��]��?�ϟ�m�aR-+�c�٢����l�T*@6J�x���p>:�TaJ�`\BƤ�	�������p��
����: (w#O2~TF@o|Y�w��v�t�TS����OG�%�A���)�Yx�g_�M�����H4&�1�]�����y}ϱ���� y�-�����Y�ͅ'ul��S����֬��!7�u2L��?���D�:4�	% '��R�!n��mT��^z������qcw��@$`�$�Ѝ��o���%F��2DTc��D�}�#u.,�遏Η{H*���`p��Q��s�qzm�1p��ӷ���kU=��o=�I�I�9��o���VPmM?Κ@W�s���XH�ZX��B�}Z�����k�`M��
��բ�R�*�����C���8р��bw9D��<%ݫ+��9����`�&���$����RX,͜lP<Q�j��i�T�z��~�Q=ˊL�ZE���{��~G
����"F��S\G!����­�ì�z�U�-��C*_FB.4
X�,��m�C���{l��B�3ր����-㕖<����(�xb�vh�9����O@m	]w:{�s�����u&eZIZB.�6,!�؃�cܸb������W�N�h�w�&����P�����v4���I���O��5�g"���$�z:�m�1���D�Izm�� �Ve���=S�_S'02)]�v���$�τ�ԢM����HB��D��e�aɸE:(i�"�r	K1.N>'צQM�HP�v�>8!Ό�-����UD�.K���z�/�i�$����(�4�+�(���}�3�ck��Y�Y�8o��rآ;[R�U��O[PۑI��482���兠Кd�fc��@i�M�B?w
~h���(��d)�M]�oQ9?)�A�(�whyPp��{��H�M�����o����2]�����I0b�Im����R,�|5G�-�H�.�J���=��̀��`�-�d?����ɑ�IElp�d�GQo�+fȇ�[w1 zݻk!~��)�%oO��u�r�I�=i��,o�M���Tʬ���3B׷TL����]�=��Q��g�Ƭ6�53I\5�il��'lk�8�G�>��ߊ�KF��2�ƀ�=A!����.z�Ґr3�I����J�6MJ�1](�a�pQ���(>'����]�������訆�W�raW�ͯ���E���{'��{���7��!�&{���=]�l��B��p|Sx'�S2v��H"�|r!$�������[{�|gk���F�4��d�+�
JK/q�5;J���V�,�SY\�����W(�Zfދ�b"u/hG�m�^L<`���y�ح�b6T=đ�����tp�cH�з��,p'������a��J]�������� �3��˰<P˽Q�%K�4m!���4`�����&����*�_�փ�&��⇯���d�h�w� �Et���i�����`��ޏᲚ��~#�7%��)[(.{y{�9�����4��Hs�r�V�����G�����u66���l;���sC'Xz+�n]���e\���4I��Z3&��d����<H�#u����*�դ-��j�'.�����Hhl6@lh�ω���ٖ�Ӭ�|��؟)!���j�|�;�����Rc>�[����4��mL�Q��A�\��N���:
�޸s�$�Ak-Y�236F����tշ�;n��=��H���&ث��G���K��c�!���咶��n��v�s�&&;��t����2��k�`4�\lw���T�V��)Ƶm�9���*�6��d�f�M]&}��\n�ո��"ҹ 8��?�$|���� ST)Q��%N�SSsa��X�bj����9��#Uu]��7v:P�Vp���2�����D��Z#��)�V��� ����3�ҵ�b�(p���X-Af�U~�eg�B������rT�g+0�O�{u��tˌ�:�q-980�v�G���U�0S	�#����>���}M-��b.��{�J��{�S�DӦ�f����T�ek���A��{��(��\#H|�l��*�X8��N3�F�����?Rwv��Y���j���IG��-t[��Dz["*��������b��b���VFj��>p��8�_��{��u\�9s��� JE��ov��g10bd���_�әJ+�C��D�l��W��uN�	��Tp����Q��!�T�r��sx �0f}�۱������UϮ=iq]�/§�8G̢[(L���K�G�����3��k�/POt%�[�eo�"P�'�M�C�C_��=�
Hf'D?	���u���K�7�JV�s9Q�%I�����Ck�y"L�(ӧ�&m]�Q��i��S�m�E��"�L��v<�H듛�U�ٿ���Z���HJ���.֑]=U��@ =Lc5@4�+���:3���8���.�M�u�d��k��j��7�R������H.D2�|�!�|Ұt�gr����xW)�rܒ;�$:���j�����=��P�+�����~����V�s��^@�H�gy*l����^��!�F�1}(:\��{lz?�D�'&��#����,�	�A����v�v���,��	�w���hl��[��1�qh;��O[u�j��8�e� �^����[�h����XI��Y��FEױ���2��0]@~�hT�
�T��?���ՃX�J�
���h���R�y���򾾠�~�A�1쏪E��rv��X�8fY̐n�&${��ZZ��Ƙ����꡻��j�x�'�a ����9;�!�s}�4Ζ�V�H��9�R��6��c_�BTŸ�������!��f
L����>��6��#��Uݽ�GIqJ�&�	��������4�5f��.bl�jk �~�4{�n/���%�V��?���T�w��!n����%(,=�V{���1}e���؉=Vn�B,e����h��`�KV<p���WL-~�t���2W��*��I;"r�ʸ��Y`��4��� ��G�MkH�0K���w��<hb��nJ�n�4N�°R�]�\
���-]1�K��v��;�3y�~��ɎXθ�ePJ�^힔���FeئQz�B:�d���
������a�O�bZׁЏ1���ch��x���G�FN�g������x+�f�U{�@�Mb�[�Ƴ�7
dm�(ƭqM��D��I1@2�9�L����b��>�V�=9�1.M:�T���kߛ2�1@��"
�f�!���y�_f{,T�0��#A|t��i�����M݊�j�T:�,�_�;+��e�ҽԭXڙU��j4m��y���J�+yH۠n.�^�!�M�I4� d
&�V�����'����f�8�؄���CS,9�>O"�@^���HZ��%�eV[��� w�bs���!
��]թjُ�#�5���$���=��J`�G5�LG��)JyP^�=��T���.�����7vC8q�$l�![	ʅ�&0���7O�β�|HM�Ǿ�z��]�^�!/��m��"�D���*KJ˓V���x8V�P��z�N���rh� �+g|�ēj�N9��јL�u�H�%���]��� ��dEC'Pt�t�K�
!� ��F��uM��A���3�g�"!1���ɗ3�y�s��:.E=��Ic��#�f/�A3=��?�Y�}�v`�Дq��Y�aG�0p��>C��������;�������tLf������iU,�w�t{�˹8� g"��p{{'��i��b,Ie�_i���] �$�.v^�/����n��<@�c�m|�x�Z0v�_�.�����[M��uur!�?���!I]�BS=p�xꗏ��
��=f<���M2|U�n�.QG^d�ނFW꿅�ƾܘ���s������`J��>6����1�}��F1��셕xF��1H!�������1bޢ-�p��ߗ�2%E��a���E��p�>)�R���v8�q��k��!���2v��+�V`_�4Ɂ"E�� ����m.��Vy�]�f.g�]j Cl�����&)�:/��r��;G��vl���[�_�	>��DJTa��M����o�
z�L_(���)ЭS�����p�Ty�����~�\5���n����2�7z�:���x:��i�C8�bzI{���ӆ[h�(`J�ہ�AR��t�Dxߘ�[�ϿrB��D�Sw���Y6��E�p��%&�
j�lŬ���2@u�0�)I�P�2)ޢ#�kJ3�E�)/r��6$´�E�8��
#����NJ:EY.�Ǧ���{�Z�� T�(������c}�ê�P�
��/�;smxW;�|�C5�w�U�\��wz�x��!ǜ���e֧P�Ғ'�H�d�5���x��Vÿ�lZ�H���f�Ԇ�����������a"�"������tY0�#�l�ף�,\��%n��ϫ6���l�kvW�W��Ci�SsO�1��J��E"����6�����H2��"�l�7�c���Ms;c-�Bb$����GG����_1.��LA�)s.�fQ|;��	�~�P�xO.��4B�X��tO�be
��aT�\ X{�������M�@��ve=���f%��:�b�Ɔu���Dl�AOU]h9-��h�;����ԗ4��L���3��[.��ݼ�h����D9`� �4)T��b�}���?J~)u �'�2_������/9���h���$,8N����_�<}_�>�K�&�$��F�q��i�ppN���`�|�	1yl�<��ZkeF��Xp}4�+kp���JN�^�[ʣ���<r�/�H�4d�O����6`�(ɒ��
>Z���C2t#T%�Ǧ��ԗ�$���Y}��oBt���DO�r3 Хy��D��.K��
]��G1s�R�m�ذ	��������}A�$ꚠ�7��}����6ڡ��x������!L��E���(� /^�v&t��}B�q 匂����x�spf��c����oeB�nF��[(~{fn�2�/�y�y� qb�-�����R娨\|�R�EwI����5+�C�Pk�;
]�⮸M��u�H4�67��6��*�����Y�<i��G/��P���]��N�?�SB^1�(�Wt%�x�|�����s��0�Ғ��u;��Rb�4ؔȘ3�Į�}�������c7���r|x��1líG\��(+�S�cs����<�0J��5�%r���ZJ(�?S�m�g�Y���y��ð9��{̲.A,�m�t�U7�_�/�(F�1���շ�r7���+aO�*�ȧ�{?gp����z���Q�N�� {ذ�CW�`곿T��-k::e��Z�H��^L9���_L�}����u���x�t�P�tNm����;p�B�y������S����w���3�	��ڿ�����po$�LNg�oI�/'��?-M�2��^H�k_V�a�І(��~+�y�]�1��q.So������X�����?��i�U��ba���$nՀ���M�v���ي��� �^�7���]�\ 4�^۝��3X�
�>�;:��@���O�v��pZ7�M�esTOE��smN�Zz��Q������f����9�"��MZJNf����^��/3l!�چO�fI�yo����������Ź�W~n�_o�&��1$�i�I���:f4}��"���8��<4Q�w$bhn�B|E���
o�À���ĉ4��"�����fe�cy�߉?̡H�<�{F�$�]Gʧ�r6J��Sj����<����%��C�}��K?u$�מ��&���/4���\�']�n�=�W�q��L�Y�W��<��m���|��O�wA�'D�-S��8ѻ�u���*k*|��ͧ#ڏ�s����v�g�����AK\'�6���`#O�he��� 
#�|V1f_�]?Gw��F��Ϥ.'�n���rQ������*�����_�/���ya�lx=����e[M�*�w\Z����Dn�s�N����W.f���@I+hVI��b�e��\:��]�����z�UZ����O���-�g���%�������}m"�ÊpV��$νl��7ڶ[Ac��uJ��$�y�^w�|b ��N8�t�:X�I6q?���\c��,���oK������Q�|�N�PV~��� �%����>�&I������KYs�]c<?���n��8/RH~02�-�)�o�$��������^��� G����q��؋P�g<I��,�Uu�h���hg<&w4R$���Z]��)NJ,TnGo�E��?��}��hgy,�"�]`�ƫ�	K7�^���Rw��V��� ;���J��XeR@�+�!)����ge�z䇜���F��b>��޿9�y�)��]���D����];�b�b�$⌏���,󶝊۶?7s6������F?�q�=˦Ũ�bH��n+��Oֺ��棂�3��]<R*��!e��"&{Nͤ��\�Ƅ�, �g�c�r�K��u�ZN��0����9����se�A�~b�&�$���6�}[/�U����T4�� U�/���!q)�Fv��<x��>%�(y�*	�є�|jM�zMO`@�X�
.Hh12l�0�Cd�J}�q�K7�!s0?�=kNK]���/�\��dZ)a��m����"/�kk<QB����܀��� Ґ�R�x&��43��)S���j����H��R��M�^M��>?y�L�Z��ZKu��f>Xy��� �%�W������{Ϩ ���K��n�������n�pwu諃�.2
�Z:��[�5_���m�_����[��f�z7�k��
�k�L�0���ģbO��f�SU�0FX�*s �������<�E���B�i�,�D�wR
[�NO�~~�U���[���̒���<uy�&J��w	��0���g�)Tx��7�>�������!i��%�1���x���G�h.|B�;�ưx�c����3�ɮ�	���;yj@�IŅ��h��dkv��Գ��� ?Їle�	�X��_y�)�\�c}����3�w&���g�4�e��-��
T�Lk�(���ҥ����n+�C�PD;��\2.�WA���Ϛd	}�G���i�b�l��'&�yN��L8��=@�p8�P0Ό��f9D4�O�����hq��3��P�BG��f��@)EK��i�G0i
C��icn ��E0��n칫������}�@Zl���QO�YV��ޢ
�����X`�����~��*�X�#V~�	�K���e'��5�[�Q)�u����� CgANE(��$�C���2A^��Z�u��}��	@�8뢳ez�`�`��B�G��+��ڃ���_��c���������CfDX����Z�����G���P�<��pu%vÈ(s��H���Q��;}��AF��mi����m�n�p���ג=����n�
��U1� �iW��T��m���_F>�B>�8]�,:_~��jO ���`��|}V���X��%��a � �5p���f���]*?��r��"p7riY�fH%�r�1�����bހ#K�§j�Y��ȆD�~ 0t������P/)4��������gʿ!��ݩ�c7�"��wR��5^��M^�㛟$!k�L�X��xJ���%�wԿ"�G���DD�k�W�0j�h�v{�du��`�c%�%'-��_��K�u�I�Kڴ*k���*�{�%����	:�Ko�	eqG�fſ+����佶����}�[<H`�w�z��ڿ�^��G]6��ˀ��/(�{LF�r��3Z���сd�	�)���`�͟F�|}�����Q4B�3UI�~?ÿT���7֯�ըY�,��	��f;��N[R�89� ���֗�v��Y�����
�4Q�p�8� v�)�"������U�?1�{;��)Uè=�^<н��7�✪�D�SՂ�gE�{-�	��@�d6�.�������D��B&d�F�jq�F�(f���2�N{�k����E�a����"j?�lG 9��9Yʅs%�k��8�����E��^j�E�`��@_�x�K��e5����E�M��Hx�T{x����@�����q|�>��JR��nΈ�N�@��]�b�cG-����/|�Aփ����vЏd��	�D��_v��*]؆�q�I���Y9&v�e�\Ő���թ�ԺhD�T���)Q�1�3>�)L�*՛�\#�_���\qzxO������#��V�Mm�P�x]me�&6mqѹ5<T��%u�ڟ�7 ����85�`:2ꢹ_Azj|]���Cxb	�lbe�鹜O[�\�ҵ�9g�q�2����=��Ѽ,��׾�SqM<�N��q׃���;��^;��ޓT'�W>a�x5���T�2%BQ_3EZ1-S�}�߂c���U�4�I���6�s�%+*�g�������0���~F�0�A�N["5<���U��ׅ�Y.�����5������S�㕂�R�Q$�xҐR���+�b����o��n�R`�1�����v�4�FJG��_�Qe�禮�+݃�C�Y<3�ʠ�A\��$�}�l���/7ܣ�4��}��o�w5���ۼ7'D��L(�:�x��7��8��M��N�@Ⱦ,զ ��0vި})N��B����1
�k)߫M���Y��	�7���J�S �(а��@r�?�pN'�Ё5oC�#hH���L�G;,�1��g�����DG�i��'#l�\��g�nZ�A{V�3=�����<����������ϖD��	�����"��&��$$1ۓ��� Kv�LUAl`pk�lƧ��o�s�8!���tif�|!�ӕf�5�{���
rM��P۶��������B�)��d�Z,�1�?��z��1���+�ϺyɣwW�˭��C���[DƟ4��!��k>S;mP"lG���{��������ᗟͷ�c"\�I[�wU�AFK�Q�xK{���N��z�;C.�Y�0,�z��>�6GF�e��4y���#R���u�Q>��=�*P^زW&��.ܯsj�u"�������뉶qiB9�g������E������M�0>BK�wSV�P%��D}��?��.8��E��y�NB�9p���7�m��O
�p�I!����V�I�xx�h�<��C���k�$I��m�����(��^m��0-������u1ѳn4�/Q�!��iL�ʣ���Xb��.J��=�<����|�#�!2�p����*�-�$�ڰ�]2]e���������;�3��x�c��]��ol\.�AF�O�	�`9d�n���?�V��=t���P"v��q؆�m��R�e�(�&�c?Teq���M�Y �f�9��A8��8�u�.���<�G��@^ E}
]	q.�o@�acu4�!�$��U7��.�'$L	��v�{(�Rq���Tcב���e7ܘK��h�d
[C\��Sx'jRq�4�R�kO�I�!�����i>I���}��}�H��q��d�4X0� �Pd30j�E-�/S�(Ri԰ea2�>��V߲P9��B�c>�u�!W.�OKh��e���>Ja	���0��؃�l����8�H��U��H⏾Zé�}�Gм��dΙO�|��8.1!QΨL��o��wd����5o,$S�~C�uPe����k<4�	y�cM�ț�WwvN�_�F�m�î�l��x�}8�XgG�&&G����q&��w\��X����c�	��sd	7��I*�G�B�7L@:��F��[tI��m|��7N��;�D"�rۘ8���J��1,\�.��&�X��;h��K�^V�۶��`�L���C ���v���ۑ��i�dWB9S�"/9�'j��	zPu#J��[Nw�0��&p��b�l�;1���7&�w�la�� Q��wo[�[�]��f��#���^)�
#�S��acώ}U��+��"�V���x`�o���D���1��b����bFe���k��s"�2�d�F�ɾoQ���e��faA�\4)0f��� �>-��ÊK��3zlK_7���:ѵk�Q8�zh���m�M&r&̦�����L~�w@�k	/�����>��m
G��Zw�"��(m��?p���+�϶���!����=42��d�s��@��:X���Um
[�u5�?T�����$&� %�9~�jԮ��W>����](|t'1i�2�=UM�Uq-��D���}�8e�K/�ߑ�X�2NaG��ڀ0�q�j/��w�S�c��,p�X��41�S:w1�m������cy]kh��U6ގ��t�A����j��lV�e��0�(�䌞ݔ��ˠ��`T�X>��ʡt�r�6a3��K�SY�?�M��7�D�����[)���yv�I���U�ۼ6nKW��R���y���G�˓����De3���#��O2�6�t�j~���=����v&t��`5h�H�a�vu���d��L=�An�Mi8Dz�h(W��K'�w��&�(� �ҧ�����Ej �X#tI#r�X����rۣ�@�Lv����L��ɶ����_�6��֣gM�=�s���%��g���	�;�7�Єw|��*���b�����O�7��g�΢�E�E9�Ls���d!Q`ǼmӁ�7����pH�G��aT�S��y f���uQWt����`��^|�K
S2D�H�J��ַ���;M���䨏kQ��Εd�	8��H��ݏ�\>}`�EBʋ���f�k ���sB��?�؇�݅��>���IQ�W)�0��[��ky��� /Gq�t���uW8���q!�f����(X����?�R>�Xr'W��R���w��&ƖO��І�%�ht����F�����j���8ϳ}W�a�X�<�)WY�,+×xT��1���^�r(�!e�1fBQ��y�ڔ��s��,iV�..6�)r��i}x(j1��
��U�Q/6	ȳ�[��Q�7� �N�:��3�O��%w+d�A��.�#[Fƻ�[������*�CA��:�ڊP(�C��gӯ}�n$��L3V_?���g����161)�hB/�-��1&�y��.�m��3�m��c,p��Y�����������;䷌Gԕ��O�e��}�3�����C>���zW�g.�z�$d�ߜ���|��K�YV,���\����;�K��o�� Z��y� %�̯�d�ځ��g�gT ť�y�J����!����#�G��he�@��[p *pw�uP`}�y�ua;q0�6$�������j����)X��l��D4u�^����5�ɸcG���i�@�3R�q�,�yfYɔ����_�w��MJ�;��7I��_����Au
7ŗ���U��9al�F̹"S�-y���l���H����!�{�V%i�*w^w,w���ur%��U>��}cr˼Ij��;�|�g^�+��|t�����dc�:Y����9��ΕI�'XS6�_�e�;��}�7��i��� ������B��ƻ��$o'�`t��M}8o7�J�)bm�� �m�T7\%�Ee���b��8�	-��H��sBA��S���ď��Y=�jxd�7�w�HK[�Df�T6�	[#b��eх��hk������J�Ճ`.�խ�QB`8B&��N�(n` �p!��T��@�,������E��B�eT]0�V�FΥ�![v/��b$\�B����*��f���;,��s��� �i1��Q���N���P��f~ToW�u7�~Z�Q�j"�1��pgM`�b��{��t?z:n<$�U�%�n�X�-��C��!vgY�
q��F�Kڼ���j���e�c]�ލG|<��$'0�f�>s��ǲ�`XO���y�����9ǫ�OkxA�u�U��a6�
�X�����}E���ɘ�pYK�b��[����Q�[jL�hq��ʱw���[Z�?l��Ǫq�I��P��pv�/M���؛�.�76�m%;��Zu5�@�����3vI��Z��Y��ڕ�]��na�|໅TU��tB�Ƅ���z������*�!��+6ւ���iۻSl��jا܌�AuՄΏF�]�N�p��ût��٬mOt��,7jd��QJ��b��A�J��E��=���R��@j�g�7�6z޽u��Ȩ^��i��5����/A�_�����JW���Z�],p���Qv��g�=����{\�p��^���JԵ���6�AT��8�����j�s��0в~�|K������VNȇ?�K���M���j���`�z��������r}�*�?b[�ॐʈ�Z:9~3�5���n�w#��<��� ��2�7� ױP^��eֵXB���gʌ�\GwK��y�~������iA�^�&���
�Pp�{��~�Gv�M?��R��#N-@���)!��%�@.�&g������r���+p��^r���H�x� %�<X�q�.;����)Z,����#x���N&�a=}���Ϗ�T ��sq�Bm�¯�X��ЇJ<w�B~���4I���x��\�D?I�esF��x3N�LX� ��&:�Q�Ҝg�4'�d�FM��%F!�sy܇���̚�d��ۅf��[gvWN�ߥ,ZԊ��"������������In�ՁN�]Y����zkd��g(��Q��2e���,O ��C���Xu3�@X�Z��)�<�K�'��*���:d*���`��\�n~H�nt #0��=-b��í��%Z&�	��Z�}��#)�Uۤ���B<V�i��7&hͅͲO0� `v·DՕTՅ���7�)re�qo��cp�+���3N\�0dϻ���6S]�s�V�G�#f�������?Pb@�`��>R�!���Ǝ�!
p
��	��76o��Gf�0#�>�Q;X�~.�QZX��_;��lp|0�[�e�T��o���2�- �K}� 
��_�G+m�Q��~�&&Ǳ�d���#%fG���Q�(&�b��  h���x_j���_2>�.t٥��EH\��xK8|t�Y3׏lK��S_�z�	��~]� )�x ƈX`��|]�Ĝ���^a*�[-5��=���y��V��Go;�� �].bt�K;���0�X���+��a��)�K7$	6i1:]��w1���}/<���s���Xy�|.�������qVz�g�Caݿ��S�$e����M��5����7����%$�7h�;#n(t��$h�{H��\�,��^೒���,����S����� > ��a��~��΋���-����R�ݲ<Z�Q1lGl�̋��H�V�QW�ՠe.p{̥9"���UIM�e�j�����#�S�~�k$�H��a�g���[t*S��Ȼ�н,r��xS�6������Z��ˈJ�w�dO<�(���{]�L�ӎ�4~��o��WJ�_�|��N��Y�gn�r�
-pPĖq�t{ˮU�@?d	2�0����-r��{n1M|��I���^y`�6F�R�UZ��_J�RK��:��%���G�\H��O�m�Y�|�����S��?�P1�^F�6&wf�>�b
<�PV\����#n0�R$V�� ��b��Z*�W/�8h���S�$���Xr�i�߬���ʦe����!�f|��M��&�!��/K�����6Y0g4�l��.8
�{��ᰪ�m���m5��r��E��/��c��𣫲ح�I'���t>:���_��@�Sj����y�S�1�|d����.����_��t&�
�~�G�x���z�2��e���G�8�VPO�+����U$i˚�4�sF}Wv�F

�����,�kj||�@ZOE��:jQz��(=�����-�	��t�?�8>��9�{�(V��8<Y<]�Lrh�RQ���Iν��]�C�z`QOc��m��aj��H3���X�̧�/F� IKW���6�vRV����9=X����������
D�����9��#�/���1��ێ��V(xXL�+���]��)���0�sdh=o�x�]FH�S9��c�!���ŉ�ڻ�`z��%�ڬ��u�,k��X�[�^	�Da�v��}���
��GYe�v���U������)�!f�U>�&�V%g��%�v�)h<��)�%��.�� �����eI�W{�Y�����Ɔ'��鹉;���դva�?>��:�?cI�+Kɵ. ���} af�]w'�7�I}6�e�3��V*ә\P��'9�°�, fL��n�(��y��LnR��5�W����q��z܏���k��V� 7p��2�b���!��Rm���{�i�������# ��@���=����>��]�L�8/��Gg���0^�/����7�f�t��B6�̉	g`��&\���t[�M1�j|H7�uФ��p�6����6T�f�J�?_
p��^�A7�A�}Χ��{,T�~l�ˮHސ���+_0)�CC(���\�#�HS�����E���p+X��$�\H2ԉ�A�1W	��G�J�y�#�͕*OᮦG%�B���}:�}�~;HZ�#��ϻ���\�<��h��2�t�[kJ�FDkw������� 	�iQ;$��?�;CY�}D6�&M��������� ���D�'�O�~��!��%Q�R�A�7GC� u�s࿞nmOh����� Q��&f��`A;����W����P�,7��G]�f�BT����EZAt�Se�A��K�ei��9m(-V�2[#�Y�Cʢ��~G�D�~��1`Cu�x�����6mJB �$:� �d�J����$�Rlm
2����98K1SG'w��#��*\�q��m�47�Nøbԏ�Y8�B~XH�.��e�d �v����fUY��'�gu�_7�6#6P��6D8hd�"��s؀_Z�p�e3GB����I�e�թrjօ���Є_%+:,7D}@X�'��=2�DS_�S�R��P�V�0��Wv��WT�sշ�A�M�^w�a��+V_vL�n��T5g�/����KIb!��p�M�6�u�7;*��4�'�֥��ز��z��̅:1��H��g8��'�R=,`cdb�G�v�P2��H��w�dH
:܊>ψ��:[\����>��QfZt�~����5�ew7�>�Fs� w5�fL.'78�T_�Ǵx��`����#��T�2T%���Өt�x6y���ٱ=I}� �s��D?ֵ؋��� .%Yv�o�r��	���C�qz�tW�2��s֋c�����eq�c��`ϸl�0��٦6�E���&dE��`Zi��C�ԇ�p�z=���� vơ��O�7˕E��[�AL��a<���"N$x;���u��Yс��t�����SO�n�F�����F ��<h�@��lq�q8��B�PY�T�e䏗�K�&;R^�Z7��S�e݊�;,H�������PƦR������;�>N�ǟ��7s9'�E���C�[��h���--�q�Y�ڭ�Ne�"rv���`����~�d�݄��zX��t{�C�2�Ј�e����9�E(�g?�%���\SGָx��Ņ�5��Q�s-�B�����a��w�Ǣ[a2um�`�>�rq)�z�4��^G��+>7�>��'��V+!�%`��F*�7C2�q'�Y�H��.pq��ݣ�!?ѐ '[��on%�"��є�ȃ���.���E��2��2�/��Eo���	�1�J������l(V>�[����ZB"c�p�{���6(<�jqO�,��C�m*�p����5�uF
R|T�T��W�:��	97dH��G���Y.#�*�f_��'��?�Y�_��ҴpYC\&�* ѳ�\�:�~# �=մ$4�Y�\��>D����v�[��<�6E/�f�>��هR�ˁ\��J��I�PP�o0�,c�����"�Y�=؂W$��jJ�Q��e��uv���6i~o8P��Ʋ�Ǖ������٬Y�+ܪ|A���u����	�)�c��-�ok�xW'&��v�F;��˴ʕ�4��0W��ה��z�ǊPr�g�m��K��vO&g�!��$ɹ�6%c�����F�h[��@z土?0�����MRV����GN�#� ��ث�U�v����E�k���҆
���p�4ٙ�����%���Ƭ����Դ��r�<��ԬoRY}������ի����Im�d�"Z3���`U_�W'�ռ-O�^��XЌ�jX��0C�7��L����>Z��ЉD�NN�:~�먏x��'T��\���t��w+"l14�>���V.zq� $���@���.�4�M/��k<�B~K�
a�Kx��"��mjI{�cѬ���v��xo�<��ۡ��DUح��0�$����Ĥ -ׁTm�z�3�����h��G��tA�/�
��F��A�n߸����転l���I�MV�JD����s�Q�S�}Ǻ�����mX%�"	3��Yuy"�#]���5�h_,��H��a�'xо�ഥyhJq�v	���5n�-���M�Υ ��!u�HlrE��5e���z� '������.��y�`�2���6_ftArC��`6�Q���ĪF��(��cyjB�u� +�gF4a���]�(�ꭙ���o���T�U�X�n��՚X�9������������!Ӵ4�����'Uoưʽ�{��-nŘv��-��2��W�O�c�S���*��&�_1���exKݻ�t�I�Ǆ�R(�C��4��|E��S���Z?�5�ʢ��%���[��X��������GL������^��b�n����b/��s�Q>���2��mb�WP��?��{��0��_�c[���\��ha��� ���.�օ�� |���f�'�%�ZG`h�}ir,P
���L�C�R�C���_�Ώ�����QQ��JQ�`f�|t+��Y[�r�-����zp��m�_g�"_�u�k��h X����q���U}�g1g��'SQ�	�K�<O���2��P�?�й"��|��C�x[���0V�,R�Tm�5M�F`*x
�ߴX>�g���u*���* ��� .Ǥ^ͩ��F�ݴ�2���͢�2�C*���Vq��h+2׏(H�����b?M� I�E�l#:�bU�e��cު����y�/\���� �o\A�0@�����5�qzx޺����zq�{��%@u����L�Qm�.\���hޝ�W���⭹�yhɥ��gs� " ������i��Tꃇ�*̮� ��^�܉��fu��p�Q	
J��i��jӏ����|쓢*:���b:�5�S��`���K�3K�]��ќ���Ƚ�/y�A�e"7mB�J�u��u9���w!�u\jc��}go��n�Bf��\0��?�[3�����23-�hb�n�cz�����@YYJ?I�拁lH��<�Oۗ��7��֖z<�O�"E��𒙱��%_��|
b���ތ�Ac���!/E�K�[��zC��F|,�H��tx��Xt�w��A����(%���c�BMW��97fV��X3��@/h��@�I;؞g��a5�1���I�!>�C���3E�V�u7�Gr��A����w�?ԛ#�sšfC.�I8��+:����7(�� ��_Cjn�(�G�sE}ƫ:n}ӻ�Gܲ�T���^�&%Y�z���'X��Y��.H�5�Q�T�k�Y�1�@`��Ś��X���.�ʾ.�\��t��t�p�Ţ����3��P=�B�:Nr1,9�ĢS*.H@|��L���:��A�:� RM�����
!����/L����E�`��ר��]ƀ��D�%��G���ӥ���K!�����(����\>b�Llg>b9�O��#��R���~)0����~
)-���E�y*рX�A!r�R.�0��;��������ZFT��i�>�98�b�Ƚ�ϳ�KF��6�$��ʊ�����h,�T��u�H�rkt:)v�L(v���u�q+iy�<H{1��
��kH��]	�Úe��ː�a:c��:���$�,��ې���׺Ẕ"f;�!A��� ���z��1�*�^���N���Ѧd��{|N�YHG�������!�xTL�$���x�U���U$��rBF��p?��O�/����] 2�n[�c?�>�H�eA����|����xέ����x��J�qD6yB@]��0�Qǲ���^�~'Կ�}r�!C�T�H���~��*M⾺�N��F㞵R�Pq1��H��(���'a-�?�|������1����(K�Dؘ!�]���y ��\��ϝ/E|�Z~���x������uqÔ��[_���6a���ؾ��:��$��_Rex"�~C�y�� �,������A��k��f��[�m�+G��/C�h;��{��%��[
��k>��0Q6���\񘐣	_�ϰ��20�N�'�)Ҙ��:�5r�l-������k9����9&�*̈Z�*�<��ʹ���Sz~��	����@
�`9H���5:�����) r��V)L*���f�E[���X�;�S|9kCI��b�"�L�b��HI�h+��b^�[�������,��.G}� ,ꩴw��|�G	��p�Ӆ��eS�+��f�V���!/?S�$��jS���.�$9�Ъ�U��žίC&F*	�^x��x\�/����":�4V��t��#�������#۞i�/�I�R���IxV�\a���VdD�ը=]�@	ޑ��G�,��:��1��$-&�0]x@mi� }ɗ��ek�����œ8{��8����`�Ag#�]ڕ�,f��� P�~A����ÐF$��z��Lf��]@#��G���Ն��\gC��xU��|�N�^�U�E.s�w{Y�B�*�8Ʊ��  �~�s}��x���F����H�O���&�?z� �e���e���f'��duV���E_6FR5����ͫ�P�x9@��}�,y�)�@c�F
�Q��5����zL`s�V6S/k[�w�E���׉�&X(��:�!9پ�\Tqs�y�m4�c�r��a1� .Ho��V�V��Ɂ���/$��{�'���P��p�,�6>5��_�H��
8Q�ȿ���I??i��t���Vs0�ꓵ 9� ������������;�\O0�[�I6�p�Rl�\��i��M�qζ�������^n�� ���]8"ߕ-�t��>�Z����� �?:ef�+
p�C�[��a���>�P�' ��,���q0�op?�Fp"h��{������yn�7묑��~���|�)y�j�Ab�����{̲ �_T�f�ݵ�Ya+�VV��>��$> �9����-0�!�A�ٿ����A�����_�K�,��5 T��
Â�z	0���K�~�0:�K�qb.=(�<[@����{Ic���v��}*A�����B������hV i�6��*���۰Q��ZC9�p6k�lC��	˼%ZR��E�j	�g��4!�����zY���eB�\o�¾Yu��_���	�a]��!`��f�#���o���He~�$�r*"/��v|���;�O��s����^�������Y�t%��X�7�gT�|.~�70�-IvF�;ɳ�	%�ࢎz�<C'����Q�y�p
,o���Z�
#��s��"���̧���ՊaI�V?d��JW�Z|�j5k/��EQuh��^�EH��
�0+�!�A�aנ���g^K�V��1�m�Lz�R�]�x�E�l�WE2���.ذ�N���0

4;�hύL��0��*�Y�E�0U2�/�m������>`H��n�����k�w�ep�%��fU^h|�]����/9���R��nkgq�S2�
��e�#\;�HG�MqQM���r�9��#����3 �J݃�ą�y�x��tnH��u�C<�}Kf�ܦ�OA�ݗ��K�b���quz�����|;@)�qXSs�W��]q�9н�Ugum�
\ҧ�ڕ�C�c���+��ԠW�O�����ǧ����v��Z�Z���̱xFr6 ����"☭;�c�*��<M�^3����Dn�M���zّ�q�.0�0g:n��ćo��&�⺑ V�������Kb�7������/���Uf�<{���Rkh���~�EMk�q0�	��Zu�e8*��IV�e'�:U˟�VW�6��+Ag��<X�95���0�k���Y|��ch�5+1V��\����L���8�Y�n`v$� ��ix`UV>c�9�8]�,
�i�a{�������Ő�!�Q�u�O�J>�T�×-���\��1O���l���'U�#,V|�d��Q"?OG�@�x�P�z� õ͏��W���p��g�t�ݘ�#�K�|���׾�^��"��U��+R��9,�{i�Ƀ�������ldL 0�u�Ǎ�i{���k�����Ͳ[�����M�� d-ю�[�|{ck�|��{�4*�ʇ��9���{�o��8�:��~���Ss����98bR/�8O����I����TX:Xe���Pt_d��3���r�6+8�"�T�װ<*i?3c�l�������+���L�%�$���C���g4D�عf)�zb�Pw�%��i��h��T𱀽�p옖q�􇍷�Y�;��ij�eJ��E1���bi4�N/Љ��I���*���B�#����(�C�ykE��eN��6��O��Z{["Dy�dI���$��2�$��6w��x�9$��ۡǷ��,��˰�e��:��;Z��,H��g��b�@3s#�G�OVL@�I�Ú�X�B�Zm�J8,iR�(W��BJ�e�� ���^��*�P��ߔ�����>ݵ��nPy��`o{,yv;�,�j��~�
���[�{'����:dj��*t6Wh�(�m�/���}����V��O���D�c�
��:{�t�����Æ��wC5 ��}�\�9��&������ �SI8}��~oT�Z�xUr�B�i'b�'&��p���
$y��&Mu'��&�2��U}�=K)&�Ϟ����#/Yᕗ'	��/!0�و}�/���N�Q�����V�@�_���5{�J�&�F+k�������Ľux�ҕ�n�
S)/!�1]�r���kr,�&���7נ^uq;�*l�a(��k���=��K* Y��������jۣC�猀Ř�O�1Y�!�
���t��H\�y�{�����<�OZ4�IxE���1������Gx�y�1R�pr�Qck�8�<0�nV�l�;��5kW�A��,e��+���d���n���Y�5��0t�(�,ϯ&OȔ�,\�/mF�_Đ���u�F�������n&�����d$�)�&�x���YoL�&>�򊢠C&�������х��n:ב���P2�w�91�_��]P�W٭�+���V��8�Q�F=��H��h���%S��ɨ�i���@�_ ����+����r>~�c$����8�M���_�~�ٍ-�]~8�xT :@���d�,�4��x[h��Dc&Uj��ҫY�J���_�n��!�^#SuU�g
�	l	ty��ٰJ�'�@w�
���O�{���P��T03�4�`�goq�����X�R`�ڒ��G��=��O8����%qQ�-�Dz�b�w	��G[�1rex��Z��@�>B~��d%��N��W&,���oUB3����.��Ĳn�9d�"`g��z�L�O�S+�E�vnPB������컘�`#��I��88�2g�,u��&���2{��f���'-�4�R(b}'/L~3�	n������Q���<�KK�j8��x�S[I�o��Ec��'Ѓ68���XC�v��}v��^�QV>a�k��x��~y7�tu_�d��>��n)�ܮ�l.�m�A�9%N�������&����M�9������CŦ�ơ�8���>D�Ȋ�βt�i�JOA�7��I	����'p&�\��R���` �.��s3^�H}.��6�Sz�]F5�p	L�/�T%���L޸�P�'n�<@+�A^�C/��Kh�� � 	�(�![�u&�}���P��2�qO�J�W�uȪ�n��{��8����j����� �*ٓ)-rA��HI41��;�GR/����;r|ͨ��x�Z|���d��ln�Q���(Y�A5r���W�̚`9Gf���Y�q�ه��� $�22\�ƪ��	��@�P�	��q���[.A��[� �zg�z�3E6T��?e��63G���ZvF� ��+���xp��I�
� �kx� ;�:�}�c�g�7��t`����$�^���,֛��Ay���%�\8]`�sYܝC�����.?;߹D�+{�3�7,A�h]EN��k6d���R��=�E;�wv{��A`��*g���S% ���[l�_�`\/���KgD�d����ph�Z���|e�R,([��[" ߏ$�%\u��B��#3э,;��2+=�V��2˙�'�F뢮k�!��P �� �u�a�A��ֲ�P�z�Z+k���0����NNn���&�`?ʪ�q{6�8�RpQ<��_�?f#6N ��;����"{i$OB�b]��t3>"K�%	��ª��7���
n;򃶯�� ��c���$]}"�6���>�iz��"��j�*�HJ�G�pQ�p��l�DE�1�8ҶV��&��L�d���3���^��;�vq�6#��g��Vy�tw������� �	k�*0��K���_������ì���]����+�B@�A�"�#��8�e��,�jl�ab\y�h�����;
�t����)��ro�?ҕ�fc;�Y}�	j#Y�z0���D��Y�Pe�8Z�|u��{�"�.MQ���)�\t�
���ϓ�Τ�NԺ�4��v�Ë^��!�G	|���L�ǟ���� n�{���\���o��DV�l,d��1�ۿ�+D��U�TD�͜7��v�c|�"G|K�U��J�TCw�=;����kp��'���(���;Ļh��/M���V��H�Xc�2)�8��))�*�U��^d�^�R�e5K7+��^%}ē�[~n�xE�>L�;��Va�#����!� ������Ǔ�W���]��/����R�!�\	Nt�M�,�U]�N`�����u��ͪ�B!(G�HR32o����x����1{ˉ	BwTBH ��Z��J�G��ʢN8�˰��У��6���Y|q��&!Y��d�|�[K�J Ի.uq�@�����3�v�hnɃ�M�d_{�f�p_6�O
���X���i{���E0�/�.��M��~�����uw��.xpC��>9�hIN���������S8>�EF!̗�c�U���;5�̀ńr��;x{�\���;��'Sy�=bi�Z�%g\-)��s�EJ:ur\�w�6��l{������!v.�,�4L(�|�f����m=V��u�����z=�xķp�%�..���؍z�H�aF�޿-;�������HP�^�ԵNe�}__i��`ST�B����R4��Y�M�Z޲�A#����"m9)z�VZ6r�%�W�}����`fJEyFDv'7x�¨;�M����f �>ݬeUN_�P�PE�ܖs����S�0>qY5��ީ, fa�^�~}Ȥ�ײ3�;��c� N��ܹZ�S}n��ˠ�ԡjm_�'J[=�Bvٷ��GV�0�ּ�6�������D^)|�6Y��Xu���d�T�E t0�B^@]�1:O�8^(Y��SO�4iG�ۛꨇ����xE�2��<E��u����/o���.iJ���~.Ԡ5��a	��P�������`�HH���k�����g��ymn��MA>��˿5�*��Jԥ�Gڵs��w��s�jM�fTTD����Z\��S�e"1���=�hCu$a{5߱��ޱF�]t�J<G`�P�[��W��=*4�HWM�8�j�%m�4�P�e���s���E�+l�Eol�:�|��!{ik�wK�:�� �H%�n�D[������>^QE?��|e���!�̻p�&�t<m3/��sW�:� �8܇/"�³�()L
q��ε6��LTsG����M�U[�N�dm�F�@@����7#��`ê�L�ŗ߽o?׊�qZ��J2=zڠ<��n[T��B�!sW��)�B����;�Ε��}w�}���b>�����%7�,��x��S�/��m��Z�
��L�G߿B}����bFr�z��#��!�q�p5�X;F�6��p�u�o �2�Kn�Ԃ^A�@����p�������_7��*8Ǽ�r���g�Jr6*�U\��G3:�NIl�0�I�}��&�G�HT�5����2��ZҴ�p���n�y�;�*�K�4�:=�Ճ�b�~���Vh�`��v�
�aTx����W<]��G����0ޱ&�JGM�%dh�S�jh��ҵ���J���Q��p�¯�����螐pl��U���D�;Q����.��$/���Ra����ܜ�H/)��B�"1�5D��ض�B�Kq�����������2JU�J�y��
w�C7��LTb�(��P�W���[ٯ	x?�) t?��Q|���x9���xZ���lm"�W��>�+͸�'RD��j]nr��bG� |�keN#�ǰ�LM�����D�Gv�:��[mɆܸ���،�	��O�]����\UJ(5��?�>u�ND�m���u^J��~��)+��ǃ4��ݦ��۝R��n�1Wh�0�n�=����x˖�mR;=CtW��#���n(p�U��4�\�}Fl̀� � [��oz�5V�E��R^z�r�>F�}�agbRd��9sQ��׀%�|A��r�$�f�ڣֹ�fT�u��Gwo���UR�T�����S���E[����ӄ�i̴�q|#u�X�5wy��Ӝ�'��-��-�ͪm���<"��ڿKnM����A��%1�ԥ��LWa�мw3R{ϮAKd���;Qe����
��Mޠ��iQr��+h/���X����x�2R{iP}c� 6h��<ۊ�*����b�� ݺ㔠Q��e�Wl��ekt:	t9�.������c��*��M6YN�({G�}Ʉ*��k��l$6�]���u~!�B�;�>�a?co�d�)6�������@�績��"tn�9�},��(B�C:u�j�w�R}�+܌�!�E4�s�^��C���p�G�ؗQ�q�,��n[���C_�Z��Ű�\zxht�Z�7-R�����.Bq��T�������s�y� ���഻b@��>B�*��V��jE[�\<�W~�މb���{�ך�*)�Ľуf^d���GT Z/���Ҁ��-�oJ'��t����kp��\1�`�|�
)��t�)%�ߤ��O@�'���.�W�R�F:��8�m��8+�բ;g��EgO����L/3T���`@��.���S��䙅̾��*��q�3�@v�̬	��U���il��4�]o ��r4O4f�������y!f�otYӌ|���?�I&
��a���B�r�B�'���tr�Al2�8nJ�K�4�����g�X]Oz%�~mX���dC�A8E��1q7��; ?�f�`Ū6ql(�^���E�R�1��o~Fn������F� �JG��}�٩��� #5��VwMZ��Nm�M��A#��\`�ޚk.�h���\,�XZ�#-��&�i]o͡d������H���k/�Tz��Zl��;J��_:
��\�����x����-���d�1#Q�y\*)WB�ЦJ��d֋8ڃTf��s>�8����) ��o����<�y�Lk?/�,��8�]0��w0j�[�`����w �C7�p5�����ii����"��߽� �N��]`���W�}&L����Z_�=
<Knv��R�y��1!󩩋�����ӧ-�{m��ӿ�z��OCa����x�=!6`�n-��b���|��b3�{��a
�ؠ�#3�/��II]]F.z��T��p��0Dw7jW��������z䪬�h���r�Aߨ���;:3�9��@���Cs/�E����r�;�N(�M_?�&}��,�y$��,[ ��h�+/�sJ(��nw���g�pK��s�ѻjn���s,�f;�����������]�j.�H���勒f�#�'n�m��̷�82�QJ�m��
�V�D�x�i�������	��:� �0��j���0%���:�;�|���p?�~g%��X��C�m�¾�t�鬓��s$�(�18��sAq��X���K�2Ҽ1~7c䆦�����7��Z�mp��*��b�˔�	ݼ6����p_CLJڐC�Vس�6xز2���P� �e=:q��Y��Ў����^��\w<�-y�MB�M����}����js�m�h�����K&Zf��,2hGv��?��m�N1�I2�=|���b�g{x���l���t�c��a��M��&�o�+������R{2p3��>�<��J@ˌ����EY$=������b���u��Z~	O��J^p]P���=��i,�����b����6(�H�G���r�PG`5|Z�Jj��."��F�ϱ?�g�}l�wbz�{��vXT����9�qOc�|z7�.nFJ ��͞��~����fۨx�j�=����"�FQ����x�+%���+�^K��^���S���߷�[�W��+���SO���l�@#'�>���;:A������]�������g���
��y��`����Ѧ{�1z^����N���t��HD����
�C����f(�;��ܼ�!�	�PA�:ƃ�"2�DUQ�
l&�2^��U�^#��ph�D���	{:\I�rO_B��uZʥa�&�<���������z�ձS��[&�eU�j�	Kx�u�$|�NX��6�b�ߡc�?�����~�S�JK�`de|�H� N�>	�1*c�F�q_�*<Aޡ�C5�	��rѭ^¿�N���gXE���t����r
yP�wRu���g(���W*��}AP���G�qD�5��7�@|���H���;�&��A/�_&?����-�'�|W�3?Ր)�X��3���T/*�_�)�;C�HO3��R�c�i��|�OgP&(;6�G���Ab���f� VQ�eƫ��r{����N��Ɖzxlnhf%��$�q$3+#�}�s�o8����j�J�%7IN�ի3�$�Kƛ�����ƀ��r�܋���鷏��
��s_�Q��ߐ^�2�[�9!�����_amKdD;>^2�u�m�_�<��?>�6;n�o�UGU�"I�&0��x��t��o>Ћp���Ԍ1#&Ģdk��B�����,A��LHI��$�*Tz��A�ȽH|V��h1h����^݃	ʟ
��O�J�t��~��|�g�PX4v< �|"�Ex��|N��k"SB���j�\o���7^6kuP��I巑����N�!�]����c *�/��K�@�����G��AfO��z8o�*b"[Ml�pf���1 P�b�l7�6@����v��AC�%���/�Nj3vֈ�I��TӔ�[M\��M�pR*J5�bha�}Vm�]6�7�'����)v�������Zޑ� ��U��`Â��_�K��;v+�}Wb><�N]Gt*�h�G�̰%.�ѰAd�>��%N�Iĺ�һ��{@(��	B$�Q(�L��a��T����C�����R���vIoa��C*e/��Y�[��/J���p/���@��=5'1"Q�|bi��]=X�����x���d=ͫ�*B=z�Rj{�o�G[����[�5l
�6Y����O�ʉc��~\����Ər��JeIV=���v��#[��r{�@`^~|����H��x���ŷKYh	�۹	��F��i��K^���Ժ�v�XbH�oRv���#8�b����ʵ^g�q&����vAyZ��LK�2W$B�;~IcÄ/�]������8���=puph���J��̓�@��|�Kbx�J�r�r~Z��:W��m�n92  �׍]T����N�˕�@a����QHu6�nXM?ЊO�@�U�D��TS��?�5�d
\�6Ƕ�	�j>��f�����?���L��)P�k��b,���� �t�����^n��x���K�Gc�=��,(��?s~sH2��Y`��%��{0[���%׹z�&����_�B,���d�b�##5�҇I�����MV#à�@!��n����y�8 �h��r'ns��We����$%�L;�;�������U�(��S��OH��V�����=iL[KYj�N��m����|V��uIǓ��R�dS�.��G��Wv�m���I`���M.�iT�x_2캙�Y�?�U�� ����zz�!����k<8 i׋A�MR-n�XB�yH��$�{��E�_�A��q?���=摈t.�'��t/� �:iB���_c1E�bzW��V~�ʾ��"܀.g2�1�5*,�8��Ը�v����O��X�M��³�[���3V l� ��C5'+�\ɿ�MQ�����T�uq�6�2坊� 4��ǳK���.w7�eo��4������Q�eo&�������:��v�KY��Bل�[���Q�pe7 &!�h��Ϸ�1�J�^�������s�xD(m��}��􃬊� -W��^����[��5ʝ��C��eN�k��P+�b�n�/:�C4�sA��}5.������֘:阰��1�)S�i4 p�1;u��W5&ó����vuB��ѿ⏼ɥl�	n�ޗA`��0VܗLnɒNMI��s"߯�w*�˨�[,�s������[�����+��G{��q�{ӵs�k|G-b��/}��F��m�?��%�8�-��w�P�5Vyw����}U�`�X븃��0��	�5�$"�����%�vA��t�T�<�=j�<���'�Î�Lx��T2���Á��(���ѫ�����S�������RCUJyp3��]V����n+���C�D�Q��W��ROHu�A�`�šh�F g
��beD�I-���sq~Re7x��q���0�>D���g��#H >���/{�������ݹ=����*�v5����+Y��B?�F��=�jy*���r��11���X��tR�D�H�Wl��1�dU�����#E��Y$ƚ?�����8�J�g�������j!ڟ�l�C��l�Z�z���n�`W4�KQR�Âw,D�㧖Na]�xg৷����t�n1ƊO�`�.�H�Du���?�����RZ|{�!�Dw��@������V��"�4�S��Ds�Z���r���,��m�?{q`$'��l�vc��Hn���M��$���K|1�J���k���v}�vP�eY�D<�D��Qx�3���4��(� ���ធ�Y��i��0p#��M�T$ܭ����Kx�>��Wp�]sod�Lŭ�_�ٹ%��>�_(���x�����!��K����d����4�$?�ut5}�!�G}k��Jq��`$yٻ�����Mb�y;����%a�!'���Q�77�(���n9Es��h��	/�yM���X�*���V�艳g���`_���}(#!��c��i5�(����6B	��޴���Β�$a��e�J���k�b�A�n�j+����Z�/��]/�^�i�_��rCF�S�}I|{�c�i{��(��H'O��c�
X3l���� Ev���8�AC��%��,RH�x��7�5}�{իx@{zs:�`����������{ O44X0���p���I@�{��n�����	$�x�±�ej󏡣Q=m<��sR�tX��_�`e�h<��,��z�ηJ��;�ݕ�u���Ty��F�:v�~-�zO�TiuQw!"�l؟�C�Q.�Ƃy��� 
�P��=�����G]*�e��B��f��b� +�*�{_��&�n�T h�7Pq�O�h\�N�F����^\����z��R�^��͢�3���r�M�=x�,N���ő9.~T���q��c>��N�Ǘ��r�1��@�z L��]��Y��,Ȓ0e|�Ў%���"}�u	qOH3#��k��[[{y�-"�`d��$����3%�^������7?�_Yv6+�}���ъW��KwE���� �MH���@p���]��ʘ��r���ь󽺤��1��:�ܼ%USm�&ݸ[��_��[��3� L��u��G��V'����1q={�퇖�|*S�tl?=�D�F��x�6��d%	JzNAz	����4��Ѭ�Q�]������ipGry��${�
~�c�<�ɨVM"�w�F�Q��'a+�$iJÄ��a@�Y�n^R�M���Z��C�]�xmt
�,k�U#�z�z*�ݭ4Ԟ���3���r�T�"3a��]���s,���"�6C�z��<z(W+[��K�C-&��C�h����&�W�!�-C٭|�;dP�I-Qz4rC��;���	w�ϗ[�~$��҉��!T$g����0��i�w6�
�c��e�/Ke�=#&�S�e4����,��L�(v���%���M��p�\�'XdHG�ؘ��N���.B� �?u*��4��l��׋���S�V2%�T�o�}�[kŲW:�4)�pTHn� �����9.ȳ��M�W�%藞�Q�3Bqt�ʋ��Q��\pxY8Σ��豣��=����$����Iu���jÂk� DI"5nz�8�CH��=���ru�*�g�n#��u*��mw�A�8t5!*7@2y�A�P�+�f�Q���ʞ�ï�.Gqx#�l��`����[w,���޿Ar��6���C��+��ڍ +�������̖.c�Ʌ��:��u���f��9{8}!��N`9DJ�dzy��j�c��ˤ��3��a&L8��L��Y�_� �K�4qP�}{���|�����0��O��u�b���ֈ��,��R�8���~�����)4�U�Y���Ku�|Yh׸^��q�Z]�o���'���L��.K���
�i�jڌ���B�qLN��v�3��J9�S\nu�]��r֟l�ù�!I:�h�!հ��S�04QTj��V4���[+�8dQϚ�����}Q�L.hM;L�r��U}#������XG��,K͜~������ g��U��;�GKX+Y3��j 4�OtJe��>ޮ��5ט���#dD`)mB�m�`'Z�n}5������E�J ��C1B
��eJfT�~1B�A��~��B��FB���:j�8���Ǻ��G��<���,�;�6}�܌�Zn^*&F�"�%����h�YJ/��� �z�=o��ތ���}"v����������DԒe��w��P�
j�X%G7Q��hb��\���a�N��DP<�T�����J��:ɉ�f1��ռI�a�����Y�C�.�R���{RA{�}m����*D*�l�%ry���<7�c˔����C�� +�HQ!�Q�`���R�t/C�6|_Tw����?w3�HTC��c�hU�{I�hi���}�q�g�(ܴm�c�7���&��*��5`�8