// niosvprocessor.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module niosvprocessor (
		input  wire  clk_clk  // clk.clk
	);

	wire         niosvprocessor_dbg_reset_out_reset;                            // niosvprocessor:dbg_reset_out_reset -> rst_controller:reset_in0
	wire   [7:0] niosvprocessor_data_manager_arlen;                             // niosvprocessor:data_manager_arlen -> mm_interconnect_0:niosvprocessor_data_manager_arlen
	wire   [3:0] niosvprocessor_data_manager_wstrb;                             // niosvprocessor:data_manager_wstrb -> mm_interconnect_0:niosvprocessor_data_manager_wstrb
	wire         niosvprocessor_data_manager_wready;                            // mm_interconnect_0:niosvprocessor_data_manager_wready -> niosvprocessor:data_manager_wready
	wire         niosvprocessor_data_manager_rready;                            // niosvprocessor:data_manager_rready -> mm_interconnect_0:niosvprocessor_data_manager_rready
	wire   [7:0] niosvprocessor_data_manager_awlen;                             // niosvprocessor:data_manager_awlen -> mm_interconnect_0:niosvprocessor_data_manager_awlen
	wire         niosvprocessor_data_manager_wvalid;                            // niosvprocessor:data_manager_wvalid -> mm_interconnect_0:niosvprocessor_data_manager_wvalid
	wire  [31:0] niosvprocessor_data_manager_araddr;                            // niosvprocessor:data_manager_araddr -> mm_interconnect_0:niosvprocessor_data_manager_araddr
	wire   [2:0] niosvprocessor_data_manager_arprot;                            // niosvprocessor:data_manager_arprot -> mm_interconnect_0:niosvprocessor_data_manager_arprot
	wire   [2:0] niosvprocessor_data_manager_awprot;                            // niosvprocessor:data_manager_awprot -> mm_interconnect_0:niosvprocessor_data_manager_awprot
	wire  [31:0] niosvprocessor_data_manager_wdata;                             // niosvprocessor:data_manager_wdata -> mm_interconnect_0:niosvprocessor_data_manager_wdata
	wire         niosvprocessor_data_manager_arvalid;                           // niosvprocessor:data_manager_arvalid -> mm_interconnect_0:niosvprocessor_data_manager_arvalid
	wire  [31:0] niosvprocessor_data_manager_awaddr;                            // niosvprocessor:data_manager_awaddr -> mm_interconnect_0:niosvprocessor_data_manager_awaddr
	wire   [1:0] niosvprocessor_data_manager_bresp;                             // mm_interconnect_0:niosvprocessor_data_manager_bresp -> niosvprocessor:data_manager_bresp
	wire         niosvprocessor_data_manager_arready;                           // mm_interconnect_0:niosvprocessor_data_manager_arready -> niosvprocessor:data_manager_arready
	wire  [31:0] niosvprocessor_data_manager_rdata;                             // mm_interconnect_0:niosvprocessor_data_manager_rdata -> niosvprocessor:data_manager_rdata
	wire         niosvprocessor_data_manager_awready;                           // mm_interconnect_0:niosvprocessor_data_manager_awready -> niosvprocessor:data_manager_awready
	wire   [2:0] niosvprocessor_data_manager_arsize;                            // niosvprocessor:data_manager_arsize -> mm_interconnect_0:niosvprocessor_data_manager_arsize
	wire         niosvprocessor_data_manager_bready;                            // niosvprocessor:data_manager_bready -> mm_interconnect_0:niosvprocessor_data_manager_bready
	wire         niosvprocessor_data_manager_rlast;                             // mm_interconnect_0:niosvprocessor_data_manager_rlast -> niosvprocessor:data_manager_rlast
	wire         niosvprocessor_data_manager_wlast;                             // niosvprocessor:data_manager_wlast -> mm_interconnect_0:niosvprocessor_data_manager_wlast
	wire   [1:0] niosvprocessor_data_manager_rresp;                             // mm_interconnect_0:niosvprocessor_data_manager_rresp -> niosvprocessor:data_manager_rresp
	wire         niosvprocessor_data_manager_bvalid;                            // mm_interconnect_0:niosvprocessor_data_manager_bvalid -> niosvprocessor:data_manager_bvalid
	wire   [2:0] niosvprocessor_data_manager_awsize;                            // niosvprocessor:data_manager_awsize -> mm_interconnect_0:niosvprocessor_data_manager_awsize
	wire         niosvprocessor_data_manager_awvalid;                           // niosvprocessor:data_manager_awvalid -> mm_interconnect_0:niosvprocessor_data_manager_awvalid
	wire         niosvprocessor_data_manager_rvalid;                            // mm_interconnect_0:niosvprocessor_data_manager_rvalid -> niosvprocessor:data_manager_rvalid
	wire   [1:0] niosvprocessor_instruction_manager_awburst;                    // niosvprocessor:instruction_manager_awburst -> mm_interconnect_0:niosvprocessor_instruction_manager_awburst
	wire   [7:0] niosvprocessor_instruction_manager_arlen;                      // niosvprocessor:instruction_manager_arlen -> mm_interconnect_0:niosvprocessor_instruction_manager_arlen
	wire   [3:0] niosvprocessor_instruction_manager_wstrb;                      // niosvprocessor:instruction_manager_wstrb -> mm_interconnect_0:niosvprocessor_instruction_manager_wstrb
	wire         niosvprocessor_instruction_manager_wready;                     // mm_interconnect_0:niosvprocessor_instruction_manager_wready -> niosvprocessor:instruction_manager_wready
	wire         niosvprocessor_instruction_manager_rready;                     // niosvprocessor:instruction_manager_rready -> mm_interconnect_0:niosvprocessor_instruction_manager_rready
	wire   [7:0] niosvprocessor_instruction_manager_awlen;                      // niosvprocessor:instruction_manager_awlen -> mm_interconnect_0:niosvprocessor_instruction_manager_awlen
	wire         niosvprocessor_instruction_manager_wvalid;                     // niosvprocessor:instruction_manager_wvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_wvalid
	wire  [31:0] niosvprocessor_instruction_manager_araddr;                     // niosvprocessor:instruction_manager_araddr -> mm_interconnect_0:niosvprocessor_instruction_manager_araddr
	wire   [2:0] niosvprocessor_instruction_manager_arprot;                     // niosvprocessor:instruction_manager_arprot -> mm_interconnect_0:niosvprocessor_instruction_manager_arprot
	wire   [2:0] niosvprocessor_instruction_manager_awprot;                     // niosvprocessor:instruction_manager_awprot -> mm_interconnect_0:niosvprocessor_instruction_manager_awprot
	wire  [31:0] niosvprocessor_instruction_manager_wdata;                      // niosvprocessor:instruction_manager_wdata -> mm_interconnect_0:niosvprocessor_instruction_manager_wdata
	wire         niosvprocessor_instruction_manager_arvalid;                    // niosvprocessor:instruction_manager_arvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_arvalid
	wire  [31:0] niosvprocessor_instruction_manager_awaddr;                     // niosvprocessor:instruction_manager_awaddr -> mm_interconnect_0:niosvprocessor_instruction_manager_awaddr
	wire   [1:0] niosvprocessor_instruction_manager_bresp;                      // mm_interconnect_0:niosvprocessor_instruction_manager_bresp -> niosvprocessor:instruction_manager_bresp
	wire         niosvprocessor_instruction_manager_arready;                    // mm_interconnect_0:niosvprocessor_instruction_manager_arready -> niosvprocessor:instruction_manager_arready
	wire  [31:0] niosvprocessor_instruction_manager_rdata;                      // mm_interconnect_0:niosvprocessor_instruction_manager_rdata -> niosvprocessor:instruction_manager_rdata
	wire         niosvprocessor_instruction_manager_awready;                    // mm_interconnect_0:niosvprocessor_instruction_manager_awready -> niosvprocessor:instruction_manager_awready
	wire   [1:0] niosvprocessor_instruction_manager_arburst;                    // niosvprocessor:instruction_manager_arburst -> mm_interconnect_0:niosvprocessor_instruction_manager_arburst
	wire   [2:0] niosvprocessor_instruction_manager_arsize;                     // niosvprocessor:instruction_manager_arsize -> mm_interconnect_0:niosvprocessor_instruction_manager_arsize
	wire         niosvprocessor_instruction_manager_bready;                     // niosvprocessor:instruction_manager_bready -> mm_interconnect_0:niosvprocessor_instruction_manager_bready
	wire         niosvprocessor_instruction_manager_rlast;                      // mm_interconnect_0:niosvprocessor_instruction_manager_rlast -> niosvprocessor:instruction_manager_rlast
	wire         niosvprocessor_instruction_manager_wlast;                      // niosvprocessor:instruction_manager_wlast -> mm_interconnect_0:niosvprocessor_instruction_manager_wlast
	wire   [1:0] niosvprocessor_instruction_manager_rresp;                      // mm_interconnect_0:niosvprocessor_instruction_manager_rresp -> niosvprocessor:instruction_manager_rresp
	wire         niosvprocessor_instruction_manager_bvalid;                     // mm_interconnect_0:niosvprocessor_instruction_manager_bvalid -> niosvprocessor:instruction_manager_bvalid
	wire   [2:0] niosvprocessor_instruction_manager_awsize;                     // niosvprocessor:instruction_manager_awsize -> mm_interconnect_0:niosvprocessor_instruction_manager_awsize
	wire         niosvprocessor_instruction_manager_awvalid;                    // niosvprocessor:instruction_manager_awvalid -> mm_interconnect_0:niosvprocessor_instruction_manager_awvalid
	wire         niosvprocessor_instruction_manager_rvalid;                     // mm_interconnect_0:niosvprocessor_instruction_manager_rvalid -> niosvprocessor:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;           // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;             // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;          // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;              // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                 // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;            // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_niosvprocessor_dm_agent_readdata;            // niosvprocessor:dm_agent_readdata -> mm_interconnect_0:niosvprocessor_dm_agent_readdata
	wire         mm_interconnect_0_niosvprocessor_dm_agent_waitrequest;         // niosvprocessor:dm_agent_waitrequest -> mm_interconnect_0:niosvprocessor_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_niosvprocessor_dm_agent_address;             // mm_interconnect_0:niosvprocessor_dm_agent_address -> niosvprocessor:dm_agent_address
	wire         mm_interconnect_0_niosvprocessor_dm_agent_read;                // mm_interconnect_0:niosvprocessor_dm_agent_read -> niosvprocessor:dm_agent_read
	wire         mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid;       // niosvprocessor:dm_agent_readdatavalid -> mm_interconnect_0:niosvprocessor_dm_agent_readdatavalid
	wire         mm_interconnect_0_niosvprocessor_dm_agent_write;               // mm_interconnect_0:niosvprocessor_dm_agent_write -> niosvprocessor:dm_agent_write
	wire  [31:0] mm_interconnect_0_niosvprocessor_dm_agent_writedata;           // mm_interconnect_0:niosvprocessor_dm_agent_writedata -> niosvprocessor:dm_agent_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                          // mm_interconnect_0:sram_s1_chipselect -> sram:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                            // sram:readdata -> mm_interconnect_0:sram_s1_readdata
	wire  [16:0] mm_interconnect_0_sram_s1_address;                             // mm_interconnect_0:sram_s1_address -> sram:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                          // mm_interconnect_0:sram_s1_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_s1_write;                               // mm_interconnect_0:sram_s1_write -> sram:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                           // mm_interconnect_0:sram_s1_writedata -> sram:writedata
	wire         mm_interconnect_0_sram_s1_clken;                               // mm_interconnect_0:sram_s1_clken -> sram:clken
	wire  [31:0] mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata;      // niosvprocessor:timer_sw_agent_readdata -> mm_interconnect_0:niosvprocessor_timer_sw_agent_readdata
	wire         mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest;   // niosvprocessor:timer_sw_agent_waitrequest -> mm_interconnect_0:niosvprocessor_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_niosvprocessor_timer_sw_agent_address;       // mm_interconnect_0:niosvprocessor_timer_sw_agent_address -> niosvprocessor:timer_sw_agent_address
	wire         mm_interconnect_0_niosvprocessor_timer_sw_agent_read;          // mm_interconnect_0:niosvprocessor_timer_sw_agent_read -> niosvprocessor:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable;    // mm_interconnect_0:niosvprocessor_timer_sw_agent_byteenable -> niosvprocessor:timer_sw_agent_byteenable
	wire         mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid; // niosvprocessor:timer_sw_agent_readdatavalid -> mm_interconnect_0:niosvprocessor_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_niosvprocessor_timer_sw_agent_write;         // mm_interconnect_0:niosvprocessor_timer_sw_agent_write -> niosvprocessor:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata;     // mm_interconnect_0:niosvprocessor_timer_sw_agent_writedata -> niosvprocessor:timer_sw_agent_writedata
	wire         irq_mapper_receiver0_irq;                                      // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [15:0] niosvprocessor_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> niosvprocessor:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [irq_mapper:reset, jtag:rst_n, mm_interconnect_0:niosvprocessor_reset_reset_bridge_in_reset_reset, niosvprocessor:ndm_reset_in_reset, niosvprocessor:reset_reset, rst_translator:in_reset, sram:reset]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [rst_translator:reset_req_in, sram:reset_req]

	niosvprocessor_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	niosvprocessor_niosvprocessor niosvprocessor (
		.clk                          (clk_clk),                                                       //                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                                //               reset.reset
		.platform_irq_rx_irq          (niosvprocessor_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.instruction_manager_awaddr   (niosvprocessor_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awsize   (niosvprocessor_instruction_manager_awsize),                     //                    .awsize
		.instruction_manager_awlen    (niosvprocessor_instruction_manager_awlen),                      //                    .awlen
		.instruction_manager_awprot   (niosvprocessor_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (niosvprocessor_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awburst  (niosvprocessor_instruction_manager_awburst),                    //                    .awburst
		.instruction_manager_awready  (niosvprocessor_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (niosvprocessor_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (niosvprocessor_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wlast    (niosvprocessor_instruction_manager_wlast),                      //                    .wlast
		.instruction_manager_wvalid   (niosvprocessor_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (niosvprocessor_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (niosvprocessor_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (niosvprocessor_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (niosvprocessor_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (niosvprocessor_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arsize   (niosvprocessor_instruction_manager_arsize),                     //                    .arsize
		.instruction_manager_arlen    (niosvprocessor_instruction_manager_arlen),                      //                    .arlen
		.instruction_manager_arprot   (niosvprocessor_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (niosvprocessor_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arburst  (niosvprocessor_instruction_manager_arburst),                    //                    .arburst
		.instruction_manager_arready  (niosvprocessor_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (niosvprocessor_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (niosvprocessor_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (niosvprocessor_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (niosvprocessor_instruction_manager_rready),                     //                    .rready
		.instruction_manager_rlast    (niosvprocessor_instruction_manager_rlast),                      //                    .rlast
		.data_manager_awaddr          (niosvprocessor_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awsize          (niosvprocessor_data_manager_awsize),                            //                    .awsize
		.data_manager_awlen           (niosvprocessor_data_manager_awlen),                             //                    .awlen
		.data_manager_awprot          (niosvprocessor_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (niosvprocessor_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (niosvprocessor_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (niosvprocessor_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (niosvprocessor_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wlast           (niosvprocessor_data_manager_wlast),                             //                    .wlast
		.data_manager_wvalid          (niosvprocessor_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (niosvprocessor_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (niosvprocessor_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (niosvprocessor_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (niosvprocessor_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (niosvprocessor_data_manager_araddr),                            //                    .araddr
		.data_manager_arsize          (niosvprocessor_data_manager_arsize),                            //                    .arsize
		.data_manager_arlen           (niosvprocessor_data_manager_arlen),                             //                    .arlen
		.data_manager_arprot          (niosvprocessor_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (niosvprocessor_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (niosvprocessor_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (niosvprocessor_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (niosvprocessor_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (niosvprocessor_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rlast           (niosvprocessor_data_manager_rlast),                             //                    .rlast
		.data_manager_rready          (niosvprocessor_data_manager_rready),                            //                    .rready
		.ndm_reset_in_reset           (rst_controller_reset_out_reset),                                //        ndm_reset_in.reset
		.timer_sw_agent_write         (mm_interconnect_0_niosvprocessor_timer_sw_agent_write),         //      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_niosvprocessor_timer_sw_agent_address),       //                    .address
		.timer_sw_agent_read          (mm_interconnect_0_niosvprocessor_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.timer_sw_agent_waitrequest   (mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest),   //                    .waitrequest
		.dm_agent_write               (mm_interconnect_0_niosvprocessor_dm_agent_write),               //            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_niosvprocessor_dm_agent_writedata),           //                    .writedata
		.dm_agent_address             (mm_interconnect_0_niosvprocessor_dm_agent_address),             //                    .address
		.dm_agent_read                (mm_interconnect_0_niosvprocessor_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_niosvprocessor_dm_agent_readdata),            //                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid),       //                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_niosvprocessor_dm_agent_waitrequest),         //                    .waitrequest
		.dbg_reset_out_reset          (niosvprocessor_dbg_reset_out_reset)                             //       dbg_reset_out.reset
	);

	niosvprocessor_sram sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	niosvprocessor_mm_interconnect_0 mm_interconnect_0 (
		.niosvprocessor_data_manager_awaddr               (niosvprocessor_data_manager_awaddr),                            //                niosvprocessor_data_manager.awaddr
		.niosvprocessor_data_manager_awlen                (niosvprocessor_data_manager_awlen),                             //                                           .awlen
		.niosvprocessor_data_manager_awsize               (niosvprocessor_data_manager_awsize),                            //                                           .awsize
		.niosvprocessor_data_manager_awprot               (niosvprocessor_data_manager_awprot),                            //                                           .awprot
		.niosvprocessor_data_manager_awvalid              (niosvprocessor_data_manager_awvalid),                           //                                           .awvalid
		.niosvprocessor_data_manager_awready              (niosvprocessor_data_manager_awready),                           //                                           .awready
		.niosvprocessor_data_manager_wdata                (niosvprocessor_data_manager_wdata),                             //                                           .wdata
		.niosvprocessor_data_manager_wstrb                (niosvprocessor_data_manager_wstrb),                             //                                           .wstrb
		.niosvprocessor_data_manager_wlast                (niosvprocessor_data_manager_wlast),                             //                                           .wlast
		.niosvprocessor_data_manager_wvalid               (niosvprocessor_data_manager_wvalid),                            //                                           .wvalid
		.niosvprocessor_data_manager_wready               (niosvprocessor_data_manager_wready),                            //                                           .wready
		.niosvprocessor_data_manager_bresp                (niosvprocessor_data_manager_bresp),                             //                                           .bresp
		.niosvprocessor_data_manager_bvalid               (niosvprocessor_data_manager_bvalid),                            //                                           .bvalid
		.niosvprocessor_data_manager_bready               (niosvprocessor_data_manager_bready),                            //                                           .bready
		.niosvprocessor_data_manager_araddr               (niosvprocessor_data_manager_araddr),                            //                                           .araddr
		.niosvprocessor_data_manager_arlen                (niosvprocessor_data_manager_arlen),                             //                                           .arlen
		.niosvprocessor_data_manager_arsize               (niosvprocessor_data_manager_arsize),                            //                                           .arsize
		.niosvprocessor_data_manager_arprot               (niosvprocessor_data_manager_arprot),                            //                                           .arprot
		.niosvprocessor_data_manager_arvalid              (niosvprocessor_data_manager_arvalid),                           //                                           .arvalid
		.niosvprocessor_data_manager_arready              (niosvprocessor_data_manager_arready),                           //                                           .arready
		.niosvprocessor_data_manager_rdata                (niosvprocessor_data_manager_rdata),                             //                                           .rdata
		.niosvprocessor_data_manager_rresp                (niosvprocessor_data_manager_rresp),                             //                                           .rresp
		.niosvprocessor_data_manager_rlast                (niosvprocessor_data_manager_rlast),                             //                                           .rlast
		.niosvprocessor_data_manager_rvalid               (niosvprocessor_data_manager_rvalid),                            //                                           .rvalid
		.niosvprocessor_data_manager_rready               (niosvprocessor_data_manager_rready),                            //                                           .rready
		.niosvprocessor_instruction_manager_awaddr        (niosvprocessor_instruction_manager_awaddr),                     //         niosvprocessor_instruction_manager.awaddr
		.niosvprocessor_instruction_manager_awlen         (niosvprocessor_instruction_manager_awlen),                      //                                           .awlen
		.niosvprocessor_instruction_manager_awsize        (niosvprocessor_instruction_manager_awsize),                     //                                           .awsize
		.niosvprocessor_instruction_manager_awburst       (niosvprocessor_instruction_manager_awburst),                    //                                           .awburst
		.niosvprocessor_instruction_manager_awprot        (niosvprocessor_instruction_manager_awprot),                     //                                           .awprot
		.niosvprocessor_instruction_manager_awvalid       (niosvprocessor_instruction_manager_awvalid),                    //                                           .awvalid
		.niosvprocessor_instruction_manager_awready       (niosvprocessor_instruction_manager_awready),                    //                                           .awready
		.niosvprocessor_instruction_manager_wdata         (niosvprocessor_instruction_manager_wdata),                      //                                           .wdata
		.niosvprocessor_instruction_manager_wstrb         (niosvprocessor_instruction_manager_wstrb),                      //                                           .wstrb
		.niosvprocessor_instruction_manager_wlast         (niosvprocessor_instruction_manager_wlast),                      //                                           .wlast
		.niosvprocessor_instruction_manager_wvalid        (niosvprocessor_instruction_manager_wvalid),                     //                                           .wvalid
		.niosvprocessor_instruction_manager_wready        (niosvprocessor_instruction_manager_wready),                     //                                           .wready
		.niosvprocessor_instruction_manager_bresp         (niosvprocessor_instruction_manager_bresp),                      //                                           .bresp
		.niosvprocessor_instruction_manager_bvalid        (niosvprocessor_instruction_manager_bvalid),                     //                                           .bvalid
		.niosvprocessor_instruction_manager_bready        (niosvprocessor_instruction_manager_bready),                     //                                           .bready
		.niosvprocessor_instruction_manager_araddr        (niosvprocessor_instruction_manager_araddr),                     //                                           .araddr
		.niosvprocessor_instruction_manager_arlen         (niosvprocessor_instruction_manager_arlen),                      //                                           .arlen
		.niosvprocessor_instruction_manager_arsize        (niosvprocessor_instruction_manager_arsize),                     //                                           .arsize
		.niosvprocessor_instruction_manager_arburst       (niosvprocessor_instruction_manager_arburst),                    //                                           .arburst
		.niosvprocessor_instruction_manager_arprot        (niosvprocessor_instruction_manager_arprot),                     //                                           .arprot
		.niosvprocessor_instruction_manager_arvalid       (niosvprocessor_instruction_manager_arvalid),                    //                                           .arvalid
		.niosvprocessor_instruction_manager_arready       (niosvprocessor_instruction_manager_arready),                    //                                           .arready
		.niosvprocessor_instruction_manager_rdata         (niosvprocessor_instruction_manager_rdata),                      //                                           .rdata
		.niosvprocessor_instruction_manager_rresp         (niosvprocessor_instruction_manager_rresp),                      //                                           .rresp
		.niosvprocessor_instruction_manager_rlast         (niosvprocessor_instruction_manager_rlast),                      //                                           .rlast
		.niosvprocessor_instruction_manager_rvalid        (niosvprocessor_instruction_manager_rvalid),                     //                                           .rvalid
		.niosvprocessor_instruction_manager_rready        (niosvprocessor_instruction_manager_rready),                     //                                           .rready
		.clk_0_clk_clk                                    (clk_clk),                                                       //                                  clk_0_clk.clk
		.niosvprocessor_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // niosvprocessor_reset_reset_bridge_in_reset.reset
		.jtag_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_avalon_jtag_slave_address),              //                     jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_avalon_jtag_slave_write),                //                                           .write
		.jtag_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_avalon_jtag_slave_read),                 //                                           .read
		.jtag_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),             //                                           .readdata
		.jtag_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),            //                                           .writedata
		.jtag_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),          //                                           .waitrequest
		.jtag_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),           //                                           .chipselect
		.niosvprocessor_dm_agent_address                  (mm_interconnect_0_niosvprocessor_dm_agent_address),             //                    niosvprocessor_dm_agent.address
		.niosvprocessor_dm_agent_write                    (mm_interconnect_0_niosvprocessor_dm_agent_write),               //                                           .write
		.niosvprocessor_dm_agent_read                     (mm_interconnect_0_niosvprocessor_dm_agent_read),                //                                           .read
		.niosvprocessor_dm_agent_readdata                 (mm_interconnect_0_niosvprocessor_dm_agent_readdata),            //                                           .readdata
		.niosvprocessor_dm_agent_writedata                (mm_interconnect_0_niosvprocessor_dm_agent_writedata),           //                                           .writedata
		.niosvprocessor_dm_agent_readdatavalid            (mm_interconnect_0_niosvprocessor_dm_agent_readdatavalid),       //                                           .readdatavalid
		.niosvprocessor_dm_agent_waitrequest              (mm_interconnect_0_niosvprocessor_dm_agent_waitrequest),         //                                           .waitrequest
		.niosvprocessor_timer_sw_agent_address            (mm_interconnect_0_niosvprocessor_timer_sw_agent_address),       //              niosvprocessor_timer_sw_agent.address
		.niosvprocessor_timer_sw_agent_write              (mm_interconnect_0_niosvprocessor_timer_sw_agent_write),         //                                           .write
		.niosvprocessor_timer_sw_agent_read               (mm_interconnect_0_niosvprocessor_timer_sw_agent_read),          //                                           .read
		.niosvprocessor_timer_sw_agent_readdata           (mm_interconnect_0_niosvprocessor_timer_sw_agent_readdata),      //                                           .readdata
		.niosvprocessor_timer_sw_agent_writedata          (mm_interconnect_0_niosvprocessor_timer_sw_agent_writedata),     //                                           .writedata
		.niosvprocessor_timer_sw_agent_byteenable         (mm_interconnect_0_niosvprocessor_timer_sw_agent_byteenable),    //                                           .byteenable
		.niosvprocessor_timer_sw_agent_readdatavalid      (mm_interconnect_0_niosvprocessor_timer_sw_agent_readdatavalid), //                                           .readdatavalid
		.niosvprocessor_timer_sw_agent_waitrequest        (mm_interconnect_0_niosvprocessor_timer_sw_agent_waitrequest),   //                                           .waitrequest
		.sram_s1_address                                  (mm_interconnect_0_sram_s1_address),                             //                                    sram_s1.address
		.sram_s1_write                                    (mm_interconnect_0_sram_s1_write),                               //                                           .write
		.sram_s1_readdata                                 (mm_interconnect_0_sram_s1_readdata),                            //                                           .readdata
		.sram_s1_writedata                                (mm_interconnect_0_sram_s1_writedata),                           //                                           .writedata
		.sram_s1_byteenable                               (mm_interconnect_0_sram_s1_byteenable),                          //                                           .byteenable
		.sram_s1_chipselect                               (mm_interconnect_0_sram_s1_chipselect),                          //                                           .chipselect
		.sram_s1_clken                                    (mm_interconnect_0_sram_s1_clken)                                //                                           .clken
	);

	niosvprocessor_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_reset_out_reset),     // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (niosvprocessor_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (niosvprocessor_dbg_reset_out_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
