// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VPOJZoVHaLfGp29foJWXYPCBO9pQ7A2Oq8bBGciHYzpcYoXuFzXDZHv+eixeui8JjAJ30eJoT9K4
9d7pYfbm0ytX2P4u5J+UjvxSa9X92MtvKQlFZKB4RD6it4UxC6NiU+SR6d/5F1BIuj6hR0fGBl4W
ArHIHu3Ef1szirc2pwYt3wKfiS6t0Fs2xuOsNAxg3olGsPPPdHYyF20IUBr59xhi8yfAoNyWgo3C
QkPgU1/6+NMTYwYtYr0CZJu/Xz0xdTAgbVljhjB9fcsFvhiR0UPiyqpWmAOIbT+j9sTFCIkziNl/
ydQnYcOUMzvWKa8WSaOcoBIkYGKTF8WR5fgLsQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6288)
pzqjNwrWghMHnyGXPRDFuteq2zx09fsyjyY/CHjEFIH7t6jrgqisUsa71HFRQrTiYCZUUguTanWc
Mq75K+aI86yOf/zN8MdCUSagZFoGjHY2XFFeKi/K4k7Ak3VUp6az9zxP79TxwakJQL0GsdLbtNem
pvsa+1f6SPftiEbB0k02/MIzUCYYGiRifVxEgcOJJlDEw8d5gxWOUNJGGdfeHOa/FZn3B/GiEg/J
r6UX9AY0QE+7dCb71ajsp2c3irTCwtNHWx5j7kepucVhkAezGQe4BINWF+lswRx9PC8oRBwxtBpT
umgw8pGC6pMwHONBmeC2H6c2tb4D7Jltone6/9xeHN64agJrn/v29yYrUTy+8zNaeLqnXPkh5B+S
OGN9NgI8o22Jpp6M/hcBFAp1Kwv0fp+kogDLz0NU11xef9MDHbS3h5YG3N59DBoctoTN7HBJ4nB6
K2FN1RoIuBP3GazdZ6BfOOQ3FigkEocV+RrBMiZJcLvX7cQquxfQrgUerUsc3w9uZZ4dSgWyDiR0
JY1kxlMWSKv0ChDVd5xLfh2n5KzQsMLKtDnw3KA/ARQ5uRQEVoBPsE9hnhnwJ0k0lEuSD9IKUc71
Q4Wf/uHSnwn9YM72k//pI+MgJslsL2p/iXeCCwJl4n081GLGxe9rPKEA3BSTVjPsmwhIRDSSsHDk
dOzfNt24qpvFhsHBAUDa9m8pWHNWTl8WGE+QO5BmE/RYP4Cg1F5uFCXr5QwCG0pmBD102Omj4hNl
eheev0ZC4X98t5bGgzCpvFcVoaZvfU1FSsDUFYpNo53AKYhalpiGYT8Pfd+jdrK32ZdHahNU+69o
nH517+BJnTmMqOXYWBmHd1i9h1QgZxy9amFwSQpIyfkcWcVOMrze5zsvc5dS0M2LRMPHNciH2c5i
cPLrACwR4QFyelkUtiM3S7HSVciZ2T0keVjPYMWlHZZ0+J8uwtzE5ZV43EPE4hAEgci6zNpyYEVS
B6T2N6puuALpUjMZ/uglJ6ayDtH53/0yC6OnWl3aaJNKpGFRjB+vlro3xffQwJnqKmReC5vZnzo6
kzHquQlql55/PZxld+uS95zVBtFKK0W+dH9bJ9dg259UZD1wkwJfTLtO4MyDwqRIZoEF2MVlVa55
6ggxBceo+VTKySADueHqW+7DEZCa5cmdodLLCOI/rTflbOx2mlEyI8N0XmaA2WZ6fQIWJKAPCTGe
Zn3vrbkyMHmZWWKmmWTpPA51y5UZ1uuk+i4mgR9beSW+Wza9Bdc7BuS+Dm67NtvyieUdmkJI78Yc
LolJfpq0jzQz5Ep+b1INGo2DZS4WljS1+vY4mfTxe7lEmrXrLDAIvOdcTp57KHz+xEceC7hOcuSx
/FCQ+gk3mf+xPI7YGJSbvpEq6AxC5ENDCzaalatBAzwlW5fKaOBAZBlWEfiQDrR3jmNCJ1yeyg8u
6fRWjrfdH3ixbTBpXOfuYm91XD7c0B7RRu3sjme/U/WGYsKjz48tDj2HdulE0VCuVvnY9li3Iy+i
fC7Ie+I/JGGAnjlTRZ0Cjhvdh2fellgOleI8vPLeinSkKuz3DHd5qeoTyvazSEORIYSqNdxg2fcK
4herfSEkllAX7QboU8k2glRq6CdJ93M5zahfCwXj5UdBW64H4TMitTnScDRK3Er2wwrfG12v4czU
lp8ZziFSbqm0Sv/0aTWGU5mNKbsFKPy7y343PPB6SyPsf5dqdhx4jcVrjzpG0kl9vVy/n7sBymt7
/3u+cb0u27owsWS7heUbWVmErzzgbiBljdrrWJ7USS5gGNRrI6wr9K0uv2bAg4WnBgLKPoX+JcIH
fAZ5rEamUzTHzej704F2XS6Wc6zH9lDdvJCKU/1mTDhE4+iAkMUgMSkQfOj9tQWRHbkc9hgPoI2u
XpophMkyKb4bkrUhJveVmPW4CKG+/Ly1TKo6mb5BLYvuJAzvN7IPPJm0/CXfarPNCs00t0tXdK69
vNncDHDf0DnjpmxkYFF2CrvrQj0UHFUuTCAjttC2CZmh1smvemfizE8rTFQyHlNz3+wj21h56oF+
hjpXgSaGSkC2+Ty8SIXTeE1rOVjKZSFxR0IM5f7P79uhlQLdVRSziZKtWSJgYC7LbwncizKMIWRJ
/V0Yc9PLAoRe+a5rGQMuOApI2b30Gau1dgJrCiEWkIv1/+ToXiBJG1LC/0X1ygoqBFLEwd/STHrW
DYMKPXNjIpJbuKua+KTZ9L6nigdMszhWmEApfnvTK9zLLqWDOhQdNIGXuBVdnpFJCxgOdtYoHbjA
alOJ78jj3wKTvbRxRy+oSo78Rj9+pjZrcgh49Zp3gAeQjIfd2fajB+191ANLOMwCPwdvdf6KbHam
uyd4IctxGLQ1Lc+p7x/yxFLGbNjvqyhLFt2dVqSJq4k4LeNuhsLwYKzgaW4Rdvj51Kg5BbQW7rQB
Xbjhh528aI/nlPyP09qRZkB/BT0Jtq3ggzBRVT8x87HynX6aHOMm6fUZZ0WrOmzRQ7h6iUuOlyDF
bG9VPziySVrKI3iYv7N1dJlO/b94Uwf4cuHrFKHNV5k1/vRfC4cFLaeu38YvYYkMaEuDUmgQTCvF
TExbaMoAVv54I8qOaI76iCZEOf9aMoLl9Yzed64L/D+ipwrg1RQ0ElbN0EHi5NMs2LFmtPyGHZXD
aGnvSj6lQCX5aKBEhZikQXdWznchJ4jvYRes0eGHZ2pS9yrZCkIIrYRAAiI9Y2RvkVvElgCEr/65
x75F1UHv06KR+5BPeXHnr7TO1XK962nqqsGochUWU5nF33Xx2VboZ4pBk3n0GiTHz/JKk5+ZA/6F
ejoiTqR8Hhav2QsoPYAVxDgYOaE1UFlD+sFfwwqQvxieLRGCjOrWCO8AG/xtTy1g4GevC7kWxTEr
cxIbh6csOVFvCEWMP0AahHG1euneY8AOJ6eR2jGl4Wxo1gs9GwKT5ilgnUW8IXs5r7LlcOW1OT2r
y1dR1yX9SN20MZXgZfl6gc1kLzDKwuWkoUsHR/X1s0CJOoKICqPHw14qBUaXNc+Y+GPdZEHFc1vY
GI6TkD+QuKCpsBMNJsFKRhqwpllFPJuPMdxF152lpqloBHjbAhg9njg6ReP9pe727kGFhwJ1x5QE
tDYT1FludWn46beCcT9tpRp6JBd1VswLAIC53ZI0RNTb1ziWHZZNYyCw6Vk5lgt3L/8NszAm2Utm
b3B1JT4hJAuX4pznAR7v1wte9fpNpWjVAVHpnQOOyH5UvnWHiW0Svt/raHpq343WNNIuTN+GmoI3
M6Y4lhOKEfiez4i5hhYul0TXrWkofEzdpuC0XoxeL1AKIS0mUy/COd1jersumsrq7Nt1PetW4z6b
AiYCVQUd/gXWYTZVVMIqBhha83eItYUyLnPPw00Y0GJ3A0WkOvZa1Smv5rTxvGKIY64lePWb7l6y
SbwQB7y/L2Z9BBbpY6axS9OoDwOcDJTWDdfle6jgyisFAgENBXRkMYHvHs8p4AhRbhY9PMislobq
nH0MXegkAhqp6O8O+xv3cmBN5FGDONYSucTdoigvEtO/ZEXzUokf6mpIAsdPyqSX/kibol5HS0Yw
7vZ/Z1i1lXwRbsjwB6aJakmHAiDg4blQTFbBhLxIexTlSC+i6PCrPYAG/XGOhzkAk2zsrt8ikxNt
GPXr7q9/s/2T4PXSc98WXKqLodiepR/1nIyZkD/DA/wrToPOP4402/kJksg7X5rF+dvCHw/PauN7
KQ4ts3rllgTl+iZdS1KFuahUwZ5rl9TaIAIIIHY/VJfiWSyB6R4oPBNyjgHZvlIa7qMWVMFpyTG2
YlLV7ZXzUhVNT1lGZ6sPOHlfCBUqhNufPBr3mdnswmV9yHLtESx6UZA1TSf8qLkMt6tS6Yl2k1NO
DBeai8oRwDsafLlhUoTWyh2+sYPDQoCcQQrTxv1qNkbn65wFN1L/3WOwkszuSZl9DeaEmdH9OpHQ
iHjr9MpCAtQakg3GDjrf71a/z6Ovxpmcc2TjF9j6r5Q+xmX7C1iMbiJyU8ecrPY98Y3UGQ6txmQU
D3tZFSIw/d6J5FRlgJvXwjRWp/gEoZtRX14PNji5U6js9a+XafYTTABTtsnLUXipAYXAgGmRORqX
GZJhb5z5cUDCu+ZGxjE/sG4CbkbPtaWte+CESoSl9HbTAuVcpUpp9T/yBP6D+VkiA8fgSv3Uzmc4
1UNsrobH1q4y3CETtWf3brgUI4yTQAGXoOfFE6ET3+OgbbcFNNFWmKA7lcFGtqX5/nFX7DQQKis1
C22/28Y83mofqhWrlFer5IPaZZYikb6STIHfKDPVOMUQ+0g/Lf3oT5VAsbPBBaKTF065Dv/DGio4
SBTzYb7fkCPNMtpvBbb6+BQQI4Pa6uNnn48/0q54YEUzJmWHf2Bzqwx1mpEPwgwgjoxDkSkdXf9n
pY4eN8JQDsHCsjh+slBC2mdlnrzvAI3vNbbAXvoAJIVMatQqUJMWQ8UdVT2xho7flutJjzE9PBUu
h9zOClaGpBTbTJyGwsCodFrLGke8KX8wCeWRnapMBZVChpamNCwXQqyjC5rJknTP5nOUJXS3MMSV
A5rug/Vo9fTED2zF1mg4soTRorMDWY5EOhIl7SKeEBt6aXxcR4lNs1EfQW/Hrdgt5dKtViGhJela
jDUd1fDfjoGCwDHYVWpdJOgRiBE5L7afxUiab+pBwFMaAKWFUnuXVDkwlwLDjn+IJbjT6oMenQbR
LpMCVrMW1HoZ0/R+gHCnVRSCT+XwZPLkYCDd70FmvNJQiybG62DfW1+Ws0amlPGfc9pwuSvbTkJ1
yZ1ca9C9yJ7L+S4As/tRy6t5D7zHpQTftkyUeaLXqD4xH8jdZhwHWlmy4E6VCp/+MTUNZU9vtp+A
dGAlq22VcRtZYBF8d1nvNI40vVCqoKRr6fGfAP52AcuOl3wCrOlrszMGHjwR8KXXVcYgdaul9Fio
qQJgQ3EZdtb2TS5Q5P78lq6HP9osf+NmFuZWSpb4ys4k9yuBy2pAAnWB02LR8Pf/Fn3Y0sQJe6jq
RXRmfpuhABIA1+OL1Kldeg1ZyLSERnVQxRZswkMdWFn/d6q9CCQYiekpnGaWIti2vF3XDRoxD2T7
lpE4jg+nvvg3ioFZ7g1NzjtufaDddJ02JEk3vD/D6LDS3318p9iiDcOwvOzqmPJqc0sAx1i+i1Rr
8Gg4pIDsNxuczTN/WvTnfcXbugvdgSt3xypfkd2xf1PT47Xewl47dFYABWX5+WtZt6Q2v/J3D6xU
aUHj9IOaD+WwulhQRq8n2zQ3/Wvn3INh6txoZv0zfm8k3jxOLOuMApaxhrPNfdWSPL70FWg24ykG
2EBrlFtDPeqP8Wpb4VG4Zeahv8Y59UsyCat9TNPSWKNI7aUf0J1r9xwzA1O+0+zYEt75fVe9hsuh
Xvc6gT73eIGliRv27Jced/TBPkELUMLKa/K6dPzR5N+RSSnbxp9asARbNc38txvmYx0IpfBttLaK
Pu2MYE9H4gyQ/nrzgUPga/3Tg90ZWXJrjdGHq0zPRygFvtRiKlk7hO4fvbXD6pWTX+ZUIHGrQtVE
TFx38+5jxeEVm8WgNxdZcy4YmHluSRjMUMYJ8x/Xw4MYrLLVkgP5HsLjtmO6jNLnJ/D0vqvYDpWs
HvhiIFlMeNCUsVwLG1jIWayJcpDQLP7tLKIJLKHB6OmV1W53GF6MXc+ArJoBz8ajOgyaN29hiolZ
mapEXylimrNIOvzN1IxnV8DGi/5cQ3HjC/F/0vnRU8nR6MUHEMGRFw27f5jYtpS2OeQdLrmwpwNn
zR9DxMFjyKPpHcthAyj0RdsQ6Rfop1fk0G9xzqcOI2n5OYAU1VOgX3rbgNODg5Bk4EIzPm+hyOjg
S2QvmbSfKX5rpLDXvKdU8GEuOoI5RZy3BOC4mP+pzTWbBgIiCokvA+KMIA3tQMXsQvvAh9XBUEI6
eR5DZFiYx04YOta9nEWJLGGwD4h3dh6f7b/Qspmvm0TtsJJi61u22llTQRYUvcRoVWaBu7hzYsuZ
xcD+USm5sRJrO7/CHakvJtCFnqqvpc2TVEAHoYy1Oio0jY4yVcSo0FzAq0vTPLUuvHgFyYCqn3rv
BgHhMJICKl8SPmC5V/AYZ8/kSbFSUPB5e6cocPjqgGinNHd0cmd9YlHEwCWgvsStwpj1eHOkIaYh
BtnBY6b4e3SCnQ8gDMHum9dE7UvX/2UXaWJoAiSgIi9DIH5QhJBQDVQfTZbCnSp1h5Tgi7SZm+uh
DHBJ0+pL07e+1a7RVqOpeGxVZlpuTQgP2TPT8hxaslHpONYiSR43T+O8nbOZvOoCM42SRpnFKz7Z
v+oMrrk4nvQuzuDn++vXgF4z7BbcsSR8KoDLx3vBnPJ1F2O5iG83BD+y/8O++KiJtIhGV6jrEqjc
a8TxqgUNrJ/zrqYXEPp4PtyhSYHFAvTLKcDIiHYKL1rW+YpQm64cxKUBEGJKo0syRdJX6XSmqww+
xuZ+zyj7A3pliEXJ8HYc+Ygh7Oc1Em1YOkcfSWmzyCBxOXEg3NDpHHXOmbGGViyVTV6oSvJPk+GB
qoOfK4pooWbCO/0znrgEiGjAT82ma9h/jOn0UecKr30/lJt1WIjrxSoZ8TdV+Qvi2NrjSUcdv7zZ
j2J75+bsxcQ84WPJW9LmuEg3povc27sG7X49UO73hGaSwKVkHT8b4F6NZ+5RPixamRWTV+tGbDI8
x96dH8HjR9PjeHinzsXEVEdmG1R+aPXaMUaAMdNMsX3zoUjUln8vsFPjyQSOrasqbxpMQy+Hf4tJ
j8a3NxlzTbUa1/JZUgfsUkaeBmI7vLeyXOXU1+6KwrgWKsO/mJ7QMrc6OklLFoW9QHcZnwUV58SI
b9svVoWm2PNEAnjN2AKfg53PdKjvRNL8y8m1mNIX+c8scPbUjd8RgAO/Q7TRrqu3AS1FuiNFYIKx
gsqjdOGFk9CX7ElrMMxX/9LNdA9Z9iQuzbkmU3zOSQs2M7aEpTb2+ZciWLiM9xYCa8Pfikhz2DT+
h6Un4gvJpVAZw/XHgwBPacvpfePv/3Z/AFrEZ37HqMA9r9h4zmY01Wpgr6MAC+ohXatgU0NpV3i7
eitBXUFqqUjiQbsXcLFZ8sxxBMVROH4Q07BHfTK4O+BbIittyvFGHAU0VRczQDhha12S2FGPOwq5
+h2rO6M44b6Em1cenkLeJYLO7s2KTmLIqj9VyqLEBQQ336bX7BwmH8A5RRdCwMH3XJzp6DQLI3CX
DjNK3+Xz15hNxsnIMn/4jEW2lTPzSzRQoJuno//dxwzX4g2dY/s9/OiS5Q4Ue0ccagh/fmOEyHQO
FtHyz8U9Z9B9ltOHo9kWyWS0bwXCw9KOhktnu7rYkabx5OHHWCrRCYnFLyEY9byg2h+x6gr3+Nbg
A8xeqvuCHnc+9vGLhqPuckMj1ySY35F2bKFQaF53skM9JEubXPG0ESKJOGPhZzIoB6aYCmPU7+r7
K2EBQmZENYP6Onfq8wgxng1zxFb5IWahkRNQ13kVUwc+iLcFzNs5iReveHnURw863WgKk07l/fjH
hdw0FMJc5egB6D+QrQw6lmE1KRsZqDHnGnrdKhh0NFwopkKHhCKT6qvp26gEzCqvxCQ8PpUlyGil
sh89dPPOk1/gUFHvv7GLXanLaLKndffrX+Ui27z40vw9UnThasEfqOvIJV6ux+H+52hS2LCFx1bP
vX+gooTCGF34ua8zSCoMJJbCGz20wvSiREUGfY4MbvTT013mxTsbF/I+DxkyoYIWLnxvMSPTH7P4
EG9uEgKuF+Tr7sVklqk0Yg7eK1w8oF132J273WDBO7JlQl/HkpfVhUu9hCUqCj1rGC2e8iibh+2m
jvR2NCXDRQEcSm+Wn3axFVRYr4V7VkQ3Ts+0AioSns5WdoEMPsoljBCk2ruEAn7focVS678/OhVJ
a2D2vst6WpH0J4i/cH5pLvgIHKcqG9/etFnNdkunsOWMiUBU5wjx/JBcNThXDC+7tAG5H58mOUi5
vqcHmaCdDYq4Xl1i/86sL/Aow2TeADWvHtdDY1czoRnnTStYGillta4bQw3J1HypUwkqOfFbLytA
VEFxjwmxTB+49TkfqcnA5uQmQxQJno55Ncwv8eOgIe2SV5J2+ZoUUKXFVR5bktnirvRXRYV4gg3O
6pHH4eJszfUylhReQs45pUjAWo7QkGi+CPUU9HMR1mSXmdJHCOQo5irnF8+1BJn/jWVRmBLqCQjS
nMKkERCcBI+LC2lpSVei4NyiTSRF/O902F6uhIaBgJkAMeKf9DXhoi4mXGPj4LESqg5awnFNNj+y
NcZ2nmzdcVw4F7bvhJfhySmM0gxTJMl+qhGGu9p8HkduCEQ/4ZziNOAmYybxsjg00/4UpJS5NKic
UEdU2ckiW8WU1eoVHhmKEb0p
`pragma protect end_protected
