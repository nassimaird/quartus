`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g4cv82Ompr8+ctF0O9WrgFoV1myD14Oygmge8NkwDh2I5Sg9F+2Gpu2M1zRaTygT
5VmnAchzh9TnSRPvRDpFVdQjP0oDMe/g9Z62w88OG0mUQyWnHd9ZhbDA0g6f0KN9
Y7VWqRDQm0KBQtLpYc0iKjgvqfmp6uGlh0I8TxDZ+wg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3392)
I/lBxmhMwgcpf9dOyw9oqFNcHltNvEEQc0d596VvUqoK+p/1y4UIw5cwUs5HCb+D
A2pgCBCfGR8g4Zcg7BlIa57sma1OYxMC6+CFqVql4FBdOeVUXt7sn+vediRB+1Iu
Jso35+DTfhdEFwfA21/Lia/VOrvgmY/uZ2XuDrnLqXN/FjoBpKSazo1hk456vvnR
ZqTYLLWNgg4y351fFwhZ6L6DKXgW8oWPv1zmJvMGifyysjuXcQHffYg3VVlfMFOy
Rxo1Z658uWo92UrXEeGsNfW+QzV/Ac6rIN/+LvFrWGyEGNH4aB5pHkQFr9yf1cwF
zEyPXDwDJgQGXikdXbFwD7Ye+rE9s8TM3JoUlEPTX6VMKV9pj3BWBCkCoLeZ1TW2
1ABFS7aXNZ3Av9RmvpGn/yTdZuJWaEELBvzJchz9yvGBqqKsxCN86V5rRT0oLHEB
ElVbx4UTKxu+4ENmHiMvspKuDvyKaXDC0Ov8jHsuPsMcKL37IpBskJtp7u8DpccK
MxgRXJhSiz7U+euGpJH16E8EXwi5C+5fKQWADDCTrnL97lZ1X2WePe4bX3HcHUjG
DYNEAfl/f01XGyrU+Quh+zMwjNmokycgy836NF5vZAuT1H7gx2qmVHgYdnoH3dk0
MiaOYfpMBLsIQ9sy3Dk7YDuIHdOFrJmonCnqWyYiytDVZiSyjrwvyUBbzbrcdtKn
hxinevRE6LbUCKoIF0xWUNnRf+0BkRsGGmxO+y8710DkD0SgDuYP4c+A4Io5voG3
lyPTI73+ir1CI9Ny1CyT3u4szpjRDw7ot6Wq/yNznU7VNFM+ZeiJjq1DJBfru3DC
dlgZ2GWhJ++4y/OugkBl4glZEVGs69kczaFjP1H/QsLkALWISEUDTQYei8/EkPty
UUFhgP80MroBYTl5UngWpBltF10JphAATtYuZgpFl0YiwC0nETfLIymvmqyMueMA
EwfUAYBFR2ji6Q1iClAFLweDQ9ZtnLgm3x3ZMq5IDB6EKtLnIU/eibFn9w/oWQYw
RovBxITuB86xQt1IFyhGKFF/FX2unBh02+Yhuu05WRMXwzuKDFiosdHglyhIzfka
3ON/AUe4heLcm6q/S04STmFH4SatWIaLRSknr4L+aZIb6AkURoOtLOAHeBWpyCAA
xYfLbKIOfQQKuDCz0N87Yq7B/9YhrtrIn3DYB/61O6tMj4QMP9+4MPeFIWpfSBGv
czVRapZWi2kcqw9e05uGsUa0cQohiy9v2Oqilj8UHPGAvRwMxOLXaMj3hhyPB9P4
RsNqhhJ9MqJ03DCYmXhbINZC/PGEBrnomXDh4sttaHrI8/kmf0uYiIUP5SQgczEk
24XNk9qgnyeyROWL6aUnKzUO4jQhmqiv59jqAzURXDBurgLAoEJN7+2sEocIF/e+
DxGVReFj8oiYh5IrUqMvzYjVTSXPlgoqi77WamLwdT7X4zpon9GOZDdkP2IHGUp6
Pu0rPBNpu85alQhtc2/phT6XhxOJziMHvOUF96UDcc6/YDXkVMIlRfOQhcNoCLWO
UL/I2BedTaRvhXMP9KnJtIME8HbTZofu79qt3xxDRcvuQr+Rg2NGXvizqff6taQf
Gn69RTMoyWnod+2B8ujxTmAKsUjlO4niJR5rSKU9bm0M817QchpgqznZWocAgpMl
98R+DYa102wOusrp3gWuG4vLTLrQpY80BPDZuiTHT5LNZsUoTL8C8XkHiwmpcWpv
6wpwsdRDMcE6Dk3bwaa7aAFF8MxH++RQPKKxdxH9XO/L3iW6F3SMPmuizrSjmpCL
Axqf/eNX2oqsO75LBPDNFbWnOgaDHdF6ilKu/2TfVw8KdihQX3GmnWFQmSauO7PE
RyEFzJ1/Jgm4ICw6ZHSTToqnlz6eaH/0U7EvvlmA59lbZE8eKrBQlkT/zaUK2dd1
qzppuS1VtFil3ZkwHZ3D8IW6MBQ4N8E346W76Euh97DKDXJf3fkjRtYJIkdxzIxx
iCBOoXspVV+nZD+DjohvaOVK/SfUzKUD8R9G8lv14egGAOPuWEpKyfXq3OHKlhVZ
I6r2jeXIEkBl+SBXRAFciIVBn62Ftzv0rlPhbcZUZV08uuWidD5lLop1im/zYW1k
LSm8VhV7sZx4WyN+Q7gHeD0xrEM7pDy3Odb9bnxhHP4n0iy6h8eOSGXDSIOjYp8h
4lbsiaNgK0fq6T5RLO41hhPXMNBvv98a1PVbeXpEfWh9z9f2HTwyXeDpOWRiUr0L
//YUY0RZSTOfdDhNIw4xjrKpXg+0CtxgKlDjJJw5GczmINaUoMhaidEr2BfO/YtJ
rUvftTzRhjB7II+rUp0zoyBlK6MSEz83t3pWmsEc3erIu/HFgnrBpXx7FdTwX6Sp
05mJn3CyazKrt2P6TO3dF4aXQhPNlApjYW4HQ8yCGFlyb1PZa0b+gtJnLKfZjM+w
3ADVW/He49JNzuYBj6oSy1zsgCi0fwhOBSKaKIkcHL8GBYZGIqww5icicneH3scw
Bt2J9Pg8rJP3WTESyUDtYVk4vl2zqanyKWsZovmRp/xh/cs8l3KypYa1zxVJfFQE
5OUFAX7hoqa536xNykrbO3vnOA0EUumXCwnQfEqMxbmeWMYXgi04AvoqqfaxFayn
IEGuG5u8mSGtJqlfqheuEIScbMhIjy8TzgFQlKf4HCNqOTBvebVS7arIBsux1A2a
XIEY9jAnmhawcQNTobE10lkdd2nuslAElwytLxS1WKxK5kcNPWPcITn2ttDuYwno
5LxEfFt/iE2Ev0/5u4uFx/ONPeW/xBvJY5SYwzs8AZYThII5ga8w85E0NS3xLb2p
xuKOllp3cE+/w2uftMOzIJNkwcbDHnMR+Rq++PhERB0koRra9hkBIPb9JdJmpE9V
0gEX0P+qFs8U6F2Xe90KJYgxD/r62jNUQfvyGfd1l6yAYlpyYLZFQ3/oArnx/2DL
eaHbZ3eoensnPRweTwg7zAap/onOi7mqHhDwSmRuKFR731zn7/ifIOnsdmw/ho5q
RbXSx5cSPYoG5wwLJb05XuqiGM6tzzeBEuGAdlz0Akx4otbiXPV5eApv3IbWP2hb
zQsZVj03nq8m1JawTalUNTdxr9C8sd9CpPsdnGHaJWKpZeZyAD9fMaXwt6cI8iUu
5S65+AR0dcglqvOzyXqOidqh+hQIgVn6kPWKbN0yf9gO0xTRy+xpOHK/MxMh+SnY
s32nQLRVakR0pc/2FXr41lg+hpzH40I9EtfmRMd5nwXKv1VLPZYTTuOM5mAN4S+Y
/R2hlRza2Ig1UUamNrFZXfFReSSIDzTDsVpvUxHCtBHs4nMVotZamxg+HCbNPpC0
dldEpTYcI5mOlaTwMqWcIL9iW6SVMkSCuzYio9K8vrbWuNloiIIqam+1WGeld4G/
kT5eYXLULoegHJovHDQRlTeRKfTQLDD4KeVaG0xW3qHLWrcEF482SKqHNyg42g0E
DIRO0kt/W6qkQomd93NaWAkQgMfaRxodU+EO1ZHD5VCNvJtHbhqVIrVQy/yyHagH
NHpBB9nzEaf8WRUruAbdPMm5Elo1O0EOI+oL0HAC99sKqLgDdtUSDLy/OiLWoe97
lR9ABdzckL9SijkXQ2PA2LpCmAYyfr2h9PiBlIoWsCJPRhkJwygLiN0RHABMhYOr
BdJqED5hzzka2ugIKiDgfYCPsHxCXi/SsAwZTGa6V8Htx2GWkIqNZ7ndJZtB3w5B
cuq+Pw8h7ay+F77jBubUYi6R+8buYWZMyxjS6qHR1SgcItyZktHGIq5ydJFZaVKt
ffOBo3NVpMdQXiYuOC/7tFDMA+BtwK366yPdDi8KYwSUgXdZt8RsY3l35vRj8fnY
PcDYJ/z5Wz6kKGqcZfOZTGXN+z9spca0kqKRD/LzQIwknkGDDMKJ7svji0XRwI5B
twOLlahvusIGc9wmUafv09Kt5rnsmKQ7myKHD8HVLdEhyAKs78+JnSrw/CRGHaml
GRCW65ldg3q+X1WOdorxMm3jFJIXevkNMRukonaCLTrXRJbtFKHxUqFkmPNoBwv5
lJC9XT0w0XUAhHFTStbt8OZy4GG+8ZFKSFl5Lj+wYivqPscPp8liIkPiYMCmhcu+
0IL5nNv9023CJ6oOlmRDgnMt27ylJzHgRD2LZUszjXDIcesH6YwrtL/c3ypG794c
fbma0/R7rCPTgDiSLyWatYagG558zxc+1nGkLVUpMg32mofv25h1VkC1jMTWfvNS
nn1HOzN0xUSSQ1BBM1vk9Brx1vBkrm9JS0UbHy9uLlJqAfd+Pv/2jQukC+X6YNVN
7CkH8uzeYdshrmzQmZYMeE8zP/yzGg40FZHFh6XxBS2BKbY221XxsPkYGYQxtxiV
eNOx7Te72Zzx+Lw/tcaEUcXpK600xT8A8BO1Xynh1nHou8ek8HtmdKh/ayFycZvp
wLA7C8DijZtNf4tSvNQv3UXfFNtAIe83NbQETmgq14DJ01q03NBg8XDC9kePwzAl
DAs1EaKFHlvSyu5vefLB9MYzBPuQ50/+Cpsnn6COQNM=
`pragma protect end_protected
