`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eWRrUuzm6fUTpSVtFJ1WZgraP1Fi/pJblB0UTVscRhcG9np1y5p4pGSp+0TUIOgH
BLnNtexmXN5XlcmDV7xXtDQkP6HP+PvFB3VLEYHGZcmbK03U6XO1NHdG/ab6yO7q
S031ErvGWJgNbXtOrRYkhbfvCI3MkHj4TgpCqax6tZU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6368)
xXEsBqGTVmc9BWuEwIvFwMrfhmWTR9E2iGM94IElOnuK8k6GLHA8J0tnVEuXf65Z
A9y9XdnOmdbqIVqER+6RUDXEptcyhvQa++sktRyUp5e/k++pFEWUKFl8bj8Xju3C
T0g41Oarv6qTs+tEvJctSnkzR2XaYwVfDUqAtJ1j718O+Qh6NMmcC0AOjduVGbAq
z0OjxemdXEUO//j9mqelJohFM8na2ARQr1158X1SEFH2L172VxikHJQLvPg13irX
DAniE44pfqk+fpxLQHFXJcMnn4LnCQhOCb9mn+LCtuEW33lTH13Z9cJMN64ojQWi
i62Vlytd5dCDJrJPoEhFceGNF1cITa/8wJs9LvX7zmXv2kMMv/qmmvQWYOE9MVhj
VOyTp3xde6zPDFg4UqPyqyGlk8Ua2ux265EiESGyInDk01HK7TvK1FFXSlbvJ7Ka
TfS7zOQ41y1MNWbTqTbJvSqKEs2UQDbzmtSNJ/7ZX33Ka3/1yu17g6BZvVeAftSQ
4S9TNHBQXaRspEl4/aA2gVH5YTqlMvsXAt8ItIlZPMtIFSB5ISSpq6ExN/p4zBqd
XstU3zPLc7P4d279WBKmXL+TwX06cI0id0R7V8UDGNfv9RYZHiPjlNPB8AUj3o6k
0IJVQmc1jyOkwxPgB+tV9THoUmbHGNOdTV3sIMeYSXCwGgA0NJ6gcZeR7Gnz+P4b
wIf3Lyh4XwvywAFdOTgTfIDp96sIJZ7mzyQAWfKolg2f3ltPLnPGmNEYxaJErPhV
SBkOM3fx2MN8n9D5FvYMGphNXBAxD6XVat1mWPuoaUhiPrFtx2dWoYZ0Ef8FVbqD
kHD5/QIEhs8mMKLmgu67H9Cnm9HhlxDjVMJIV/AmTZiqLlQqrOfh+q1q5kGyJIim
Fx4DOQyNalTSX3RDhYXa7PnxLorh+1e1zvTNgKInaU0ELJeEQMQSvrVfr1lhwzRq
ok8AYxhJDNlv/uknXjCYB2EXCljGsdZ0sf0IOc7BQFNN43R9f5pDJW6zgxGutfZ3
VERjPive9p8NqQJPR9gK9Fnw6a//FL2DcE/ugWeiRwMi+fK67PEziJZMEIiYxw9W
m9j9qHmNHnVP6gdg+vLHsct9cIhZZd5MSXoDNq7JVLMEs0T0DBnUzBB23J7g3M37
OfxrpmZocsYZR05kNpLC6EeJcemajDXA/aRyrXb96rBl7+NLTanLrHCMvt7uQ0zw
vEX4RgaEGa87etds3/M81rG3TW5/PK0OTgjRrw+x9T9YVDVc7Pwg/U6rh4GydyGb
dW3a1ergDZKA4BvkWKeif/pdcPzGvPC+6TUeb/AdlGMfoE2E2gLtWWL29Qk8R/lw
TtStVgyZPbBmPHm87NTbc5/5I+JwheZQ/pTOH5SnuV/YEP0Z2MRDMp0C2pqFkj6a
fvkfmanznPB0rfMzA/Mq4MVAp2llTPmqgLpic9TeQ4nKOiaP/+0BFta4r49L6wH+
xl658oKPfKTXzsBIViRGxanp3kx7G/7YY/2qGCCZJu3s+2fzqVcXhIjjRCpoYKZ+
x8+ojSHdBGygWyEjvxxrNW5SNnkcdV/IwaozYUwPAUqFgL3j4hpV5RI/Lfgch2NO
CrPIhdxkeeDYBqABG9OJDmPgGLSVeZ3teot8DxSGFW1maD02mxtm7KjJm2/gIuEp
hu/TrodisVDHase/qnEVtvlkX/8NcBcDhxm/oJakhCF5MkUgB6dwvmIt8uK/9YH7
Klm6/P9JWGJGvdvRPtEf5zSzhMHVcRFQHYk20s1U7SgatiaKRHF6F6fRmNGZvS9D
uBosQB0Dz6BoIYf8BpCJEPcHliz/Ld+wmnR7CjiRF0v7OdFgFhkMRZiyfDDmLCIf
Obufr4Ismaq3vzFcaYKd8fbw7OxEKle6DskBybVe+mN0JnUTTAIPi7JCTvejTE6c
ugk36fHULahhlzQL4QdaJytLmIqmw4akmt1Np7Y5/fswL2Kki3NZwkTFP2XRazXa
iyOjmLRHRbsHb3muHAI1M4SR1Xtk4Xosqt8M7kkadPuxss8iVv7g0EG//+ixoFQM
m9uyn3gxCCjR1oJzkNbQrC75IpKMM1VUF29F6wrCAqlM821lL+1n8T2mChTd5U3C
wbYHO0wEkdGCxom6PwYleqkJuTW0iwexmOju86NmFIzW9RmrAi3GyG2Uig5aheE0
BjigaSCBT/xunTLHBq5NdgvbKGYn+zehP0R6DkfJPPbld9LtWYXD3ESjjqql53oc
i2bB2ekS0WXSLtnc3QNSvC/sqznViTQLOcZPnp+SWkyYJWaSr1ElJpVzqrJYvdXD
VFiRXTkqep2gFe4AswUR4SlE5vNfN94K4gAmW8AjqTkX4Ad04hSXj+zbZRg5jQaB
e3QiKZiDUJQQEhfZ1MLaLG7HPY4A4wwuAHACWxs27BJRa2VN4uq9I2j5WtfGFcr/
FOR5oIYTplfaH6F53K83kUeIJHtFX+Go+KWQ4vPNCrDk//Dt3L6lDorN4ohj0CkB
HZMAuBJk1uJtj/W9qqCEaNZnRyTGSf6+yKxwJeQx/e7e2jLK37uAa0OvZT8J74G9
GgsJkjK0CY0pkgWjeVmJCpu5amAt2/t6RIp0Nln5dTIjJJaKabvHJH/XQ683rv/l
taFjFOl8tkfNPRI+zkGVQEgg+dk4MLn9XsW+sMCesf/etYIexFUUDDAeD+3x1kY4
y0A/nG5RljxKxNi0TSgU0U5mWjOadaFxxRV576qo9c/20vqt1aeM9+xz74k4j/wk
eC8z8GhRfLrQvpTP5L5UF3PNc5BisoarnhqrkILIFZ9TeRkeOWgZV8Z2b90uebtw
zo/9tpRIAZye++jGxwLZJzbzWdEZtZKGpU9NLHesSjw6LgpHqpL20jhiKFUqYcGA
Hb3gCUst6hTE49l5RHdhPVdwtgVFKx7INL3+V3DBkb7D8A3Mn4ytwXvTTooerb52
++Maep5HAUUk1ueqP4tEbBQx6wcrnFtQpeuXYt0JdqlRRsHTV89h4f/2ZWjiH63I
4OQAfL4pMuh462XWroHFdD/EyXx0GgssuyJbYNfT8v9uEDoyqhIU8BXRR6q6HdT3
rUcBwb2YJz/e072c/G23JIYpXdLiNNNmeZxnmFNuhqcWc8qD/QH5zukN2atkWaW7
f6V0cR3daaS0ImA1jzPMOj8pkRv1bUUu9zkrDx1ILjjxY1WaZBP/HGxh/TF/HnrN
ZTnzx/WLLWH+VyEOzA4DMq/+YYK3j66O3LdVlCHvNyi558k8Kedn7BgbMgIvsfpn
ZxnlPJr8aHhvxWYCkh0IY5he/mHt5EuVq+uryou5rQrijr3S8t1UDoBcmwsHT5en
7c3O0UhaHqsl3iUF83XyZ2NMDosM7zaoD+pGOusypS+4v0bouAd6YZ/PG+LXarLI
iLDn7M+OEgSa2NNn7ju3LyyzGDcBb5U6ohhbmcLfOz3nZ1h9tSfE488vdPKxeWzi
nlq7ezXg/ANck7pt4rGVJpSOaJ9HY3Zw9F1Co2MCHhBAWfi2u0xq/JSMp6Xznz32
YsVs7gg5CiZviyQTLXpfSMhcFptCGOB+2rj1TIeWpKD3AJJNKl3Gx+DMvGhxx1Ni
17/iqzg/P41Add9s3RJt8stgmXr4tTQNPVtkcB9UIOjz5SVa6L1845js9ingTuyT
1QFYjgx75edLrrZIHVXICxVcVFWGXHAw+jqksomR76RUV8qsphP1UYJi7ofsxaQ6
Sg57akwIJWPALH+674l5XYv70I5E+eRKP4496obdt1v/u6nz06t1XKrvDkMfbHIc
b94pBk8mLn8ed6uTKJx2XBd+DJcdOvurQ4HR7qMEtr3d6zMOrNSClVPhHR7vS8ny
23zV9eY420S1ZCei+n8wNlgC1ueHmWB4djF6sdnNOujN9tXj25Tb3yttmYWFG0po
kOdDmS1fE2oSQQJtPFszHxCxOq3UNY41K3eLrEfDTy2bWR5lYJCwqTFIayu2iqTG
0HLXYAzwnez/1YW1nEBFSNRn6EXBrpfQ+/kRzHhdk0kZhHPiQJYA6l+b36GMqgzr
tUEgzQq0hP3L1M+PJp3d4uY1lclDcKv8i6OdwcnqjhnZgWDxXYNnzeCFMoFfEh3u
tZCU6fTc9tvVYE0Cmbemp3313CpELw/JBvvryMoycXlIVfrro+NnQ9QlDYvy2rV5
HG5vKsTjTIMiRVBq/J03F6IbTR6B5Pj9++E5kZ41ftJVI9TnchXUKKwXLsdLUvn4
90yaRosJaChNrTbgvPbdZwaQT3GBulugxEP9fB6aYlZjCRojTdWiQfTlgkXlhIv1
FsLo7uLiv3JDjOHTr2yrjGFFL5dSM4R1sVvvrk9AmyJjL2srOOBmS10lq6BZCkc5
w/qpi7eZ20s8Fe0pPgbYfMioWIhdQJi16zxY4fVazzSZ27qys8hu2l+67kIsDs67
grCPfial7qZgOL2sSVkxP8ze11by53C7vJrUhJRIgGQld6YJXv6FxSnezgfv0yZB
B/cSKlx/QbFcFDJTaAEzAlrgPYLCZF1z05Oa9+iHW7ml50Rrge764Jj9dBXwY92N
AlJxSU8OrKYIgLt/ojlhqBeepHO2mPxuPFXRyUK3OL/VqDrAxHhHu8HWMqoJs4K5
ERPxCObL7j3zz20nvu8HJ7hFlB4voVpyDHWhAcM4MWaIks+KsTMUWZ2km40e/Lbu
8TSjTQ7qc0EJWdlje42Moztt4iy952UHKG7l/mgG/sbt20/uF7xMTnurkCvYfvYT
mm5Pj0jtYQm5vy02cam3mOVh43ZhVPBh8LXyLMwmzk2GPVbU8x8UyayibF5cmhJq
uioFiRCnJxhSTh5RaXLyC9R16Mg6R3CrWT5zX3/aQspLsVlP97vJLXZ9UsF+m42i
c6PbUXdrbsXPDaC0KSpzkpjijKp2yl2LHbqzd0OJY0QPvmDyQMpsMWnWmnTDNBTg
3JGIiQ90uAeMBKavi4Z3Oh9afRHN4cO8pHFdpsEoJaLuaa8qUBseoj2wGNEqGojX
oJOJZZOypyqikuI47nsVrQxZmTgi18/diDWnojfPkLoUaabZ4JZbQ05jklhUMCTc
6hpQ9Wwnqa52c3FRUv+bmMfG0l+b2xZzJ+uJVKOrXO+HUWipsU6wVThvkPDw2zkU
jlELSPEn/y/GnaikgRwq0IuvRwJ7f9pAcittP/tSlrXDFHiDglUFM7lIhEfa4Rrd
ob19slM0UEU0T6v/Jud6I4tWFTuiiTiDrGBGcGkfBHULu7H4UUg4brTzspjsoMDA
DOqKseau+YRCpNNJWM/DvDwJN0eN4Rrs/81uTkjpHOKRd9Nd5r2sh4ytNerJJ4U5
OQC1BEdldwDyxwGZhQWGB0XJXafXgB7Pslzua/t4KZhLlsBBJe5OHCp+R+HZO83g
zXRpD6mBYD+ic7T+C4ZyZWVZAJYUluW6uUP+M9+Jr7+QJhd8sKnX4YhwyaCRgV7P
S/zT4Y+nrvzci78YIK/Opv/eZ6rckpm751fLj52fN/bjTgGvBsUt1e+tK2jVNMO9
hsMvyyBvSRhAl8TxVVM6YmdlgTPcBBspcJm7fq2RccDD2QHyTN9T6sLNPeFsY16H
qKu35MOQwhUk/oIiaVUu9KTgqPUTMXlo16U8m0Fx42uuwPIOW0foAsLB7mQjb6Kc
Rn6W+yposTY2DXmcjizky+qy7YbrG+PZxeZTNbARDJzYuBRiAurtxMpv72kSJxDU
ul4k+E1hAhv9/dEbJKWbWYaSVpRjZEZiVsVBVG7/I2gtzlpVIOoGiOvx7RgDGYZa
SSBahDOnIMRZmFOEqIwes8nap7RSUoctH6clCSQMA+qqtIMTWkxxz9UTT4VFNFaK
4yCtniUrXjLnz0HXxEk0TJfV4arS/xZaoIdjtje83iTPouvS39Nn2uLZNbTTtOHn
uOOqDEX8ESx8joZfqYehqgm7BNvWZXLfLs+5NMlv2lHFdw4+7QmZ5sa4xl/kZDd/
OObb40hAbifDFKaPzRwvMJ0LEyGVAy/5eUguRE4S+Xr6R3vxEJbf4uURd76vwgAx
KiDGsL4RmIZTYHcgoQ9JDoenyIc7lPtlnKPcIb4nspTo5gU52BguoyDKOQhkEOiL
aivXorSGj2B4HJVV8+mv+D6jNlajiETTvSAPaV5yWcBjhI4IzjIW5uzn85FYf26H
CYtZ19QUPoWCIi6Vwjh5fp3q1UpruNggFh2zxru5AAziuc7tC4DjflfElffmfRc8
VVlpG77SrnGIUDq/+u5ctlQMbMkKQgluH3b+jcrUhUn9J6CGpuLHvYbfRCh5ns5E
HACz9LqxesLme0JfcPN7Eh0N73PLIgRdxq0mQ3up9XQ4dz+8Twfj7kiJ/yd3kO35
Ecdd+Le6UUY8/mLmM6PtUTHbcWJgZWFuXaOvme/ecb7JtvD2+cCq09rSeY86X4ap
0OONXVktxYYMXPhzSxuwtp1L1RdZdShOU2ytyDbW2Q/7p82PYKrLNo6fsSEGM8oE
mSeD62yxsW+B3thSC2Ve/iQ7nOrjgd0kqiADDP+xMCcM/ilZk378rN7yPAE1ogDY
03hVUVbLe7ZlL26ZNAwElggFzy9z236a4ioFUHrJ0529lmfeAFaV1eD35erz9w2v
bKBG1Hc6tqUQHLcV3ms3fsQqyz+Z7Hr3fo09yp1QIN6RfvIr/BzcrDxpmCmZ6wtq
ueTUtc7I1pYT/OD+U/8ubpdXagcqPLkliCDCr4jwPS/gjOYEuNgvpyAO/jmDmBcR
Rz6FDwtSJkhIOeFa4/KDL2OZfQqQxU4pXxEUYeedv271VsXzHFGf7zUW1e1e/O5F
uvfYb9vaDJTZnOu3XkizOUofZxgGG3Cj++b9u7uvJ+Kw0nx+uMo1Q8sYxvCl1G3C
Xu/GnjKWH5ZcXA3LRw/16+fNO0LRxL+MP/M4HAJkUg+iyL1WT+gKcwGLTNJZy4AJ
KXPGalGLyp4nxcsKT+PoVIe1/DKWO2eAduKuAmJnElrAWe7IscWmNuXmA4Qv3NtY
eLJ3v1VmQ4QFhgO1QZtdyvzJ0DczbtVU/J1FBbACpmqs8nNFAvPTtiDS4/CPNpVA
glK1FnWZNrBRw3xice8/NyszwBKHBNWnYL9W1BOIECUubpKR8/NyMWLkDjszQsz3
6jcoP0XczUZlRiXxqFFROs5cqdLReXeuhgqLX257OoqGMkroDc93EFJS7UIap2Cz
ebkuTmDk8XpVEcmoz2s4wbv9pvpug5c7w+E3Yol4XiD0wcsssq3RrThHR9nEUXR0
UMTkrlLQ1oTdPhqAgGtXqdcnlNWaCr4J+ovET2NCSFwEgeFLNmsQ2u4YdUqkqhaj
43ohSbZ1lpRod5S+wShgmL/5GyG7H1gvwHrfEUFfKkikWw8fhZzFNQE0j3SZ1FgU
5n97BcobO8UUXcc4GRcj0dqQ1VdsFDhqovpnS0n1zmQrR8rcf6GPyRXozCMkxdXJ
Ftl8bkqz4EmRwO7h2NDkU+R8wx/lkuEo9azn/dQnoEKbs948VaXOBA9ev657SZr3
YaClPZYcmfNc6HDbp38jql9dDCFKSndI3aj2Jtinb6EnndOzvXx4l9aRWEZApknz
O5m4YQp6fK8+/kjJK1HYt+aY0QHWZchs/rflCl0dNugARYSikI+GesnffZRAbJ4f
nhwFYRcWP+Fs9/lehEUHlTGwJ9rkHilU8PHCCaVZyathB7o9Rea34MjtT6nW7XhO
d3yViJT9uthhW9yu3RO5OgrBuuQT6K2M4IfKLicuxiw1melulslo41E27L2zxrMS
SlWrmfIDN8UoEF9RrMRuV46se7DNnozzeCaosnvHu5LjUEwZohjkGa1TbGRCd6+Y
3SM+3MHNlsYNveF7W7v5lh/PbBVB1YeqQ7uN50f/tDz3/kN1n7Zu5awjHe1LXzQj
BEI0CsgKy4CHaMGvAlNkD9G58tX9Shg+IhIzH1AOm+DmtdJSuWoutj5d/h1lG0ie
grCLiY9DN/jCX2NSZdMfCxdPV08BY2LwZuVo12kyYFU95vR57o9Fl+FahvgyW+mr
X2FJ6PWIBP/1EK3Q4SAcrocZHfGmIoGXk2+OF1bFWamvcNpMaBRy0uR5raqHPWpv
pn/evtoA52iNl3GX62FY0X6FBPOTSy7sXVlw2UQmXm+GfXu6EJPNlBeJ0qyPruMW
YxN0PTyLTyTkJpvLgNS3nazFtuyuwxztZY+yS0SF+W7EaehIZG89yUNyQRl3pFhM
IzbZPwXHBo8piP5gaeIBaS6xzAL1mtwgc4WkZDWTawbYNDucZqQQt4vQsj0ikJ2j
xsWtIhicJOlks3TqKZdD4VHmtZByA3m1Sl7OujP2uCJbcQSqCEv2MY5ErO64gPo+
I6h2n+LygUpobEeHkqF1OZwt/JaF/xhkuSbCA37pvG6Ixalvg2hUJ6lPRiLTrtu0
jmIxFEoKRJTBnsrDGlwAPazGkr4hY6o1sjrdVcpssxn8x+BYbTC/5iBa69dscQls
nFUFU9cKrl/fX5Xxd3hCMBGc91xA7XbHX8yxb5q24gM=
`pragma protect end_protected
