// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
M3dhJvGvEpha2gTYwjoX7R8tdish0lIeO19w2lTpTKL67E8jEITA/dPU1CJCGnRdWPXiPxGs/BdC
zbKjd61rZX8/kiyi60wbDvFelcuik5cEPHceDNebwNcHIC0mwf57LiIDimiAxgrZfTIGBkrFH57g
/9m1Tlv0XWkY/GUIv3AAM5N6zqLWDhfapivxNOAfTLRPLpR8FvZ1vg4NyEQwWyPbWu8wGn8w29Ac
PZte4mKVEhdGOU1Dul7ml5hk+3wAB6KfURx1LidREIsdz/2ouCwvr9TLBZWcW2DnCvKnTmiSAcF6
H8HywXuEtBd3ueQEoVMJ0LqXukIi+760VUy6Nw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6704)
b4ycHV4VbZTqJImv0YymToDn1Us3SlJ8YP/790f0H2pMqxM1b4cj5tfA46EKiYAWXzq5d5QAX8Pg
6ef3hj9/ZdkMoX2EkTY89VdhkSYsh2qx9+UCnV0Jcz2W8PnFWerR80xXLbgfVbTF7rx4dQNa4uLm
JPh71rh8tgWHVoslB8/RYQaeAnPuq9zDlE23FH9t4J8D8/RnjEQFrVZT9R2cZuW/E2wfWVyfU/tI
JY490gJgRE+0C2x+RGVFTRGHe7HQMyofQHNH65QbrGe/1Ex8iZE+mFFGztc8M+g8ZpJhN84wxV3h
HXu0zXscBZFgkUVHn5HtJCQpS7reJRtAhCeZEo/Rnzi506gpKsC95ltziTU/rz/8sMXNpw3bph7u
7GhDGGCki5MgYkPm6a0nWhhylhG+Ic45ghfH9sUVsalyuQtuclEgsfflChqYsvFY++w57On5VK8p
4Jylm2we/tSSJNgev7EPtAHb7lIJikjfIC8fpEqbND+60mk9kOZUJPdU5N66zovrn7fXjXSaYFfr
Gv3Chkp1veuUsUFU2sQwP/GM96Df/gh7LWYT2HPsTFZ7Ba4u47jMUXIdkb4V6pTHM/pXcu7htwoR
0UYyB+VzclG+zAGQVbErZVC9KJmOPFPvrrARj89WD8AUpFLIDWIGJpLZhRVB7m6tLGKrBrOc0KXZ
ixIWH1ZzrBkWyXceOSWzOouMnctDy8lWGIfQF432C+5WOxWI5Nib86GIFe06MmxoPSfxup9IfBuE
UlO1twTlJIQ+iWrCY01hczQ8Pr1uNsO9OgA99WbZYByiUUr4dLxLaoA3jRn3iA/tUrcYd02X/577
W9/bldF6SSOqTgi8F+EFkL4QJ6frlM5mdea+d6zfcMwFkpfHsbvT/lPPRtEg5J0LNh3q84cuMgig
fRzF62NuR8s3aOkDLLFgVAaDyKbSrPwW2uvkfMkNtHmR499vX9OruocXvo2iz6NaIi7XrVA1C12C
InWfjfG98zkaJde02wi/kHdOIhKPnj+EmCNgzIyF0IkQPRXKcFrHBcf/RBrEpJtUfqKzMG8klauc
9gRp2ZUjq7G99ab4xleZbU/b/DvJ1nYc8kCOgxhCzAs5VvUVtB9Ijh1ujgg8uPOCVhGOrU4DIlxo
3qNUJdw390BQYnLdqESrTmlji+FSt3osmBxi3lpbk5cdXBWlA6B4XkZZWVsiXctiDBPkc6ZBAjrL
APpijQl9oIFclUEthZwaZ1i/UYP0j2lGblr3NAV09sDzJODz8cxpCiTJs6xlfD4X3pcq4bcM5LQr
LddstoXJOGEWxtJ10/OYBCkWqWljx4MhPV7x0AMH+xKsJJy647xRZKVXZEyKYyQaH6xlplCpBVtS
Loy6R86rAgcInGYiv3uZJVB2nlgZBxKEwKU9W6zguET2oja66iLVD4bH3Fh2OmWg1vP281aZ8Umn
Mxhog+LSRPDERZfHhsmc0jM1cdr2j6yRaPFl9nUORkYCkhaW/qfwrq8E4gvjKKsdho9o+SW/UOIf
dwl79O1bAr/TB540pwGW5xQlQWXH1fqGUByoHoJ5UzWr/zHsVQmoa2VL1/NCypCFwJdPRHu5fgQ6
A4QmFzgope4tCb+uCk97DIX1z4nsUEB/F/lKU+zHBq7Jrh0ywYWrwiPonZIm95iN621kcojx18rl
Yutq79z+8bHnHE5ZeQ/IPZFJzprxzhfOxljs7VHPZHxPl4/eK0Vw2XF8QVGSxYHGGBWJsd5Ql8Jm
cilhrxcZxun7jeOny1IP4DhaARxVFSDn6O8RGu1WXbmOOtK0lS5QbaUpjGcbCayAYgTASwa/2hN4
q1slqGkdJzZaChpXSMId8o9QK2yak45Bh0Tg7DtEavCb+zW39X4tCMHeJQOYqIz8PZcnluJuldm7
erTS1KvhkKPDeViRW8p53PJ/K9X/gpuRMS+GSiSPsErxm8TPrJUWPPh6sV4ioVGnFO26gPVqS1Pe
JIWgs2sq5+VFwvftKoY2xphqLQcuBEm06twYl9H6AV9pcuPo1sTO7BjhDlJNMLDrzifu6ejZtiJZ
f+a/gcY4FK7Yx4iDHZ4NQemjoWnwPM8mUlJaBdE6XODCh6WXJc6SPRtWN7wwnFKoNKAM9G9N3XLQ
GR7vC0N4SpLJZ3x+dsTH0l2KMTSarN15kuIczIzzhACWXaM/JlzLXzsZKe1tW6KcdH5ibnxeyscQ
9vRw2N39OBR7GYBqlJRXnUAVGu6FfnXVvFZYvcxsIIoZKlOwKC+1G8QEkERrJes04RHsj/HGpXrS
Ff9GZwzkB0fhmsDlrR6bqeFRMBKMTs09CBo4mqAwWNqnp3wT77dM/Cml0Eq3b844enQPquCqS7vX
oasdsODweRwTm/pAvXvN3lLLWYj3B9AefJna9WVYWur7vHKUs1uwoYB1GkHc0NN1NV42wR9WcKsI
+PlfQhKCbIRTMJhYMR23UNoVD8FTs9+NtngrjwSdIOGM9236Qygw4ZRKVWGRHQ8/qEwpwjriSa/Y
1WWX+NBJZDdN4f9GL9oL9Hp9fua1Vtw9KAw1Sgw3P5hDmrSWMxNOg3jHfT8r3H7Rb8PAxQo8braC
ZqmlGdlO1BOubnkQJasE92PMkPK9xUfV4lmurAWhv1ZKty1W73pc1wrRKinw5zfOUWGZTd1f/IFJ
NOL58ERUZ7NGpV/ulC4kBAZhG1IOhLoOW+Xa7rhZR7iNJ6D17Is3LkfYYAHt71IE01Sl1qXvB/1y
qaTdwHYwfQz+TSQuoxsw5JAIqNcfVlw4K1EDy2qadn+bA4v9Bd7cZyTK3x0DUZv0MxUY14IakPW/
8YAL2KBAf+KgZ1okC6B29x9+JnF8suTdcAJotxYez6H63MekPVAMM/4RdF+JWivyZ7wAL7Idvad6
rb/Ndga0vbyQkIUEsbEy0lrKgpHVAxz33WgK2tjZLqxHJSnnVmbF6b9bzr1Xro1IoAkwTacWgvdE
HhnHD+ADxUUlnqlBwUL6bQtPIF4w9gjhIgbPUI8kBKjg8SKNt7/vMK/pIL7rh3LR4IewH3ZQpkWq
pJpKxRQMyeDCj0DA4LGLQLqBrYlT/3niDYUZLuZsehoV1NCYfT/tyaU7eIXvgARW+7s3QtLuFlCg
6Rc/WgohkNWk8p+PXrTkAewteektBP8mEudjX7Vl5Xx3GECEzlDV6Oqdm/6BqpW4I2Ne9Ou9Onxq
F+U+t826YYyezb/eRh8JaxYxYpX3ug3/FFHq/UfEH3bTLShcpSSWJK1+PsNq6qcg/lOW0Dt+w6Jj
OnQiTpVAXSDCMxv7KaAhfI4XT2T2Emq+tiVwcyUNK/2ZPs49Af5+CGFrF3QP1jpmreuqPF3VNIZv
icxwsOP06b59Y8ewQ77EzNqDZHShQn3QknvN0AWYHo5KmCnt4ktwGlJAKzQ0GWP1gJ00nU8eoOIB
IlQgc4PHcQzwCLb+jYPWCd3sC6djswoZb7+DzGgf9Byll8OC/0CIEfUep58tUYMNuVxals7B3xEG
SslzM/rpdJyHGesXgTwrEs+zYOywVBj73dVMi/h00riiE/TRamck0+qJQYJ7BMYVId6tpmFULCFF
O7UGv43PemBGZA7Znn1fFjrICdS40et2TeL2ft1VRhpa5sf33fPWHk/RnK7sHGFi/91qX9Hm1DND
1/9u9ID0VKzKhMt3PaIIBDlpi7q+ZnIT1aW5V1E9ITJ6UbhIDpUeZjgBMEmuX/h4asiqCm9D3QMa
kwam/+fad1Cj/6huLjs1NVL4rQglKuSf21+gf08p3Bu/Sntc6DgfoHU1sa/Z1B+ODEHnz4kwSZiy
BVKs35ZWK9Ccq3jT8l49HJGDBZ/j1j8fqjh8Bs/wQXy8Q/mX7wIf/lNf6ObHc0d1kJh9GwG32/nv
y+C7NahI6qsj58GbzE79NMCWOe+ZcoL/3dkNSoNgePa5WsL2pMNfyUaZq9SmxdbG4qKKxmUyP7bQ
IeqmAo46BY1QLiRWxfFMNT6GkipvPG7Nm0//2ZbB8+nfaFHecRjyfTReGVhJ1RBdTodLJYDJipqC
WVL5lQloxK8iIELFRYx3BnFS8CiCc3bdQGuq2ipvfBQY12VhWVggQHy9rn6+h6l4hmBfTukTP1t6
0ClRRlGKOhTm5M786ccyYhKEELJiw9WgqUB1w2hr5Do8R7/dw/piEjCVsP6e9hpxpelbl6sK7XGB
6PuVCC7iCYlWj2ItNFOnUr9d2S4pCyy8HVMiW6eGZG9IsLfs6o8JOvlLsdtrgnT2y6u+U6dBm4d0
hfRY63lC1UJwv5nQU+vL2Z28q3MwvTSFR8cKrC/C8FT6AqX9UOywj+xUi0fbSdAXqfbNQ7EAmhq7
5Mt0ADx2mTlpHZzs9V9gjw9wP29A3kqXUyWP6eEv6rXw6sr/GQfTd+AFyJ+Cju1aT4nheUc4g8OL
9dCyTbKZ/JhO7MC5zdaV+dpuznNTVk5z0aqffiIOsIkuR/WGkP3T5DCMcJ1v2NQdiitdfUL51dbj
9xErmXXCDGdjElLHgc8CQQl8Y0xbPRMaZma0jCuWRwfpLFwsnxgqiy71sbqqdQ7eCE9Ay72/ayMG
AgQDZE3rYx5BCaWCnJKWYKFH0wvVmM5e3uG80bCxe1pw2yyZ7n2Ysgyx33WLxBfwv0gWD9oIXZRy
ZkeU+BV70rOMaO0ru3hBn4MPAa5sfAQpV3RRX6shztr0NjhDoMESJ07LpvK053Liuz0rI8j7ykAc
0Z+2XzRWCe1eN3XaGpAOpw0shIPsjNL1mnWQ88EvV+PMQ6uKxSQn582V9+CKo/KJdmyDl7KjuFQM
Qg+yxEjzR7Ja5n4Qjyf+Id5yJz9MCL7yjeqi9oDe9Fh6bzXUlW/Za7Ks7lrZHbGgyc5xOBpUYkDL
ILc+PrGzgUsgvHEWiM5oWd9seSUYf/k6sqEL4WjqImL4E+C6xwyA5DBf+pvYVb1QBps/3e9WVdYR
A8l0tW6biQuDxaCGXXbT9kMtycV59bvCHbxauM7YePzdMtjysdN++TUkFitOMS3patXKbD8TlpHq
i+nmIAWix/ngY5jd7MiMLh8UO3rHdP+cV5C8OutGBHRtLXnseaDt7puU1mg4xVEJE5JN7nh7cLKi
krWl4i/ADExmugJexhx5/fJkJoNZjvYeIqABf9lpau78pq3O9ZEC7tmunMHmal68+AmAgo8+IO27
oA7ksK94KdLzW9me5qxVGRKmaIe2rmVmawZt2WtuntSoHyP5eqKBZDqEp/jAI2lf48gntAGtdPwi
TG8eMv7+4c0jrxuk9raOA8WSgPOR72EhvZo3FR6l9f6lHwwB2gf6r8XRIXTAJPnukRsmJYj2H5g9
bWgSbthQ6XmINvanEx571tOILb3+K9R7N2ibwQiKWU75Z+Kz4f82dsqgh4XSsWg30wxfYj4/jlbH
gDs3eBCDouQfAtgYAoqF3x2v6xkP0eCUgWJAa3E2PxFI3SvAV7krETZZIMaaIQhEX7pKxU9vP+7Q
VBp4kF5fFm8t4F7EiUxcb3C/8HWLUPGCVU30BEpJK1D0VqihJr2tuOCFitfnNsC21NXkpXWHNbN7
q1+1fxUWyPAheCh7RiGtIY4sEiC0JNlNoYvIrq8iqbmjBxMiqlroHCmy4/oNW4PKqtmWhSP/orcg
twdnuZK5WX7ssaa+DK7b1lZe3MSX1f6aNex56KjbD5D2tFzEt3RntYQr5JqZEli+3nzSmRonXpRw
Mh19X8P/WowxqWP1W+YQ67X7morlST77V4SmiV6mLd19WffCU61H7Imnw8mweJsUcGxq3IMtC6h+
hYr1zXdVSEdvQGE23cxhCuuPPh/4kz2d4N4R8XybJE15hyRxSOk5VtWAMjF0/OJN9KIxT0e6IiUx
yZINf0prUsZg3Fy2o7jNGvgt41M3oaDvW+NjJR6W+3Bis3QHkAjJTYqJArsqAu3D9ItIm8ZbTh3y
FKLk1qHDCWL16ZFfNpUpT4qE3FaEt7sE5YGyuLulSJqqIcQq/3alYb24MU3bxVefVVA/szjZnj0V
SSuoUL/VtQ0+pxQiDwAG6+R8XB7e6dx/VAIchSBOc7o6EmjiSvOzw3Mp+3/yYszB1n5bpJVlPVau
WkhzlpMaMebyJeUeZOhNuupBNkgB0ZSIoqaZJEqqQvQlB0r2/7IEWieF7eZjomOmyKO+S+frW710
jnY59k72gJhriet05nPlz0tPxa6tKVpb3Z1MbpuZ58MpZy0IJfUZIZr2LKOui25DY+Z9c8stnvok
MEFeMi7gXLOcEyYjIoGZGlZ+Whhh1qC/HVxlTUT7YZYL9hWxFUYh0H5r6ijc0JTHzGYOIv7g7MQy
0a3D8qFEQKtfTeRpEeIyPS8KzmJMoaswGkk3E4rxDtOwgf5ozZ3l32Of8nL9D7+7zCP/FbKA7Z2A
5aYPMkuXObZnaajF6mTgPIahL60rN8pMKAbY7dH++DQThq2e0tuzLgyUIcEjVimwliBxt4rtn6tk
tVHogZS1qYTtO7McIqnRGMBQwCGWg8nq6t0a+Gur/uOGBqAJjJjuKTMIBziJ1ssAaxK8BodhJcv+
zXwTYarM0H2hc47LFO74ANZZ1PQT0T4JCpHAwnconCohsYvJKTcBwSX4kJqZFHJ5+29S6lFuVpjp
AulTiBSX8+bvnmuYmJHRtHgDSC4aU6bA73/gVsR9vnpXVJMhb0RoSXRbhTQH9swnRDaBW9ppRl7A
JG/QWKZdBTeoANbtQvLx5xy7WjVnMLXoJOy8itaDBFvnYiygy+xNbvysj4OYmCjh0YsSWfQVG9h9
s9Tm1Tr8soC6im5eKfSyx/4YrXAGqjEZkk1Vj6cdJI/ZkKEESIdldlkO0oOGr6ckI0x3XgtkRMYq
saEwQ4JXw+l/QbjXFVYNXDaxJtRf5CQsCZ6CVFLAH76NNBsF5fSWg90pmko/eIOQ3k9YRPFWNVLl
oDfARvjaY0eslokoLkxnYqipNzKqOd0LI8qNE0Zzn+WlqKPBeajI8tu/7AlU4jeEUs8I8MwpOfOw
fD1zJqHvlMNB95Vc/zmpOQQA5aD9FrnefBpnJkfvTCzIQ5DL2VE6tsFbbgAaBdFJP34cstPdq2wO
DokkIBwjodeGXH5GfP9uKYkZsx9+9Yt7wKeYUO6//kFGVRZihjibDZ8IstxynXawqALjrkZa8uL5
1FL+FhEII5xJQC25mHjG6ApuSxHAEVdj1QppzqYX4bXQ4n+AdQwA7Kd0SeQFQzocq79Xw6o9pk+K
r7709eCgQNuj9FEFwrxh85Bs0lpdWsSH2OjCKyb14yVXZH8AhkvKCmz0k69ibKbLVW5CFhC5kRMt
thJ6zTMirVxXxnSfpg6njY2Lm8xJtPjVnXlVAU0L234LanA+HOPVJFD2quRM4xD2CXwPMeZtaAyI
jGZAackBjzIMmiFthlI2OpDg4TodWWs+bXEIIwlh+WC67HiEPR9xxxplMrupA7kmfVh4XvynvsXA
nkf3ZuFCL9yMw/Nenz7ETrg1qfU27Zg+ta4hFweANQ4xji37LUGU5BkRYHNUAYEeCxSY0irht9fA
e08FjbxHt4SwcJ+OR+KA9JrFjm2/+UCWwsGIoEFL6APv5A+BOdOxKqupeLVWQCI8i8xWtmU/ksPR
bgSu+E+55qUXHk/05oVRD6iOjq3InaceIwamOQqlR+98f8cPUjehwyeo4E9Tb20Qs9jM+l80LS7R
ILWQzknv5TTDziVzmD3SNS4BUXUo8o89E1eSOb5BM5xPh/lOKqN7BO4i1zdwWbhAQzIy/TeSQwDI
gzK0W46shq3fyYQtWwhdbjpDHUFR1Oxon15Ly6vla84wp5SkS6SFqS3rvPEfwk06mPl2IOMLDDkq
i7HvUPy/IRCdA0USZ+JAMBbdd2coFBGLSmIP0AW3ID+HyAK76gWATQEAOyP+4mTijfBOD2+rSnFF
0pv8s+PUqRTeabozRHTPoIjlLzJ0VLn9CEQVkdHjxopOsz54uoMJnj6QJRazPvvxaO4o8ubqnSZX
8WCeVX6+m4QNwpc3zt//JO/3fBIsdI9iGWYHIeyJmaimuVTeRIIwE0P6qvyf8na3Dg+Tuh+kresg
Nc5aDvarNT6iRlaGsHRqM1eF+9VLQIN//cjYaa/8opfc+k+lwjApQLDssWdFpj1u5hjcdmIh7O3j
z7sYUugwFi1GVHFsw9MFc33PP2q6cBP0uOvt+8MsILi4i9Qb4SJOav3AyZTLv+J39jyBev22DkpD
xrm29KWYxS31GBNioDvAvRGBg3H4uA4ieJxPS+D9sFiTR73YQDU/bGOCkAf+I8VhV8mt0fppgTYt
iek4n+Jw4wlgHP08M/eTBI6059EMFyNupOgsivkL3pysTxR6KHVJ9q0gt3TZ6f/7E1HQzhz6WYp1
PLdXHp9jlpjeaTHl8xup2JtYFmCg6r4Q++ghma1Hq7s3s6C0cigPDyvSgmFSJeRPKWt0QF4LVujv
n574EAMV8HdAP234dfZcTywUJA88QXU16uS5uHjis6wkWaWf7I8RLhyHVIfrnjDeKfsiH5Yt8VCx
JztsU5LZNgr0dzkjnotIZKT9XA4ruuGH3J+XF+lZINEJFyTqJVr+OtS6S8ALCpZMRrHwKFpUZ7Ob
zQFhRCgWE6+K3GoCjL34wZd15UI1dEDrfsy4ml26w/449boEXQ6cnTszaJlZVcGMUYp2ZiBlbfcL
zueYJ/Jahm8BDRo5jAmdOi13bmTMzkF1ximghLC33tAHjg1JobktrWU1rU/d4GUDIwi1QDR41YNy
EgNA6aRSKAi2N5MoSmi3QdpxD3r50lpXJ4sJp3aGxOE0RQr49xJKmQ8QXjOse1xaVrUhw9vr42W8
0THOn9TF3J4c4EyUoHCu7oNiH96tmaE2N1cZMHUaIsM17PorttvKqaWEbo/1/nXSvJK/vOxzHI97
cDFgaOox4vJ8r1GI9o3hAHYjl2mWy4VCdeAJINZI5Rl6Ojw=
`pragma protect end_protected
