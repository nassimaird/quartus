// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
b8yHDcg7CBShExUz3XsuT6d0ZQ34DLGZJI0cozPaeLnFF8dgF3acMxix9QiZZCIVwRJ5P39ypVKp
Em7xfUREztDJRLNWCmS4KaliJ5NrJMuXQlc2hjb+ihjwzVZ+j5Q7cRA+alGjTcXDG2PmGorDC7mL
yTK6EZ9AZWwzN8GaQouiYlbTAgFC6OBYbUOSb8CvtM3TDaF8609j1MDLGCuwDMv8gP5Tosl6tr0t
pLroqLhBLCfzxUMeguSCBktEvWcKIN4iy4qjhLpjF+pjFYtp11MFmIueTqT/g6uGebmV8iGaZqDk
GgFyghEMxh2hk513UrvuUxWjKDZvj97f4so0nQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10144)
jY11KUgn3Gbx+3U5MmWhAa1EI3I0l/iVeZ8LEOvJxjZnqLvadDFfX/3pftU2mC+yWEkqMbRVJS7Y
Ql++ZkFZfnHEVMwlgOt9qUq7sDRlKc8oTF3ZeVGgEOFiyMuPk0XttQfMpifYkk0Q9mFGzyCdkggm
nBPrPbloy5cNZYgZlEl3ObKNcM8Cud4x7+7ZgMUXNnHHPTYFy4e67zKenV5om8BAZzMdKrAdOAxo
g1skG9816zcPLSK695ueXnJOeXqCtQQB197rlf622EmlERi9Wh9xUg99cgSXrvkmVxuWWhw1EWmk
B5bXzOBSLFXyG28x337Pw5nv0MFMPMOs2JHezxcM5JGyurdH7rzbpbQq0Cc2entfHcHuRNQVAEQA
lvCDk+Td8PEQ9jitR7bq/4rIwhxleVVg5nYKOW0Q2y4dMusLWPw7BA3bcrKBLETd6p0mXXaW59pH
KWKMp+ct2/QqVZCeR1fnA0KeCaq5qDennAjhpp8xIcWcpnlCy5uV3CliqBI/GeMupyohVkUfy7zN
VWL46YWXOroIf2+zSN1ogmcHdaVX55M6chR/bEMldSePcQOAu0P17NNn1R/8iiJ9JftPUlxeNzmP
0hnHlhFAuDmNC7cXLGjczy15YG1DoOg0u4srPApoNHHXcTL+n5Z+LfxJsPwIBGnH1MoQAQPH6bdM
oufhBcbLIeTHvtUI/RktPNsM1100anwVNDpyxLL8OyZ4Zak8v/YQI1wZhMOChYWRCRyM7OhtWEw9
TTkh0G3cKWEf29n/5wCijWISV5+wkN/xE7x9NU8qTjszMQRsjiNDPgzcQvhqIC/HdeSVMDwlOyTf
d2Q0Vv3ml5DW2kBn5rhKnDJexGhp3eyHFdShiOca0Mcx3UmHOjjTPrIs2hPMJRjXr6cDSvLWdUWy
WMRMZ77LXdf8i2a+6LJIm6v3v13pOWfKYWNBrACKkgk3TdwKCtN3CUchh0cknF3UaNhNi+YQcQz9
WmqPv9Fuoy2khU61wib6TpvlIVnt9tzCYD7qq5ISCw0XRGUDSd7t7xgqGXWFJp6BWZeaJClT1iwE
I/nusCmOjHo2pLhQJlEgX+oYmDmHq0JTx6LMFb//5/cdUzQl3sH15uktG5UIVBuxax4/PmJPlAQ2
7M02L0cnoLV6d6BGsVYrNRg4dX8fqFujYS7PmdT/Yz2ya2MSDKTcb78oy/6XeRP23Tt9mhg2WheI
dAn6o05lvMQv18vRzIJddrcdpqxBcVPTFplsWLWwqwq99Cok+IrA3JYrS0bm252gpyDf7atKqhAk
5zSivulbozy7b4UPTF1Zk+c1r+0Z8Yuzi4yFSneyJBbLOuAyC+2gvPeverNQqSe0WMG2vrSyrYOi
o3lynzI1G05865FIDBhhqAs7lLzMypRFNI/fClI6my38E1nrBNpLhDz2LJfTmmGqwM2U3gBy3mP7
9eP7CViH2IVvkZs8OtSXA7ejmlmWCAvjVQMOP9Wmq7B//CmQuyAxGhHsfMvclbYOpLxaljtqsov3
MD1QcyA6V3fyeQ/mUgartiqskNMYAtXGFxFaHF0DMAWcrqkcWJnIJ/3iFOzJOg63lvGcI8CXP4zq
JI5nJ5ic59MQD9MInk8KdzEIW6Q+9FjxMzu9A/4rADwsNQSMxGvXQ6eK9lhK9l4ylVr+7CjQ5M4F
bBeSdR5GCpFJdezccelcqOAkQrv/96cMVLLH3JYLW8FesGW+SFBnEj74vJCuOnI732a/x1Gj93z3
nX+yiasYXNICWQXmu101GUw2eSIp5yhxfubRQCRgP94tkKc2e4XGR3kJczovWZ3VOqMTv/4Wu8py
WfVjACSpfv0R6QNYa+RpQme8ULFovnJaQLWrxl45Ra9TIR4d0/J3fJq8mkc8eP/QINKjOubLD+Dd
ivxuP+5omw6by93A1HudPLbIcdd7tz/f/Vgf9ON6Y/wpOzv8wbmw5+wKetjH5cB/YG0XDYSg+XAs
v3jNbBk4PnhTC/Dl41W+Jc9oFFZX/zhkEdOOW8sbKAjXbUSXu3aj0PdHGhV17a2inoIWPddFP7VB
esqibM1BvjKVvU9K9F7lmycdVJsbGQUqITABtTXxeELf10n/JkskB5Pn8HA2TOhHfVy8kV1EezzN
PpvO3ZfnbIQUjZJjWnBcnKSgwIOVEFMjbCdMIc+FRWwfAy+JeXOkrwot6CK/flMSCCESNqy1iQMz
W+2U/ibctY2ajZWVNgf2+t4LaMXIbiM+o5E2FppfS+clRwuQcIP946BCShJ0b94yNs3s9VFQUm47
sx+x9fGsL1SFfZOYSV6duk3vvMpbcWIP7rsd01gxXFLWXoaQjBCbb2CRKxp0Vl+v3Z3TcOwYEY1Q
n42btqRz2KQVNq4a/ngopk+Sa0m3SzHRykhtdETkofdhSk3Ncx5Z3OAjhc1NO8bA7WVuMEz1ddyn
17sZAZ9XORiT9RpOay90bZWap7dnIy3GYBOxbJfU+jj9LKG2guZEGaEC2pQvNKwboYF40iNaYf/a
q6y3YluJYZDDFTxYu0Gih8WhdMTcpJOIA6qjCi5cBqrrsetFjddupT1inu9VvoDL8ECJtYO1JL2t
JWcrHJLxVyQjrwpG7PBKkkATflm9Bn7fjS12A9rBEQ/5iKKsQ37ftEc4YiJmFgNHn/+91PDuVIAL
7kCkeZ00RRExJD+shlVcsaI2+8U0+xL7m9U/QAv+8KqgdOHpUjQVo6x9oq6blZeRsYUSUp5oELUf
xklelbatep6S7RISwCpSehTCmsHeVm/nwB3WIcwsOHKUyWFfQNLXYZELxZPwX/y8YNuactUV553y
bu3xixeUwiJ6PlYqOoD5Cw3NJrubWNVr+hKuks/Ps7pcM3ZVcukhyyedZphLCLyuvTdkHxeafcno
ZL33JhmZe2yap4OExMG8BEzuRjF4e08V8xFP4ZyMbrs750GFLxJR8D6kpofnczZyIvLSifcdj2W4
cjy15BvIY5PyQC0Jfj3/GvFG6cHwLN3xz+OzgmstBUHn+q1ofV+8P4lquKDYbYM786Y58Ag5crq2
ZcMbboqxeuK/X2TihmvAEgFfY8sS4XQTSPxvSKo+94e4Tdm7IDAQgp5RB0O9fFKhOvrsb7FB//7N
5CnWgfnpFuyunXRimxRHNAZcURYFBw0HNi6EuGxtPFGslD8m+c/LDf+bYzLp5d0EDGffJFr2fX4E
1zA/J1urZ+ZBaBCVM/jUBSfbtzpQ7RRDOCZYNI3b8M9x9hDAqmJ9zcQamysIepPlj30x4D6KUkLm
cArtZ9cKe2QdLyj+p8zkXkPSQUiwp9o9f2UfKaICi6xjIBo0MrFlXxjcJs6LJROM6sgADZ4SzKJ+
0a00QUtWoCWZnGd7uBkgVVRrG97eLe8DfEAP0rgXJ5YNlSfwoTNOkQnLQw89brluQZ+mV6fxj4l1
Kve82wTeY6PoEW+40L7zlBzn6pvqION/DPbWEYi+zb+6csWFnPrDZ93FaPwyYWMpttik4v2uPb2/
E76hi/Ai9wwIJHXprtOEopMvH+W+0LLH+k1PLhMvLM+N9HqcaIZYTutI4uNUJRUKoM0zswB/1EMv
bc50D0ZapZYJ3XA1DueiGRorc5cC9MKPlyxiqNhtgh5mJx6Y0oAl6jeS0zES/perWH4Ypa9kJxOm
2dVmuQSc1NZ0J3yEkibZ4UxhAOe11Guml/tDny8RzRBYSMvM2zqb0O+wgfkIY1ZZOwIfzLq4VTqY
sUIte942Nux182t3UdMnk0kxdSZWbRskqg7YI+xh50sU3+1aV8bfSr8OYJ4JuXN2hrfSvWGHSx6o
pKFUBdcgx/vZgegtKVdMfgF8rrulqKkLnC/Jdq7rYwtbbxNk5EDjj0ewV4Xf5OaMIpcwGBzghdWt
3Vlr5KUOTtS7Xo4+yTKMUk2M4kER9WoOvdQyo3sVZB1fZdF5jijoWJnXL/gTG6JQa9n8c42g9FaT
a2J+9mmFIgVUqCylzO+yToN0WXoaIxUYD820lsBl6LXVzlYehTiTi8/flBx3DBEm6PU4IY6Ke7DC
x4p/zIkNa1uAno0wwy9IJ0m7najI0Uaz0+jnkpZMB32d3GhCQDCfP4eA0UVqqCnWRj9+g7GGYrAH
UvNy446awTTvyOY4VmlceK+v8Lw3SG41f8Y8j8jCaz5pR8qZ/qtthBuUzu26tH/3V5KNtdz4Ylgh
YmdAphGXCAeqOgapYtP4wucStZ5Fp8J1H8+GU4a8y74K6UGB5uwH7DYveU2UNKceLj1gEAMPSCVE
bhGiAD4qHbsjJdNuMJlbi1x0mT/5Zj0QwnHsQoLE7h0AtC+cil0Er1u9olAtKwKeaFbiUi4YjUkv
iJGqygE4tECja85QP88qt78ZdZWLN57cJ0LNj0cZb0k9re3M/UjznfnntJy8Gz+X8MuFIk/zoCVy
fyGa29lPjYURs5nn/tWpsaebDeU9N8uRn+fWoqF4opvRgFdJ8L2GdUW6eEMNsh6Xp0ZwkyK3FrjU
4AuXt2iDOugBgiX5pMgfEA7NugrHM7zYsLDy5kcE8SpiWH6LTuUNlkO59XTJNpc8NzhosQejHecH
xX8hCtiBtQ6sc8Z9pYDIENrFIZiDIRRlyroMe+fjgGBzt2rcUvvvRXZ8S9Lm0W0wDgsrOWTabH95
PZTpx6CQcoAx3/iXsnQBzHazFpYF4ZHjsndZN3UEURq8jw8UpdUFhZEIppl5vsonogU4vX9PoAQZ
KldoZCTLPlUNGxd3vgVOt6aHbWWWFOtbRehLzJgZkMbV7XYgnlaYrCRC0OPr+c/r/D+QbJxydK7j
1/6SGjmXQtAcUQEJ4XXKeFJkkot+ctIuc54d9unM36nOeJo6X79gS4+rsIXeT6BQmFj+oQ7C9en2
w0c25SCwASq5bZ0bVuhpo5cmwUpY/iOzc1vVUqZl2xO+aG3DkxDzMVTmDNTZrRdpuAIRR08A+Hbi
Zvu90RnVg8N4ABaznBi57033Ptb+zQgZNx19JJQ4R9JyAuLuGtgpmz4brwZ/tDgHOqB/sZCTSxnW
m5njEl+Z+6CdX5UE5fXpQZnmFTP+zMXOJ/G6GwxNyIwI/WCagyeKyotdSEc+GeN3iyXZLg9rmpdo
USBMoiUkf4+Z5VbEGP1G6kAhnc3yFDjlEmvUo47/XP4GWTx0n1mZrzUrS55W2lci3x3f89ze+jEE
h2CNl58vp+SnfkGRzkbOLeG7+HPfl+fsm8qJTlzHe2Awy35AJolFIZ7/SOgWPWEBaJG2VH7/eX7U
t+jh5Cu7x1C176I9teW0cQDf+uR5+EqKYmxoCkR809L/z3AUNHKAw7KCXr9d9TlgHYjhAq8H1lqF
NNFDkc+OkLkSqoexZWy3/JHMfZ9LoyRKtyOlhK5KZIIAo5ZJOpIOywR0355yTM95TtwVnvJB+AXo
+v9Rs/UX05q65XMg/8R3phypzBbssdv/S1czxKSQAPwXuC0gy4ar9Lo9scaUlT73VjcJK3s5JbO3
2vuQU8i8YKVQWGETZCuSDDEJRKMlXaNGxZmMoZW1LHoa+g+T5CD4qkxEB5CxVtbxXQZhhZH+7PPH
IgELvc+GnsMwj/Aai3h2fqOou7mIh3AKlTdQJkR1NwePbYsGG7ljjjUzVYuHRlPIAXrXIAzLU18L
lMM0RZVvfkPXih2h1QE1xHZc/utSsfFgbFXShz7wxl062rZ+UmSSwePwfb3B/dwDrQt7vd74SKkk
ZOKjN+I4J7IC4xlIXW+OwQm08g1jZSpNBQGKRg+y8SZOxpE551qN4LiMFzXM9Cy3Sb4nOtJJxxcG
YgSxSM9RO2sbKL3/e3tX0jDZb26HIgiHdTecu6XBkwd9NpBtyuFveBU2nx2uu+XtgEDOJw8SipJK
iBm/lkrKlJ57fbQ/eMMEjhCsLTfwacr/u9X/BMDur7/ns+/jC7b0TDVS/cESaq0VOrMZjdPa86mJ
r9rOY8yTgQjHioDK4ud6yWIdV5OVHv7H4kIyl3rj4F44FpugFZkfZzjwGHDHD71FyCGtwdTsQkOD
t+qXod2jm/IMQEOwAm3f8lgp+NWZQowqeWdFKnLtqVsY3P/m+V0J2MpCACS8qp5k7iC+fuOxyBPI
6ImlLDrZ+gKFcREncJHfmG2W8uadzvuWoAC7nKmtWwDFm7tfXlNg+kciUnsq4AlqJNsvFECIc+hR
ijoEGa1Bav+ouspIeSGxLi4yj1eJLhswdhWsJHSWoPC+YEJJMFTJh0N/oo0BUGrfIRcdB6di0iHA
Q0Q7Xt7Rs2ETaTJI0L+9oW/QKbEr7wHyhDSHyG0bW+SEcOOXs6QS39LWEAwUbkel8tRT357pbS+J
zQSsBAgMeYxunUo5qHDdvqoAnLjiMMQ6hVgV2UFjO3Dr/3Ftlc/w7mecLvaxFnyGuzJSLCYDQvBc
F0FQxt2HJQgtIiuYPxuy+uQeHAwGqZU2SXxvRlCkqNd5y9F4+JcVC8cWyqu1utVwoog/0rPg5GQF
2TdOyiS1dqIJXDkpa6o8jqOj1KZdy8JGgac+f6ld7dbSAszLmBDSQdp8h552KP/gfae0YiZmEt00
j42sOBNfMSueAUzBygMoygdmddC/BXU5HbRjLGaBtNGNLCVjBdjR+K6uoz6AZkKYrLA+0pq1+0oI
+dCeJvmjlUv3S3WwdMfJWUvLV2Wr+0s+CHReZWNt2Xk9+gpak7WT+gpShYFAy7LXedtoGOe2DigD
kZHs0jjpv3OTjJTMSTzIxl+KH3vJckEPGT9OxA9wTajn4swfwiPfi1LMAGHR/v7NyR8//SYb3v+e
J52DTbI4r6YaSNlIRHdOymKhPC/F1up47Sqdgd/CkOBIYkRodbxGv5HifbtlnpsNXFQaDV17YAre
QimLjWsyz5ajwWij7tOZ191efwIP/vtvo8GdM9bkrdA0+MUDIg55xGj5o9Wd7gpPZe4YuPuFF1Lr
ZzHYbRfAEbNKOHCm6MlHPoMol/5IJUvdLGN+k1sdZyASB7xr0tHK3f63JygWIgEV2f0ksUxy6hX+
uXvvYFpgXtYQ8zpLb8dgbIXHfTsT1osila7VTb9pvLY8Udu7ARsjHV4aPQSdEuuS4qBFho/ifCD8
v1WPn8OSH5Md6JAHm270yePXj8SULQyEFJXCl6N0WNuVx86r3hXW6jfPqAvRHIusbrRO6YHk02xR
vVtfbPKTjlAPAYW6L0xRz/vKF/0v2g9ctuN07M+T/esMIm+4N6i7Z5LrFPkkWjwBX8goxVez6g/D
id4FKNVd/LEVCY4svjYInfcYe3ohx9Zxhf9gYvsh9o6XTu2njJ3+8UAfLy0VnKKHGjoy4ybZb4q7
Gt80WJHmH1Thuha2VIpMtn+GYgaUXNSrN0wKokFRukikDEfYgI8/zYUXT8MeYDBaQLKsIQfoXsak
C2fCZfKI/ceqOduw2B4RL2pr1Xgi1T/T9ekYk5M7qpEBjnhoc+mxTI6sJJ9I1Io38eEvifq0sUHQ
A+DEgWkGhzdLvxpPYGCsnVTSO01GnTXjRX44IzINX5efpVgv4kfp9d9ws0EAJdBs6E/+Am1aOiu/
y7CBCtjxn9/QtbXXGXgHcb8Tcly+dZG6bj3FYZZRGJcTfB/JuEr1EmlwF8r+52DchlLGGr4UHagu
7OZ0X22ciIwDAp+acSBdmjRYXR7lGCv2WxDLSdOYbGc0avi/1bhwSN5g4OFYlHjLVpe7q07yN1IL
6neyaLca+wLwRNJXElB70Jz2zebbXnsKUPR9ZGxetLzbHJq+s8ps5JNsqqH9jKMzfiqhxi8hcdJx
I2jDW6gXhnIqD5TKXjyk03ao5xdRPZhwRGAZgB18EkEpRokllm/bJGOYeui2AayoZ88zsbgM4jod
ihwYxH+29C4jUQ6qVDIjPVtP82gVmRyM9vVEkQWWiPLzRW62ipnjExhQOTyNeTpUYncxHm6vgS5W
pxZbPSqZHIsQI2fr+RHl0xx7yChB7GM9Vf/3nPFpsvxoGYLJX4UTsvIcLYXyVSzjMrJs48OiGee0
8oYep1oxj1gpT98BLYHZMFCrXHlJZIweY89X56kH3YOXpWpXVpv7AQlMjeQ2ZVu4iHnqStudzjed
e6ps1g/7NjqYcS2vNIyJiB1ZOIdmi2EgkQYMkcNpJzf2BkSYtUwWufSJmXLR9pVERkzS6A3Nz0Te
+7Jj6tcNuxbdiZXQmz1pYZefdGdhfwbs8FRsn9yBZ7ss+Kh9rH0oygmyqfdqOSnOtGAskpqAOMcS
sB/CnWXzQI6mm9UiSVJDUM451DFLLGVvmvA3M//1GdW74uAMAa2ecjKm+4F7l2ofKlYCONPw2/BF
3NLRRo/N2rNm8+XYthsDWpWveFtEBRHgwxzuFRmRRgEFKJLiiB4J2J3wXhSdTQ+tl4SQ1EM/Z9/L
L6cCXzIwVOkL48dz0ForBU1CEQlzoIkM/jkp5NivFV4VhJ2vI70aQJgH9+yXIgPZ2wNYr7YgzqyL
dPQWFRwRaNAQ/WJyWw5/WvWmCVy07hBqy9YXEMvo6cmO0dRS7hH7mI3PvnC2teVNUgNqFbLP+Sqw
jxe5FjWxkxsylOTZSmkypngJlj7MOR5epSvDfQdH6SH7ubWcTyg3Cfoo/p7eocOT91z+CIE1Jx41
ccjwMSTQFkpIcFcDXwfiAvYQurimS6p6E5+zEFA4rpIyc8qY4NI0QwbqWmSB1dVlGvGQAF/m8meL
10Ha8qFS8QDuZNk4xpCVYBBfplvJDqSZYk+z1CDR5IMJXeWLxuPi2W2WU+GLJ4RFNFLqLpcTcxcY
X2ltQ7z6MrU5CLdSU85XzeWyX5fZTRimGRbiSWeKY5hk8tu5LHYoOdnNBPMO+Me+Z6fjcOmKhEFy
RPFfzO3S8llWzBfg37rloAhp3DEwvMtQyQ3qRvAll4qLIaLh40BaDU07piB82z/0gT+vAi9iqPzA
ao3fPmsIcxnAWI+MxUT4pcyvqOu2MzazwSUo9pLOnIU4ah76QWbJ/BW6TezouQ44QOYJeE1wDGny
PT44xG49I1NXlU7kInRxkdXnGvPp9eMyHmxKz9kF4dyxKjAj+f6Vq0MrZlbdsQ70ElFaUBURrBzA
cpwumACHqXq9JHKDPE1Kx5k/JII/vvWMbevoSqrZSJBW3sNnEJleqhi04v1ApuINGUnZOblG/wnU
UAQy+tDp0tXdA+aGMo1nxPvvDIEWafLtQPWujd3gASHxv81EnZsb/BQN8q/QAoOXRD0A6nknGOiF
A4Hsul0onxisp79/YvOivIRTEulBUu9wPapzOchpa7VefnJX1y+69Uu2dp65c4isLwaMS+k4tAbq
g0j6Aul4B+GFCFpHVpsmHhhy1CnsEH7cS1E22+RXHTcSG2NbfynG/8f7iE3hypIRzd7yHdu9IQS5
W/7GbfmIcEFsEMMVt6WyhSOovZkWtNoM2JIVCT1bZeNhALrz4Dlvqony+AHx+Ct/JVuOrDjcEZvF
F5jkZcx94uulktRG2tLEiGtM9gUZHSOxRuC7WhSDuuG7fW6dbBB03O/eWH+LTvBgHdSd+ED+/IsN
MhT+NWlkDxdJ0ZFjJ6x75Tnqc9wVuKoeyEfQQwo+tGzD73/4bLy8tOcqPExoWEgI4EUlo8rluubg
htF2Oo6q1EzCOh7C4eZqtRwI0aRJOavIXd8C1rYrNJiGLlbQlmGmPSmVp9mOgyHagoYsDti5NTPS
uFnXxkMALnpr8v8ifI6MK4mpM9CAvyjm4AAq4NizOEhcfV3GkDw0/LtJLiwsIOL/PP1cgQBmJAHu
7WpqJvb6OGYZx8N1M4DoDmuI/zIBahwbgxfR/5KnKpSPW4RcQQM+qyB6Fatb7Gt+lkCOeUUfr/bM
WvMULOv2mKZWeK9s80biPuygnJhn6cLrmOx8fr6weDk5JdPeqE65U4Fngxb6GhA8VzM2lh4ZdIOk
4tAsn5AbthTMLyIwp48VbcojwwbGmsCzt1ltHC+g9muZKiWPZFvMzHqOuzXwETVtbUVek2dbTXqZ
iJuXcI1kdntt3agNF8/aXoPIZHBliaplGZe1cDLsloVn+U6LkSrh3ywLDLT04w4cqj98Zk03YbqH
GG5XSDDTWYzVr+Z+d1JoT35eCL7rl3r4/NGabqKrCRFFYbmLcmE+pH/OUdIYD1FTDHgxMK4/iCOC
VbNQfIBx1HYbHLqBwSOkAYqMWGqtnC9cpTUAM82b+6WPMCa472pdV3joJ2JbCFxq0MNLpmyBXPT5
RsMz0oU2pVO46SPiIQ0ajmJZiZan9zncgvyUZQ9OGSlDida8arGwNwxg0XpaSHnJvavnu2/uBmIX
XnY18MOmxzmjBw1YU3n7vw5qZDQNWJx9fpAxRCRqqsWGe77LFqSr3tdcvLnnZv0AKlxkecwyOM+u
WNbwxUfiDvye2sxHwk3d2XhtWCm0ez11Pw/B5HiZ6FqlOvUxkjq2LT+CzIvb6mI+FSn9U6QMEvhw
YAP3WrcXvFjlTgv1xtTBClF5DgDcCt3GvSiPxuT1QK/rtGTORYr0rNSaJEO+aayZWUZEtuVsoNbl
o6ASNQ5ED3u5KQs1kkWho/IN5E4Sl4cU0P51T7i7djojr+VZVnxiyyA2uNeFNNEwNgU2LmrQs17V
8oWvcFPxLrzfG5uLDHlgOUD0GbmCdtrEiMmliEAUdOMOArb5UE5v87nLIz2+T2j/DrsF3tViEG3B
7kD7UQzTwyaVtFrx0iii40UXkm/3jDh9NMkKk/ZmvcyLetIZI4m3W2Rv6OSDZTyaJoIIynGcJUv3
XwO8HcnzYMFdh+/hSMaifCGB7Ns2otxSXaiy9uUyjh2L7sIYmg6CAIL83vFNJuhx9fw25R1Fb5e5
bmBxQyif3YKOISEfrOcpSsk0WNY/4bdf/4N3UrpH9ixEO+txgC9tHLj4exAEUSeiFP5EtsBU54Rf
tdP4mvAtu04oSKqMmCvXMrqln06y9VcxcXtI2SDy8bdaLWfoRep5reW9osC1jnP7KnWs2Hvzkqr4
+o7VfjcJTZKtENRy/MyYiLoh5BhDl/03/ZeDi8n0Aw8EgytcRnr1lXDewp2nswsM9UHgg2cEfndC
Bu5QRFVIhrHsS3dER9hlyqUt5wMpN/Bv9nW/zWVY24EDv0YbSdsdrWulCnLYfCU1JzX7JKWI1uMx
kEP0TMkgRk7t5Gray3VAHBO/PVSulMsMRQnSB5psjIdYsKy5TUe8FdYwxECXYp+QcTNlJgjpL1zu
rhzDJ3IlboI1QFGoWlmdZ9Wm30F/sFiWMOqra17EHN5KWBA/ByqbpKpDumbk9hGo5EXJF8zxJbF1
m/gLrmn5dLWC60ZuMmP8ioa+VGkExxTh6xHqvmZD2qy68qB+Dn8p0/rT/qNCl0Y1yDyMVeTkh4js
uG38O7fVsiTp5or11GPjxIgGQFndY1w46lmUcHS1orT581qdxAqw+qlPfpjGRL69KzFs9/aP6UWE
xz6sjh93nPrCsSThkQjoMIgeHGqhKhvJq2mnCCAvIjqq+EqhmaBU6QbR6QOBQ1Tr6Udu9446gfUW
nJsK7pD/Iqu+lH8PZMA4lNIn2RyGGAOus7FRhLoF0U5CWUOSYw2QG3V6wzniSKMtXsjLPKL1MqW4
LxUWV8qmvEV7F4mFU7oUtOK0PEZe8pUus1mS5EALn+XU4qb2qznvxYNQXKzL2lK7MnKL2klYC/B2
6wCdGQ4g50hxA4eRlY5ovNiY8tLx4bD7ZGotWMhMg2HJnCSho1wJwnD6RmlMt2Ra8+mi3U1S9VAC
rleK8+HnhhzNLSN4MJtxBTIxodreVCNwNYYwmUO3DSKpyXHJjgCdMm+CHQ8QLYlL332ZMhvBD7Jd
TKEy/WpoXK586V4E+mrVyCT2bOXMiuTef4xMVP2C6SyonE1rfplIVzT3cRtz3uSfoVkCL7Y3gt9d
olE2UJ4pPOlbjitjsAmxSkafdboH4f0vbKD/leBEzvUpyLzTfc6+LPFZRLTZ5MlEJ9JQaf0FXY9m
JNgQ9p7AD0peJf62+RG4wMT7ZCD6/dKygBRzSuAjOeSjltyG2QI/6CTG5QtitA/ebkBrI3zr9FTO
uiumPwQbYvwtR030eOPk2ABfx6kCkGAlJRkTCm424LcoZVhAco6EWtLiouNByC63jkmOJwwzFXji
R9tFoeIXvfQJuVxX8RnE9aTtKAevU6YTY7wbPre1lBjfapzgrfaQGr5PTEmXm4UP/3SlZoAS/sMR
JldGWZ7WeN2sraB98ap2v398KA9nHy5272a753Ai8m+6/povgV8R7QKYubU4H9ENwpVs0BbIUORl
GUFiVf6ECocEVzCqkIBvNDlnKKGVjOdADk12VqJsq3tUTIiDEc/6D6mhD9ZkEzucCudRziw3rSA3
35pLZY5DxoVZ6y7Bv82en3tuny18PRs38iUuN1m1KSrKcwjEj127CF+nOGnGbT6a8bcfjgJJPYm1
PCadULC/GeqrrRG0Ck3oyV2U8X8LtZ2BxU2KkdhnZEXEL6GB5MsTY4JhexIB0CFeKKDUxrp48mLp
1hul9OxkmTVGL/+w1TVs9Vh3n2L0FBOV6aPIsjzBtUQ7nmEhY65u8paUYQ6uInNwfg4iqnHc5OSu
tIOqarPzrsCiFZtlEFeit1TMJV5EMpVIcc1ZcEMbTsD2d196W2+KMn5eWxpNJYnOEvXkPGN9mF3i
eCjTbqgBKy7f8MGpkfD17IVrgtmdy5bsJAGVqG+MNJ0nS1YPNseDmN+Iy+69CF+EuQfVherQO83p
giD5QkeZWfwUQAcV4527B2i0ZRVkuZU4UxXaRxxVWeo3D+j7yoaxxwe7v3pTjvY7zJhX+lnfWS2W
hH8E2LJS4aGSGt9JvoNMUUUaxbWFzEl1LjdEpg++QkHnlW+mkMXxxzDFh/bmUUXBFaSUaGqEvefw
4Mo1sQPPqLVezOymsCldBSeyr5hI6NgUBKDJIMRy5fjxKIO0ktdz+qJQdo4UC0VSG/K4ga8FXQF3
EnnXtmmru2vfg4xDKhCUlDg7S7snfnb10GuBIfOUUZRdh0lbCQl6FfLwzpe8y+w4SPznvxRcw0zf
7cZ9XNArlGM+j7Dig7AaY7ZjfadClkBiR8ctMfJc3kvKbYogs92LmSzryKG7oWanRJAREb+vpW26
AVzmby30TnR5euwt999GA+Uuzvqw1e68b/yT0U2d4HJjK3oxxcFglnDkuA65C2KaAUeHJqa111j7
SzX8FFNcMfB6L/dq0P3P+WCRKHbdZfQHVsgA70lK7mF9dethDoygvgerf3bPawBPHEjqGhUvYRld
ExeluD1Ponzy3xdgY4Ij/sPFlel58sTK7tNHeZ312/ulMdvCGAg6P8A5AUNKr3iyz3/WITlscbG1
INsh9RUnVu8a9US7cKYsCCI0pcvZJc/GdEu7R1m2TrbqJDGz7WZq00DVFPb2Tcefl8KHMyy5ITxi
z8Wl5KjFslUzw+ad3cVl3tYKNFAa+i8R42mG90qmRJyP2l1mcRNPqVacGr1ouRy/bsn04iGibMoN
FNioJX+3FxRV6DNpcyhgWwGWxowyYt1p+MYzksl7SHvZYqtFdApJP3xNLUvmf4ZxDWwl+hN3ZA==
`pragma protect end_protected
