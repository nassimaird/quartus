`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TRkWrp5WXkmjPY9h6boIqPrLQCZMCl/l8Jgv5AQJ2JaMDTtkzsWn9YIKzfYB+Be3
zE9llXm040lsAQXib4TiNyTFeIdaxoW11TrjJSs/uo9uPC2aG0gerGWWE2fdEm6s
55Le5nJikHZQX9Ot1oNjCHBcceWOSp9WEfglQ79I82g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9936)
HpbL50h7vjNMi/gPRE52+cexilJCi0wJafJy7GWYmfUwvqRwjObi+yylD9aa01FG
UQ1DcwUFFFpXLfBO53RPrmar0eDiQ0h0xflAuw30MTZgvl4ctJD5vmhHN/OcSJfJ
J4mTHudogyA1Z4zy92OMuCMv3r0o9jswg4AlIZIA1IJwhNzBwHNu+2PmPijzgMdR
9s9G1rfiT4W7RFD6y+j2rH+MHTGMjJUPiancy3Ap5mABbJqj09+CyArl6o4bHKmh
j5JUXoNjObkr7xYazGqaOPL2rbo+SQO8m5JAjOsJuhoXgqzxxYPla+gtGed4M1Xt
5ACb+mHUM2xrBtVW8zPnmul7DwgYT4vMEtF1NEOa5opC32zDbQ9QiyGu0KpRY/PZ
54hj0NND5YL3MieI550k0Cw6Qwwo8JHTuFpJO3YJXkq0f+JyL/ER+QrT0dNy70hU
BDmdnGv7yFcFHj/WZXdOrYG/n3CvFS1CFiqAwnKZKXOTrKU1meP0vH6iCAeNMlXZ
ErW7C1AHoDyV7GJT1qRWLjHul1l32n0nG3WebLs6EHm+HoeHGcqfu7Z0atS6MuHU
FsbT0AXhc2BxD+sXviEw8ciMgyAKtWpZEA7Su194/ufDXYiQ6IegpjIOws4NHHaN
tQMrsA2m11wJ/cZH/HAqv5HgALUk5Amy8V/7gTVOaAQBQE42IsYabYyfjQkCI7fe
uwHm6lsGXRHgbTW4JDWp3oL4BpjHCzjYQdUb0l/7Vs1k1RBl5NqNNNU1LCnRhuCG
mzC95hJ3HaY4ctd8QDI0RYoKRRftl6kT/Ub+Z+mNRbP+2I29SsHMGxqhI2S1rb93
uocv6+KhB6zDSNkan7Y+vjwvXpDqHfLrCbhudNX9gMUEuhg4zaCVeG3Jrm/MhlVI
jh6udkd2Q8d7pIW2Fd+cmHE0/QL6LGx4xuIUhleD6dbJ5suqiFhxQ4JmVnl+GY/Y
2fzXpuJIK9VG4JKUzHwgezixjNm8pbX2ai7kITyxjAE8Ww4jvl1xeU/8q/CtGwOX
7E3N+ySg9sNQHwtSa/n3LKBe3w5uWRPCLkjLNrMGFfJ1+L85730kBG0tV//5GWLF
BVGI2KJOM2UyD7Ye0gHrqqhj4UOhRw9pjuf/b4UTUOMYsgDY/6IRz+aNgk65U40+
iBifV0rReBUaR/9bCK4ENCtuiArhzSfloGdSQgDM2Ua8smPwajAzmKYkM6w7hxt3
VOyMik7TL+jgZ+Mk4FX8Liz4xBHkCs9FZ2Vlh6lTk3qpHkY7Y9zsDJvVLM2R9zyV
h6GVao+4l2AhBxJ0GaOsvXWdWfPF2BX7nY1wkPziLSubX3bQV5QxJfeidE8pkcMq
L5xkTy4Q0K3SeOJsX3lMhcGFqT8o+sMhLCj9smkyOCt7aUrJ+eBn+ytiSV+DL45X
04/0uRWHKPMURzYl8FxjXt71YH9ihLAKJ/9sP+D2OodQh4JCe8RpempJmXnVtuxK
uDeUYIyOrMYzdXbfxGGMVv/tm46ASnJB46R5AAItiwVvycBIp8Y62WpiutXTMc2o
zr9Wew1psz9k6BjlGGGChYJ0YhyXiEZ5LWyGXttMoOAwCuv/1LBlrzp6yS/pLYhF
g1MYPjyQvwVsbTIGzeYTYXYS8PoHQzBz8eKQ/5PKZOZA0rvB1u8wKv8o1BeuuBK9
cSs6UjuCTBiIQKod7tjV5vyTbzSP8ojCnCclTEj/PgXoltX1NuztNMdQgOomAoGj
TMRSgpP+OETDQ/RfGsl56dF1rNZJuzd7sz92KcP8BTPC+RmW79siM2s6q0jf8B1L
HgWJKNKrqjvfL72jN6pPkue5r+y3ITFu4Hf979hMnk/ayNx7WlI+ozEWw4sb189N
/ib6QEJ2EzpLYUl8mdi3bUBFS+2eXokDhHcq7aucerK+O5vkxYQiUhaagzjoGLRL
QYXxMEKkN3axxnMcF8jvqgNJZtwB9gEQVDm4dwOXaGq+vHxAAHP0lMIM/4Tbwgfz
FVeWgPAdsff2Lffazo3lxUsTpbqeF+MBfhcL03tYb1nOzPLCPoBUKRAh6Jm5vek6
gZ1Ba/WEwdinKV45BS7bZp9JolZtx6QzNOpwxhGm2MLOyFgLbCh0YeSgqn6mhIdO
lQLrRfpw3QzE8wEHjH0wiOVfFnjGht8169g2o1qyc4yfrNJCVBd/Lb7pGpmhKkHW
DqjRRXMCb/Xq5X19mBtPZSt/jIbzLlQvUidoVYm7upKELzSdwhNj7mFBAntpKAYE
++0RwdCbfrb9hUtmPVpbw7vEbgEoXVBGDbfJw67DboBym6o+vJRAwMKIeIjV0jwt
P29UhJEB83evW1KbGZM422yasrzRbYY7h+xEnARQHoh++9TCp5LlpewOP/+PhTaX
VHBpPWxBBigTgoAiYL+5R5u8JYtqyMqIKG+DiX3IDLKIHOvzbChJDbo9nv8u22ZT
xHhn4E24dZIfmY2HM/5lTg0qyeLdjX7ZrLjughhe5z70Hd+Glj9oDpcqI/dg+wvx
fH8+Ye0I30DDkolwLlIqxZ5zNSqjgwupYmHJgSL0d/J7Xd9MxJ1C6Uoku+AlSEGk
JgaiFHhSEB6vAGQ5pkqEd8fSbAOc0/PWBhCS6jyApbBqa6DU0bYkIxuvRoInOtII
/CVyE1TW7rgYkUNUbbU6RZgAuBh9vv49ZcYmsxkkvkCEQ3HZ/eukZYcNJN6GmA2h
z4z74EUSRZa6OYjufqxR6T9IKKjVfH8FuiwvLN2i52eJ1j999/2nYIjM5EDtn8WO
/cvEarSGOPvefUHrD6hl+rJttUDs4WiLhmF3LUpgYMNBxIMo3CARIoHda7WxWDKr
RIHZoLoGkPD8es3t6aG+orrf54HRhIHmbacINLpXp9AVYEKEAftLoYJ284gzimS4
8uPV4BXaJYN7VzGydjcM+30yWq5BJZqvu8+1pz5twhFHTHW+LnB02k9sve4ISIjJ
4hd2xvHJrRVc76xrzFdw5FXSGwvp57wnIgCG4/uDRcmKdfK+8sOSMPKm1U8BlDXu
1U7K/NPyzXF3F3o7np2Ej8vklPuQ6UnAULvQGha65Imm68ge9s9OG41SojlTCO17
VlPVFtRNyCXx/RQZEB2HMjdhrONKIp+XUyzXBDacHHXt7wlBn3R0DIMMHcuDCF3Y
icjotzCXg/+2lAFyUPtmFBy5d2cfU34Mma6K7xYdjyjWml+3RZQSv/av8KU8Dd3/
W4gB1hrgyTHDiGGZbHZuoxr/PC7FESwOcQzMU2C57VC8APlDHZcacRaMPUBETSzu
EFP4P2G1w0hP3RJijz+3qJinlJteQyUzEjWEhZc5TgQjtzWwOpLSrcTCG0RJaqHY
RqBbchzFADSNliIWAFmUMDl8XpQX057gdg7QAGBCQKJ4IyxnNltohnpoOIHK5091
xFCzz5aXuqtEF68Pou9u0NC42NSbZEL4lRQIwK40W0/GpFF1aiOPExxn2bkPLPua
LtJ+Qotmvi2734z9Hm4gQtkAyH+32v2n6EkARttdw6DM/wj4sTELYezLxpQEU2Pk
CSzXLlgEuhT+CSJ/UQcs4NneSOKm3lG8fjD9B2n5ztiU13GjoQNAJqF7v3xnmKZc
cPlWuHUta8fIHBgXZ5h3pS/GhcD/mLIJSPUIeXMogfvUHmd8BcLUk89fBBpudYwW
JaQ4v+eD0nznC5rgzi5rhG6pgLuEeDQvwk1AVDxwVLoXXW3UcsvSdWz5aO8TZGjh
Okja8TS7KgdIsgnSz4lQAyXaSSXAgiJ5wxGOZ2EwKj+aHuxpWyd5I45vfhJVOqXZ
1qNkAFHHvoTWfKiywd7aVC1mAod4ADobntBGH5ITqNGopbg4SyrD0DnfAasfHznx
FChnN3e0Hp8MW4vlLjDZOFGjJaniaLK7v24+IVh11TdL3OOKDdbXLLzLa53SySif
+g0ECczSiMulTczkorMOfTB3rKGwWFtQuJGI22kFKcGX+idtF7LLm6xl5x/PmTLH
0t1ctrLgHFK6+wICg02/BkrmHsOr/LSJz4Yugb33K/4tkcGJnKadcIvOxetcXDB5
PEP8RzcFZsn6TrkqFFjceRDRMmeFQ22+vLIbe8ajngs89xO1oscqV0om2wVVVxOu
Y0zynW3UnVoSpaojBwWXEXm+YqniJoA38F5IA54YL78oSVzODV3UpVx+YskcqYIf
mR1CUUPPl4C46YppHG2962hHL+5vD3Jg1psYEPeNelUV53DxHK95fCLNcayWaAJy
XbwosKNuy9SqIgg4nCkET9VkXlccigowRqtMjiqEBHksKM+/jmKCsyRZB8WW4V3R
liC4KQ3KAD3GYCDPgu52j4Hu7I+lTkVoHsYLFngto9I+/ZorXdhvF9tMOyV6wl8T
vDVn6CSEoV1cZtYssAoCneBgQl4jePD5si+3n/WrkCK0aQ+ZjwUzOi1Hy+09A6xL
7hk7HcPCXNc/T/CKG0DRzRqQJ8QwA7zM79TaJd10qFknRYSXLf+Iy+oxd7QiWMWq
P3FlG+4nP1P7NBDc9cpxqCidhZ6nz+KBWCgMLPBfzOLN0qv4UBjVWflpvUqPpMhG
mBPcLA/gQ57ich0x2nuxAS47BC99q/k6/AXtn+EN6/kNx6NSybl4ZBnALemu6kmW
kXZgWnsNyEYNdIhE/k7W363nRdJZl0HTjQpPeAd82S2D+5ESxduHBn1KKtCczfrd
QeDgXZubnpweCOTM39q7RZbHzOw6+PNqmm6z6cesCwEDXxOBha9B1OD9+7tOKe3O
xKEGyWPJI1KH4qAng3J6jOb14H5OtbrIzHay7VaF+x/GEFlPn+B/YbEjyKATYxy9
6kMQLTdsq68JPFtC8gcOH2iyxD46F49HrLqhLpiKzwYAycxi+VeiFX9E0J9Fz2Wq
adgQHue67P++abhAqhPMNj2jzijmsnBCuWkqYKuvuwOZh5AJB7GCMWLjLvA9LjfK
kjz8At9kbGPTKJWW6Rcxhwpx1zfgXXOgM7oWWVKYQOAjU3PPbMm6XmI4iMWi18NV
t2MK4BAoP51MVGmCwwghqdYgJEHywBeta94UZoE5+1GhFhYVV7cmjPPA9fhOSIcC
PzTl/79soBaW72iHuOEbkhtXL9i+kc2ief5OQqNegnGsn+EHr5q/lYBMb5/oDOB/
B0D8QvlJwKwOWcwUiPgrZLTjTiGr72yhN7NlIRFeGRC26Icyu7KCN5BlJ6ZCsGds
/iSLY16NNuZFHkpuwTzyEex50EKyBqIGn5xGg1QfJW8Ac7jAZbcHlUTCbfA9mJFB
lGqc4fJEcvXL2xNNx4ZblJ8qAl9WemtMofW8BL/8G1iQAs/CFT5FLGJlPrmpLvAO
82b7Yd2o3k+eOm4vDP2lCeHdtaBzlQkkuLp/oYwXvXihu40mmDXHODgjEclAbNZp
2iBBqwkhANq68jN7VT5PH7huCd9XwNwn8rZnTUrtGI5HRLDIO9ZU94UpRrztrwDx
PNGKeCOQfcwJRtMKzGaSm8TWnf4ihAKJaYxJ9MahE+V+OIJf/yLy59cG+H9m3D8Y
nnqQmrKKkcvvb+HuT2uzRybbLWhpFbXX9T/+sBkG5WN6BNPsk9c3dhbGTgP08vOs
WvmY3X3/PVhsesHcT8F6XR6B+/xp8LAJnNTy8K4V0AV4hhQXzoX/SEoH5Wiaq9QZ
6Fesl8+1f/d8VrMMh+QGmX3NCUmFyefYfT/D2Pru2DJk1LzRux2Rfi6x3HPk1qMV
/FmH1z9tfqbnHZCjSCZv++SbNGIewBO+Kf5DmIL24e3PyxTLQO2nVrb7ZQ2VFoCB
wQrWzJP656CfQyrHcOFvv1rvqiDuXylPzHQ51GG0gpSg1c3qeoHAtt6LxjDIGdBy
tnKCMJCRcFP4dfC8f4725MPvPDjQb9dUXgwQW43lDPrqkohhrWe2qlOM5gdAJrfu
aY/AyPDviqI5JG9tZ/a4JhCJa34uWKoM6kg6Kz+WpHEHHIxpBzzTpPBSn4AEeOia
awyc7J6LCLFU362HZh7lDA2d15hik5/PshxoarM4yr7LvsCNYH5oUPQauGUPAzcY
+XUmX9niq3IlJF8dHEwr3rvb0dHJjBrpPNhzxrUOCFsjtS6ZcWtR8eJcT0OPoycL
sFGRCNsXDrIRq2y/Z03rQ2Kof3bSS5ADvThZyRDhXzbq9f5RMQA3OTAn+5AyKT6s
9YxqnB/YeBkyU1OkhKRz+orVH6c7049ph3doESTCDjLhc4JxDWs6rQVLE5UqnY5G
UXfkNkNz210wKBz/t+cf9mZEG4FLsw5K9fgDwxXJ2GAIJWLUPLpDP/22SiL/mS+U
TnHW23QOtYIqNLcELfbKYg8TLR4E13BfH24+fRBVDS0eXZZI38LySczgGm+Abjwp
/Ja/LsLPBOxFqwMfbb475pO8cFfP/gDZ7KDfszfkSVCzLMy0fmnbpn0kXBIdUELd
Bav240oAS9UrwOgDW3bWgaBOyyqqAl7n1+JHlJjZM/1sDRFR09IgmTqQOuKUqzM6
wkyl0Hpv87v+P9GLBF7u/rEM5Er8zNOiqnL+xua6j09ZaLq1tolxzylzo8eJ1k//
3Xqs8HiUT32BvjEO9bdjkfh0klbQ+SLJItUL9PLPewnBF3QWNQz8CITOnbJGW+My
5Z4X93joVwv7/9t+ogtUkuVnDVJnxxERWcjucZp0WkTarr91Ogw7LoQzT7+nt0bp
ziIvosHw9ENB47jED94NscxTUw0PBVbeRwsoCyQDchRMQx61lCryK2b3YNFqmLFq
StQriPqE7nXFCIW2udOVPNJQxvjGysLw51Lna12LzyKCRFfgHHFFY9U57jzQ31Oo
lgWusbIqoA8+l7Rla44/sryOqdsxhtpighwxmsbUc5MnJBv996jKOIkZY7RQXVl0
RnGLow+FJXvUVDE3aq1Li6xtslSNgSoQcx7NXUihYAL3D2U6XL2GLvMD7wd9V6Yd
rMencDPpIXBiCiwWblkY1lXizJ7MfjlpRQ0kd2miIfrLwyqI3GNbbeoTbuamDF4h
mYdHilRkm6h/YA+rREgUK/QdeDXOOrA/aLDDRDFiFs/xDKcc2bdkVVGYgdBYejTv
ZR0gusNHunkzhPsXXwGmC5jzIIHC6iEaHB8ZXHTyp2mJfIAWZqgiXpRkx6HujOHF
3H/YizePzhJOUL1UmsxSKPDWYBp8xnuRj3kOAECQFqc4GVBOd43grVJBG3WLhXm0
T4iM/aDxB358+5MuO11UF8tc6N7YUM83J8LuZeYVSPOIfaxwz1Ah+p5A8QsFerr2
i9sPBnlBBOtEKqX4/Jj5qxeHKu5T2oMNsAB3cRbzaKhJ2wqoUoHHRXgVRC8P/ohA
vK2rlX+G+6fW0X6bWGX1Qezzt95Iy63JaXDmVSxLY8MrVNBWcx6qZ1xLdssD29CN
xvVTHa5EV03bbu1KCkLkEvIBpjaTsZ4PZTzC0wuMf63JnEpLgg1lEWgDA856T2cW
vSObpjItyGZkmKIUiS8T5Hy4Ta8BqZE5YQr7++SRy/yqX2eXTr51vGNZnmyEbQKs
bl3VidhLOHjXNjgDZtklE/ZqNGDoVoMT2FS9Ak0ZoJ/STRi/7PxKgNxuTZfoHse/
15jCrlpgDFDiCIJS4RiNTRsDfnlbC7csY9Qo4G9BsM/SHmEQTF6n1FcBuKdRy55c
hPH0nlHn0bbu+mWWUugJ+hmsmObQCLYKnUNcE16b8xxhZV3xSOyjwDXRXmtM8CHz
l7ejDquCA9N96tpw5XCFeiPzDDi9uwXUAoLFe1cVNfRZe3HbFhFW0Dwf24kxQzZl
QLDS1XdwofNYibGGu6tnmJmVM/wokzL6JcJHAyYDAbb0beG3YyNfkkGxEYTdlMJy
4/C6zPk9PLw4LD1+3ld0fcKcrY8KLv8fdTWDaw1oNihHEBN4STm0IDwqUTluupDZ
4oqD6mW0gczrshc5gvMlKX+ibE9hupnb6d0QIitdsIGdFxIAXHBbvKYnAaPvAPjJ
c2MBPCWaR/S5yZ3kI0TUSo04sL5ZWTt43wkFt+Hlx3n8byWsiKamaN8i+j5eXy8w
VTWDuqTuOKVZSVn2eoKhs5UiZf390+5B3nO4s2yyYZnEuBJ0FbF+yUXIcqkHkZLp
nyeZqG9aycKlIl/hQFgol53WjWqSi1/pd0ZxVyhRkdUaC4TlpSKXvYm06sT0+epp
tV0Dx3tCjN5RsgSJKq0C7Q+oWY3eYdP9X0JDmXDaRwSwv/0LAm/s6Tuk0YX5mEHF
QAZppIsx5zrygXMGQD7ughE5OjNMmKrQ5v8Rs+l1tN8xVJghwM3B49WBSR+t2cyd
9/Y+Db85lrg4WAaLmABgVae5pNVcWXK52BYG+SZosAm78MxMacEdF5OWGrCS3CL0
b4UMKSvgrtdpCcBwm8WAUJNqY/qIsTuG754iZuARuu36g5xNFjR1ay9pVeevyx3A
1sERCKoaAqn1ZEnzKJoygFFqEAWGPJidHdKjDuQiROk8gd/YI2xV555Z8GqB1nbA
qW4FAnj1nPEP1+3JoB8+w4AtRBa3YvY6FzjDsYcwT5FH0ZqIL5Yqll1ISLyP04PN
Wr+8OOMvrKq39/yo2u6ftn7yw9ruhrWiolHK8I8ielUviy3xmvrJiVHZBKHEOPM4
36uwFhS7OuuGln0n0bYwt05mOV5rhZwkwbTf/d1DubR619YKY5CB0O8xWzOISCb2
CCQyVrq3rWrXhPOg8ugcXxfl7Pt6u+0ThaSkqK9xjfkgNU3cJ5D+owNDxoCuAHgs
GKitEInclmnSznStFq56c7CWagxbd4JAWS4YjOLiLsTAhy/Z7b0IcQ/9ikEYSyic
nG8p4MV4bCVasIy2mG4mvUPubDA4bXQMTN73zxSUzhPWcT/SjE6GtNczOmI1USu7
vVjYqr30qzHRVh7ZPgt40lb7XMj9b/2fx3VvV2hfXwtVMxFwyzRGdV6XO8ZJ3Xb1
ce/6MgH3rrfvyINOfy6TsTLOiFUzWL8AwY3G5ciiBI9JY+9Tf9uydNvwLu4f8t05
J8DRFA326F6+hKK2eTew3GxwmNU2IguGHqwmGldJat0CyS9HJm5iylbfu68FEdn3
EtCf2qbDUlpUKgzlHAS7QW3kx+Qnn7okRbZZedLVdgNnMCGiylqwE1YmfvrPZLMt
5gngNwNiBmrvUgExIKxsq1uxbzHKIlR7pOGbgT6f3wkvSqf/P7X2SFOtWsaKh+ok
6tP5wgZV/ryMIq1oOWQOxyZe/a/J6PB/UjDkjswoAbo4UFyRVaDA7kHXzcEFOVvM
5IUpmHnjLNmr4t1tPnOzW/JgHF2VslxCCrJuFFeJIXeSHkSPiXqAme4PZMwZNRvg
5prZNvYCfazr51SMyejnfZ18akKebJm0kJ127HgdETc8Q4aQUmD1u1GocS31GqrP
cJj63Hw6HWFuSB/k1Z27W6aYJI9Jow++h9kerheQKLBUTWEhI+ouofApfsQohs1+
V5SPHAuxsFWmlMgfj9vZtQR5WJ9zOrYukzxGdrJMRAob8B+EP0Sbj/2md2ZMCZP/
py36JL8UTuWMqM7HfpdRu0mFcqZFJxOmpP0TYGrrSwm/A3cNWEEY9F8vhR0D4zt7
Dm58gQQ1SdrULWH9TtnhgVsAPQuozB8Mjo2EwLawZEUIKJCr7PQvTqLVfkrVzCZQ
7AaCQDDKNgZvWNYg43ijeUrlXK6DfXVv2VNLCtdegmk3tG8r+fhK42lFqBVXduVI
80XAewl29oApk3PPhfckXYZAeFFHwqjwE/2tar7d0z6QN/84O4F+5op1Uf5USH/m
Horf23zcAuRM2dQha96P0ExJECDwTDXeTJ+KwE7+F6m1VMtx8UW8cPaVostM46m7
cCH0ACPvXHZrKqWQThp7a8yci0Hu3IEmJbWDnn4jXqQHiGhWijz/Rl63MDZ/ECd8
3xypRsv9ZOPp7OzdandVVmTbL26G6iU/WY1Ed1mZdcmM1kDzHvSyZWasBLIzsCj6
/mzgO/qcI3rvGE1dMpZyfGp06MhSx7D2tknUQ6kN94SpTKvjBWOdkzUtaKuX3BQO
A/cA0A/mc8Howfd5JSu40z9nVVMlNnhYRVhhVSbgvnlfjb9PumZ4grX3wegRnlOV
5qUofrM/fqGYJumqjGZNue0gq9DbDfWX/0S6EzH9s5MEi0CDqF0YDmyGqJQksidl
Esq5IGakUarETZ5zoh/X0djVH2CxJbqLlpQ5fTEKHIrqtW8iZWi2AKNxQ0ag1BAK
EZrYRMYlVRKneke4mdAypQj7TzcjMfIzoJooxAZZZKijgRYsdjG+wTDiInn1XQBx
Y26LEgxmhB02lt0J2F1/eNl0MTvofmF8A1fNmfxsufXHYd16sAIQnBc5v/WQ/Gn/
Aq+oJUWBWdISqvIV83j4qrvjhU4yh85BoaR3mtMeVTSrmblaRiyM42G3q3k0CcEc
6PIaWKI9j0bqx41nm6bjBVDKfdTpOnopdaWxepoX2Wl9508vCGg73loonhnUURjw
SQBw077y7LX6UeUjsYaN4+7M4aOHoAoUMUbP4KtcE2a0JlrMeUPHYqqDoV9H6FZT
nCWp3Q2ljEQJqkxPgIFff/nMOGeLqWb1bznQnW0qVCnsVQhNKlOrWU4i76DkM3DI
6i6K7Dd1eenyCgPgcvNjzr6CK4mbTkRez+TM8cHNpPR8tMLFeuSETWQM8aBXC7bE
r7ehfnJnQRHpzyTDgIm0KC9Mj9G0VM897qnIuhCIGBiJedMRa6MUco9N30ei1NWI
qfOAojG1jvq0dF6sFHkX9TlrtzQCkSQUtiHUmCFmX5OPGLjk6FJwNELRgMY8LRXi
LuI0hZMJ1Sgfp1FdNHE0uy8c4y66Cx9gCwGOAvvIlG5U1jQT/qGedFGyYYeBKUMw
oPl+3x6HiS3+n8uAX+s2HKroalFkqWXo1ax8yGaTrnqujX456mI9s05RbtrZa3uG
Es6kz+TFaPIcpnBM5kBLGijp+F7W67Gt21R6NHetrfCxxO1IM22aIDfMAkmSmLzF
OkdZEjHG076yhSUb6LWdamZ7u1/wUwm3l35Lw/+/5DQ5tP677wZnnnHJWj5m0hcd
YnUhaLHMiZkzp4Qwq800qskvs1tMjBW+FmukXg6AMgCyVD90FHc57QuD0ti8l1VC
9J6TzL8O4OUfzu2qfvXANmhCy0wbcfx0EbNylE57LCzyzdv4T2W4TDe2EvC2MCIg
CJ+5+y/+6F3klSmwRAfHDGGp0zDEkeMWNCKAOx501I8tGqncdyBVE0AC2pgj1NC+
LKN4M+qhtuCmrXgkz4MZ/5TaFjgDL2jw044VEbmQW7x6YtEH7KAKRoMOPI94hr2t
7x2c+ot42drsGB8KOua1KxfB6/L+/p0mw16QrwTFBZ6wZj9RpPwUWAyoX2DoZrE7
Awqc8dpHLU9UPYhMEpX5tmCJ0IGcxnHYoK+f7BJ8aqyNTSWZH5VRP2+Vh4iLwEyn
Gv90DqCyczsmbpgYtqKEVo+c852ebNWE/lYzyhGqQAm1XxMJBmsHKYDSo4gd4Cfb
UjdjxWJc93vMV8gY1FDJETPBK2lCqsS7CaIJg+dmVAnOUAMEkijqjE7NbztwidaI
Nwc8gbvkDIfTzmMhSWsN/7o3hIA9Svl10O5ugT5vDUuJcq76Jh4jTWQqT0odXT73
QeUQSCGXdP4dYIMi6qGmxx5VRNJPloLsFsBa66mnAr1RGoz4sHSM7HRp9hM9hlsc
gKjkOPn8ztZ7sZ0mRNEKmQY694SeSF1GwB2lY2zEYm9yYSCswKawOOEjmOSOPcLH
MvrPI0q42CzSdaU34WrOilOrCXmXmDiJv9SU5hDkuKdpJ+oKxA9+MNaWc13AfrXY
Bh9390nmj951yOjfUwWDFUwmTg7IMlXFbpuJYL4Jwl99G392IZGEgUoeqCMd2Zez
CeacaSmnLqceNZGYk6wuEoM4Vvzb1U5C1tA6cU7B86Kkro6WBnVGHzzPJjm6+u03
eVH2MKbp1QVVWWOEHRNVpRs7hl50hE5PLR6U7GwQsSnvLBa7Pce2zEy+P5ns/XMg
+HDRWTxM+juBKAr4i0OGJLn5EAPI87ZQBNK9uATN2P4HHdATzxITon+E+0K1Y3eO
ZnlJuCBgCXmW8Nj5Kaxm34ns5HnjeIbokxg+HqDq+sMLaJmU0achamO4wlB3VMAd
wAgyvsodok9Zqz9vzYI5Pt9/pbtFix0bjqyzV7LYbJ2H7wjgDZZ4FyOtV17WEinv
nB8NiSrFmDDoNWCTR6EW/c1DvpUFf8eUXO/GT+6+R2XnZCNHGVP1RjDOj5dk4j9Y
7sFE1yByCJk8kbYiZCT3T8EtQI4cjC3Xv3Uu7cpR7vdZn0F8uMte4Yzvlszh6B4D
TnpDzZ8ESqUu7nzAVDNJjhUI3D96//iERv1oZPWZfNLa6059B6h0DHM9mkF2IcmA
dJjZ4kjzDzejvHxGHvCk4A45+FoZZjcExXwO7WWSzIAHFm9kXtP2ybFTJltY3Jng
+ZMvIJ7W45cssMdmnITJHyB+JKLdBcrE9x+M7QT59ZGTFJDbO1KHksKZW57KzuAy
hr5C9NDz5e3U8F38ZzT2f+OoQqYyPsevohCCyuZKbwLLSln71/2oFOGOqkTk0m7F
AyRBcBhBbd2F8Ne5yZZWCkcItZ7Z1Qd2ySah9I7iAOtB5Uyn421yXgQooNaZHvTF
q3Or1sEBuKf+8spoHibEgPbgE4jT2x+Y0U+rz/eHM4pXu/jetSpyZaeclIMqyaPm
8Gj8Sn6367kkZuiZWmgNrMhlvMpjoYWWT4fdSQO+j0+AIzt701Nld0TQcJrqMyj0
+3cQEcr14YzEfrDSuSErzPmLL+W/yhWiyqtqmUjT4x3ZOEuI9LqFYhBgzuX6iuRH
t1WJtt7WpryKDmADQWpp7w5x7sTwy5mm0YVy4RzA7Mm7A2QbE5sdw7KeGSxCS8Me
U/d+xGtvKBpamoxeHwnqA2kw3ikJs6vhKqK80XzSPBkEB5kgXoOidffcCaIYb5qR
9ZKYKP90wB/u9+HSF0GwDallRCVglcfvPRpamPUZCO9Tew3Vs4bpSN6RVvorlGwa
M8Eq9Frs2AsRfMWl4wEotVWcmLYyBy3gxqrL8zoMAk2MHsg8drj5DvAqAM4UB4KE
aG/Fil/sLgR2sHukW5gPnHaxYVgfebASWZxUUQk/l1Rk1uo2z7irHA2RqN/BXUK6
JlSkieaRPpWDCTLyv2RBPHUe8i5JdgJlKRhD/f978ftvH6MZm4nLdqKQPfhZHk4z
8/Gu+A/W6Z9ah1a6eYpQJGfL4+FFgk2WrohEC2z7PZtXPX8c4vc/3ZhIUvXCMXb3
`pragma protect end_protected
